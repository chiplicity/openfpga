magic
tech EFS8A
magscale 1 2
timestamp 1602874640
<< locali >>
rect 41095 47073 41222 47107
rect 36001 45985 36162 46019
rect 39899 45985 39934 46019
rect 36001 45951 36035 45985
rect 23891 44897 23926 44931
rect 26927 44897 27054 44931
rect 37691 44897 37818 44931
rect 42257 44251 42291 44489
rect 24271 44217 24409 44251
rect 33419 43945 33425 43979
rect 33419 43877 33453 43945
rect 36219 43809 36254 43843
rect 41095 43809 41130 43843
rect 33051 42857 33057 42891
rect 33051 42789 33085 42857
rect 23891 42721 23926 42755
rect 36219 42721 36346 42755
rect 26341 42075 26375 42245
rect 41889 42007 41923 42245
rect 21275 41769 21281 41803
rect 21275 41701 21309 41769
rect 15393 41633 15554 41667
rect 26467 41633 26594 41667
rect 43303 41633 43430 41667
rect 15393 41531 15427 41633
rect 28635 40681 28641 40715
rect 28635 40613 28669 40681
rect 36495 40545 36530 40579
rect 24915 39865 25053 39899
rect 40794 39865 40864 39899
rect 28635 39593 28641 39627
rect 39123 39593 39129 39627
rect 28635 39525 28669 39593
rect 39123 39525 39157 39593
rect 40819 39525 40864 39559
rect 19567 39457 19602 39491
rect 23247 39457 23282 39491
rect 42291 39457 42326 39491
rect 32499 38505 32505 38539
rect 32499 38437 32533 38505
rect 17049 38369 17210 38403
rect 39497 38369 39658 38403
rect 17049 38199 17083 38369
rect 39497 38335 39531 38369
rect 39215 37417 39221 37451
rect 39215 37349 39249 37417
rect 25363 37281 25398 37315
rect 29871 37281 29998 37315
rect 37783 37281 37910 37315
rect 40141 36703 40175 36805
rect 15439 36329 15485 36363
rect 32505 36193 32666 36227
rect 43671 36193 43706 36227
rect 46431 36193 46466 36227
rect 32505 36159 32539 36193
rect 22937 35479 22971 35581
rect 28457 35547 28491 35785
rect 18883 35241 18889 35275
rect 22563 35241 22569 35275
rect 33327 35241 33333 35275
rect 18883 35173 18917 35241
rect 22563 35173 22597 35241
rect 33327 35173 33361 35241
rect 27295 35105 27330 35139
rect 18095 34493 18222 34527
rect 23615 34493 23742 34527
rect 16399 34153 16405 34187
rect 16399 34085 16433 34153
rect 39899 34017 40026 34051
rect 23575 33065 23581 33099
rect 19383 32997 19428 33031
rect 23575 32997 23609 33065
rect 35173 32759 35207 33065
rect 41889 32351 41923 32521
rect 43637 32419 43671 32521
rect 46627 31977 46673 32011
rect 16899 31841 16934 31875
rect 30791 31841 30826 31875
rect 46431 31841 46558 31875
rect 20085 31127 20119 31433
rect 27997 31263 28031 31365
rect 23575 30889 23581 30923
rect 23575 30821 23609 30889
rect 12667 30753 12702 30787
rect 24995 30753 25030 30787
rect 45971 30753 46006 30787
rect 20361 30107 20395 30277
rect 34713 30175 34747 30209
rect 34713 30141 34923 30175
rect 28819 29801 28825 29835
rect 38755 29801 38761 29835
rect 43723 29801 43729 29835
rect 28819 29733 28853 29801
rect 38755 29733 38789 29801
rect 43723 29733 43757 29801
rect 19843 29665 19878 29699
rect 32965 29665 33090 29699
rect 15203 28951 15237 29019
rect 41889 28951 41923 29189
rect 15203 28917 15209 28951
rect 40635 28577 40670 28611
rect 31780 27897 31848 27931
rect 41797 27897 41981 27931
rect 32499 27625 32505 27659
rect 39583 27625 39589 27659
rect 19383 27557 19428 27591
rect 32499 27557 32533 27625
rect 39583 27557 39617 27625
rect 30113 26775 30147 27081
rect 34615 26537 34621 26571
rect 15611 26469 15656 26503
rect 34615 26469 34649 26537
rect 27905 26401 28066 26435
rect 29043 26401 29078 26435
rect 30055 26401 30090 26435
rect 37875 26401 38002 26435
rect 27905 26367 27939 26401
rect 46259 25993 46397 26027
rect 22753 25687 22787 25857
rect 26887 25449 26893 25483
rect 26887 25381 26921 25449
rect 21499 25313 21626 25347
rect 37691 25313 37818 25347
rect 31309 24667 31343 24905
rect 28543 24361 28549 24395
rect 28543 24293 28577 24361
rect 14105 24225 14266 24259
rect 14105 24191 14139 24225
rect 21327 23817 21465 23851
rect 14139 23137 14266 23171
rect 19659 23137 19694 23171
rect 28365 23137 28526 23171
rect 36587 23137 36622 23171
rect 37691 23137 37818 23171
rect 23213 23035 23247 23137
rect 28365 23103 28399 23137
rect 32499 22185 32505 22219
rect 32499 22117 32533 22185
rect 46799 22049 46834 22083
rect 21005 21335 21039 21437
rect 42073 20859 42107 20961
rect 17095 20553 17233 20587
rect 45293 20383 45327 20485
rect 21275 20009 21281 20043
rect 21275 19941 21309 20009
rect 18613 19839 18647 19941
rect 45879 19873 46006 19907
rect 22293 19227 22327 19465
rect 24035 19159 24069 19227
rect 24035 19125 24041 19159
rect 17779 18921 17785 18955
rect 17779 18853 17813 18921
rect 38059 18853 38104 18887
rect 22569 18785 22695 18819
rect 22569 18683 22603 18785
rect 40884 17765 40956 17799
rect 25455 17697 25490 17731
rect 28123 17697 28250 17731
rect 43303 17697 43430 17731
rect 22971 16609 23006 16643
rect 33425 15895 33459 16133
rect 28215 14909 28250 14943
rect 25329 13855 25363 13957
rect 29929 13719 29963 13821
rect 37375 13719 37409 13787
rect 20855 13345 20982 13379
rect 19159 12631 19193 12699
rect 19159 12597 19165 12631
rect 19343 12393 19349 12427
rect 19343 12325 19377 12393
rect 20499 11849 20545 11883
rect 24961 11543 24995 11781
rect 24955 11305 24961 11339
rect 24955 11237 24989 11305
rect 38111 9129 38117 9163
rect 39859 9129 39865 9163
rect 38111 9061 38145 9129
rect 39859 9061 39893 9129
rect 18739 8993 18774 9027
rect 47259 8993 47294 9027
rect 42257 8415 42291 8517
rect 47443 7905 47478 7939
rect 34799 5865 34805 5899
rect 39675 5865 39681 5899
rect 34799 5797 34833 5865
rect 39675 5797 39709 5865
rect 25455 4641 25490 4675
rect 40819 4029 40854 4063
rect 32079 3553 32206 3587
rect 35259 2839 35293 2907
rect 35259 2805 35265 2839
<< viali >>
rect 41061 47073 41095 47107
rect 41291 46869 41325 46903
rect 41153 46597 41187 46631
rect 40877 46529 40911 46563
rect 41521 46529 41555 46563
rect 27972 46461 28006 46495
rect 36068 46461 36102 46495
rect 36461 46461 36495 46495
rect 41613 46393 41647 46427
rect 42165 46393 42199 46427
rect 28043 46325 28077 46359
rect 28457 46325 28491 46359
rect 34897 46325 34931 46359
rect 36139 46325 36173 46359
rect 30205 46121 30239 46155
rect 36921 46121 36955 46155
rect 28457 46053 28491 46087
rect 34253 46053 34287 46087
rect 41889 46053 41923 46087
rect 30389 45985 30423 46019
rect 30665 45985 30699 46019
rect 34805 45985 34839 46019
rect 39865 45985 39899 46019
rect 27261 45917 27295 45951
rect 28365 45917 28399 45951
rect 29009 45917 29043 45951
rect 34161 45917 34195 45951
rect 36001 45917 36035 45951
rect 41797 45917 41831 45951
rect 36231 45849 36265 45883
rect 38025 45849 38059 45883
rect 42349 45849 42383 45883
rect 25329 45781 25363 45815
rect 32873 45781 32907 45815
rect 33885 45781 33919 45815
rect 36553 45781 36587 45815
rect 40003 45781 40037 45815
rect 41429 45781 41463 45815
rect 28641 45577 28675 45611
rect 30205 45577 30239 45611
rect 30481 45577 30515 45611
rect 34713 45577 34747 45611
rect 39865 45577 39899 45611
rect 42165 45577 42199 45611
rect 35541 45509 35575 45543
rect 43361 45509 43395 45543
rect 25973 45441 26007 45475
rect 27997 45441 28031 45475
rect 29285 45441 29319 45475
rect 34989 45441 35023 45475
rect 36553 45441 36587 45475
rect 36829 45441 36863 45475
rect 38117 45441 38151 45475
rect 38393 45441 38427 45475
rect 40601 45441 40635 45475
rect 42441 45441 42475 45475
rect 44051 45441 44085 45475
rect 32781 45373 32815 45407
rect 43964 45373 43998 45407
rect 25329 45305 25363 45339
rect 25421 45305 25455 45339
rect 27169 45305 27203 45339
rect 27721 45305 27755 45339
rect 27813 45305 27847 45339
rect 29101 45305 29135 45339
rect 29647 45305 29681 45339
rect 33103 45305 33137 45339
rect 34161 45305 34195 45339
rect 35081 45305 35115 45339
rect 36645 45305 36679 45339
rect 38209 45305 38243 45339
rect 40693 45305 40727 45339
rect 41245 45305 41279 45339
rect 42533 45305 42567 45339
rect 43085 45305 43119 45339
rect 25145 45237 25179 45271
rect 27537 45237 27571 45271
rect 30941 45237 30975 45271
rect 32689 45237 32723 45271
rect 33701 45237 33735 45271
rect 36093 45237 36127 45271
rect 37841 45237 37875 45271
rect 40233 45237 40267 45271
rect 41705 45237 41739 45271
rect 44465 45237 44499 45271
rect 27629 45033 27663 45067
rect 29377 45033 29411 45067
rect 40601 45033 40635 45067
rect 42441 45033 42475 45067
rect 25053 44965 25087 44999
rect 28365 44965 28399 44999
rect 28457 44965 28491 44999
rect 29009 44965 29043 44999
rect 32873 44965 32907 44999
rect 34161 44965 34195 44999
rect 34713 44965 34747 44999
rect 36277 44965 36311 44999
rect 36829 44965 36863 44999
rect 39675 44965 39709 44999
rect 41245 44965 41279 44999
rect 43545 44965 43579 44999
rect 23857 44897 23891 44931
rect 26893 44897 26927 44931
rect 30389 44897 30423 44931
rect 30849 44897 30883 44931
rect 32137 44897 32171 44931
rect 32597 44897 32631 44931
rect 37657 44897 37691 44931
rect 24961 44829 24995 44863
rect 25605 44829 25639 44863
rect 30941 44829 30975 44863
rect 34069 44829 34103 44863
rect 36185 44829 36219 44863
rect 37887 44829 37921 44863
rect 39313 44829 39347 44863
rect 41153 44829 41187 44863
rect 41521 44829 41555 44863
rect 43453 44829 43487 44863
rect 43729 44829 43763 44863
rect 23995 44761 24029 44795
rect 35081 44761 35115 44795
rect 27123 44693 27157 44727
rect 31401 44693 31435 44727
rect 35357 44693 35391 44727
rect 38669 44693 38703 44727
rect 40233 44693 40267 44727
rect 22293 44489 22327 44523
rect 26157 44489 26191 44523
rect 28733 44489 28767 44523
rect 30297 44489 30331 44523
rect 32229 44489 32263 44523
rect 32643 44489 32677 44523
rect 33425 44489 33459 44523
rect 33655 44489 33689 44523
rect 39589 44489 39623 44523
rect 40233 44489 40267 44523
rect 40647 44489 40681 44523
rect 42257 44489 42291 44523
rect 42349 44489 42383 44523
rect 29423 44421 29457 44455
rect 29837 44421 29871 44455
rect 33977 44421 34011 44455
rect 38577 44421 38611 44455
rect 39957 44421 39991 44455
rect 25697 44353 25731 44387
rect 27445 44353 27479 44387
rect 27813 44353 27847 44387
rect 30757 44353 30791 44387
rect 34989 44353 35023 44387
rect 35633 44353 35667 44387
rect 36829 44353 36863 44387
rect 37841 44353 37875 44387
rect 41659 44353 41693 44387
rect 18756 44285 18790 44319
rect 18843 44285 18877 44319
rect 21808 44285 21842 44319
rect 24200 44285 24234 44319
rect 24593 44285 24627 44319
rect 29352 44285 29386 44319
rect 32572 44285 32606 44319
rect 32965 44285 32999 44319
rect 33584 44285 33618 44319
rect 38669 44285 38703 44319
rect 40576 44285 40610 44319
rect 40969 44285 41003 44319
rect 41572 44285 41606 44319
rect 42625 44353 42659 44387
rect 43637 44353 43671 44387
rect 43269 44285 43303 44319
rect 44164 44285 44198 44319
rect 44557 44285 44591 44319
rect 23857 44217 23891 44251
rect 24409 44217 24443 44251
rect 25237 44217 25271 44251
rect 25329 44217 25363 44251
rect 26709 44217 26743 44251
rect 27537 44217 27571 44251
rect 30573 44217 30607 44251
rect 31078 44217 31112 44251
rect 34437 44217 34471 44251
rect 35081 44217 35115 44251
rect 36553 44217 36587 44251
rect 36645 44217 36679 44251
rect 39031 44217 39065 44251
rect 42257 44217 42291 44251
rect 42694 44217 42728 44251
rect 43913 44217 43947 44251
rect 19257 44149 19291 44183
rect 21879 44149 21913 44183
rect 25053 44149 25087 44183
rect 27077 44149 27111 44183
rect 28457 44149 28491 44183
rect 31677 44149 31711 44183
rect 36001 44149 36035 44183
rect 36369 44149 36403 44183
rect 41337 44149 41371 44183
rect 42073 44149 42107 44183
rect 44235 44149 44269 44183
rect 25007 43945 25041 43979
rect 25421 43945 25455 43979
rect 27721 43945 27755 43979
rect 32321 43945 32355 43979
rect 33425 43945 33459 43979
rect 34943 43945 34977 43979
rect 36093 43945 36127 43979
rect 40049 43945 40083 43979
rect 42717 43945 42751 43979
rect 19257 43877 19291 43911
rect 22017 43877 22051 43911
rect 25697 43877 25731 43911
rect 28457 43877 28491 43911
rect 29009 43877 29043 43911
rect 29285 43877 29319 43911
rect 30342 43877 30376 43911
rect 35265 43877 35299 43911
rect 39221 43877 39255 43911
rect 39497 43877 39531 43911
rect 42395 43877 42429 43911
rect 43545 43877 43579 43911
rect 24936 43809 24970 43843
rect 26928 43809 26962 43843
rect 27445 43809 27479 43843
rect 30021 43809 30055 43843
rect 34840 43809 34874 43843
rect 36185 43809 36219 43843
rect 36323 43809 36357 43843
rect 37013 43809 37047 43843
rect 38485 43809 38519 43843
rect 38945 43809 38979 43843
rect 41061 43809 41095 43843
rect 42292 43809 42326 43843
rect 19165 43741 19199 43775
rect 21925 43741 21959 43775
rect 22569 43741 22603 43775
rect 28365 43741 28399 43775
rect 33057 43741 33091 43775
rect 43453 43741 43487 43775
rect 43729 43741 43763 43775
rect 19717 43673 19751 43707
rect 16497 43605 16531 43639
rect 27031 43605 27065 43639
rect 30941 43605 30975 43639
rect 31217 43605 31251 43639
rect 33977 43605 34011 43639
rect 36645 43605 36679 43639
rect 41199 43605 41233 43639
rect 41705 43605 41739 43639
rect 20453 43401 20487 43435
rect 21373 43401 21407 43435
rect 24777 43401 24811 43435
rect 26617 43401 26651 43435
rect 28641 43401 28675 43435
rect 30757 43401 30791 43435
rect 34253 43401 34287 43435
rect 34713 43401 34747 43435
rect 36277 43401 36311 43435
rect 43177 43401 43211 43435
rect 44097 43401 44131 43435
rect 17049 43333 17083 43367
rect 23213 43333 23247 43367
rect 32137 43333 32171 43367
rect 38209 43333 38243 43367
rect 16497 43265 16531 43299
rect 19441 43265 19475 43299
rect 22201 43265 22235 43299
rect 27353 43265 27387 43299
rect 27629 43265 27663 43299
rect 28365 43265 28399 43299
rect 29377 43265 29411 43299
rect 29653 43265 29687 43299
rect 33057 43265 33091 43299
rect 33701 43265 33735 43299
rect 35357 43265 35391 43299
rect 36829 43265 36863 43299
rect 41061 43265 41095 43299
rect 41797 43265 41831 43299
rect 18128 43197 18162 43231
rect 20888 43197 20922 43231
rect 23924 43197 23958 43231
rect 32321 43197 32355 43231
rect 32781 43197 32815 43231
rect 38393 43197 38427 43231
rect 38945 43197 38979 43231
rect 40544 43197 40578 43231
rect 43336 43197 43370 43231
rect 43729 43197 43763 43231
rect 16313 43129 16347 43163
rect 16589 43129 16623 43163
rect 19154 43129 19188 43163
rect 19257 43129 19291 43163
rect 21925 43129 21959 43163
rect 22017 43129 22051 43163
rect 24961 43129 24995 43163
rect 25053 43129 25087 43163
rect 25605 43129 25639 43163
rect 27445 43129 27479 43163
rect 29469 43129 29503 43163
rect 34989 43129 35023 43163
rect 35081 43129 35115 43163
rect 36553 43129 36587 43163
rect 36645 43129 36679 43163
rect 41613 43129 41647 43163
rect 41889 43129 41923 43163
rect 42441 43129 42475 43163
rect 42809 43129 42843 43163
rect 18199 43061 18233 43095
rect 18613 43061 18647 43095
rect 18889 43061 18923 43095
rect 20085 43061 20119 43095
rect 20959 43061 20993 43095
rect 21649 43061 21683 43095
rect 22937 43061 22971 43095
rect 23995 43061 24029 43095
rect 24409 43061 24443 43095
rect 25973 43061 26007 43095
rect 26893 43061 26927 43095
rect 29101 43061 29135 43095
rect 30297 43061 30331 43095
rect 33333 43061 33367 43095
rect 37565 43061 37599 43095
rect 37841 43061 37875 43095
rect 38485 43061 38519 43095
rect 40233 43061 40267 43095
rect 40647 43061 40681 43095
rect 43407 43061 43441 43095
rect 15531 42857 15565 42891
rect 18981 42857 19015 42891
rect 21051 42857 21085 42891
rect 23995 42857 24029 42891
rect 24777 42857 24811 42891
rect 26893 42857 26927 42891
rect 32321 42857 32355 42891
rect 33057 42857 33091 42891
rect 33609 42857 33643 42891
rect 36829 42857 36863 42891
rect 37887 42857 37921 42891
rect 40785 42857 40819 42891
rect 16589 42789 16623 42823
rect 19257 42789 19291 42823
rect 22017 42789 22051 42823
rect 22109 42789 22143 42823
rect 25053 42789 25087 42823
rect 28825 42789 28859 42823
rect 29377 42789 29411 42823
rect 30526 42789 30560 42823
rect 34805 42789 34839 42823
rect 35725 42789 35759 42823
rect 39583 42789 39617 42823
rect 41061 42789 41095 42823
rect 41153 42789 41187 42823
rect 41705 42789 41739 42823
rect 43545 42789 43579 42823
rect 15460 42721 15494 42755
rect 18112 42721 18146 42755
rect 20948 42721 20982 42755
rect 23857 42721 23891 42755
rect 25605 42721 25639 42755
rect 27077 42721 27111 42755
rect 27353 42721 27387 42755
rect 35357 42721 35391 42755
rect 36185 42721 36219 42755
rect 37816 42721 37850 42755
rect 16497 42653 16531 42687
rect 18199 42653 18233 42687
rect 19165 42653 19199 42687
rect 24961 42653 24995 42687
rect 28733 42653 28767 42687
rect 30205 42653 30239 42687
rect 32689 42653 32723 42687
rect 34529 42653 34563 42687
rect 34713 42653 34747 42687
rect 39221 42653 39255 42687
rect 43453 42653 43487 42687
rect 43729 42653 43763 42687
rect 17049 42585 17083 42619
rect 19717 42585 19751 42619
rect 22569 42585 22603 42619
rect 15945 42517 15979 42551
rect 21741 42517 21775 42551
rect 31125 42517 31159 42551
rect 36415 42517 36449 42551
rect 38485 42517 38519 42551
rect 40141 42517 40175 42551
rect 42349 42517 42383 42551
rect 14703 42313 14737 42347
rect 16497 42313 16531 42347
rect 16773 42313 16807 42347
rect 20729 42313 20763 42347
rect 21373 42313 21407 42347
rect 22937 42313 22971 42347
rect 26525 42313 26559 42347
rect 28319 42313 28353 42347
rect 29101 42313 29135 42347
rect 31953 42313 31987 42347
rect 36277 42313 36311 42347
rect 40233 42313 40267 42347
rect 43453 42313 43487 42347
rect 17141 42245 17175 42279
rect 21051 42245 21085 42279
rect 23305 42245 23339 42279
rect 26065 42245 26099 42279
rect 26341 42245 26375 42279
rect 27629 42245 27663 42279
rect 41889 42245 41923 42279
rect 42901 42245 42935 42279
rect 44465 42245 44499 42279
rect 22017 42177 22051 42211
rect 24179 42177 24213 42211
rect 14632 42109 14666 42143
rect 15577 42109 15611 42143
rect 20980 42109 21014 42143
rect 21741 42109 21775 42143
rect 24092 42109 24126 42143
rect 25789 42109 25823 42143
rect 26709 42177 26743 42211
rect 27997 42177 28031 42211
rect 32689 42177 32723 42211
rect 33425 42177 33459 42211
rect 35633 42177 35667 42211
rect 36001 42177 36035 42211
rect 36553 42177 36587 42211
rect 36829 42177 36863 42211
rect 37841 42177 37875 42211
rect 40785 42177 40819 42211
rect 28248 42109 28282 42143
rect 30573 42109 30607 42143
rect 30849 42109 30883 42143
rect 32045 42109 32079 42143
rect 32505 42109 32539 42143
rect 33660 42109 33694 42143
rect 34621 42109 34655 42143
rect 38209 42109 38243 42143
rect 38669 42109 38703 42143
rect 15485 42041 15519 42075
rect 15939 42041 15973 42075
rect 18337 42041 18371 42075
rect 19165 42041 19199 42075
rect 19441 42041 19475 42075
rect 19533 42041 19567 42075
rect 20085 42041 20119 42075
rect 22109 42041 22143 42075
rect 22661 42041 22695 42075
rect 25145 42041 25179 42075
rect 25237 42041 25271 42075
rect 26341 42041 26375 42075
rect 26801 42041 26835 42075
rect 27353 42041 27387 42075
rect 29837 42041 29871 42075
rect 34989 42041 35023 42075
rect 35081 42041 35115 42075
rect 36645 42041 36679 42075
rect 38577 42041 38611 42075
rect 38990 42041 39024 42075
rect 40877 42041 40911 42075
rect 41429 42041 41463 42075
rect 44833 42177 44867 42211
rect 42349 42041 42383 42075
rect 42441 42041 42475 42075
rect 43913 42041 43947 42075
rect 44005 42041 44039 42075
rect 15025 41973 15059 42007
rect 18889 41973 18923 42007
rect 20361 41973 20395 42007
rect 23857 41973 23891 42007
rect 24593 41973 24627 42007
rect 24961 41973 24995 42007
rect 28733 41973 28767 42007
rect 30205 41973 30239 42007
rect 30573 41973 30607 42007
rect 31585 41973 31619 42007
rect 33057 41973 33091 42007
rect 33747 41973 33781 42007
rect 34161 41973 34195 42007
rect 39589 41973 39623 42007
rect 39957 41973 39991 42007
rect 41705 41973 41739 42007
rect 41889 41973 41923 42007
rect 42073 41973 42107 42007
rect 19533 41769 19567 41803
rect 19809 41769 19843 41803
rect 21281 41769 21315 41803
rect 21833 41769 21867 41803
rect 22109 41769 22143 41803
rect 24685 41769 24719 41803
rect 26985 41769 27019 41803
rect 28825 41769 28859 41803
rect 30757 41769 30791 41803
rect 31125 41769 31159 41803
rect 34897 41769 34931 41803
rect 36553 41769 36587 41803
rect 38209 41769 38243 41803
rect 39221 41769 39255 41803
rect 41061 41769 41095 41803
rect 43499 41769 43533 41803
rect 44189 41769 44223 41803
rect 16681 41701 16715 41735
rect 17233 41701 17267 41735
rect 18975 41701 19009 41735
rect 22477 41701 22511 41735
rect 22845 41701 22879 41735
rect 23397 41701 23431 41735
rect 25053 41701 25087 41735
rect 25605 41701 25639 41735
rect 27997 41701 28031 41735
rect 29561 41701 29595 41735
rect 30481 41701 30515 41735
rect 33977 41701 34011 41735
rect 34069 41701 34103 41735
rect 34621 41701 34655 41735
rect 35633 41701 35667 41735
rect 40186 41701 40220 41735
rect 41889 41701 41923 41735
rect 42441 41701 42475 41735
rect 26433 41633 26467 41667
rect 30941 41633 30975 41667
rect 32908 41633 32942 41667
rect 37933 41633 37967 41667
rect 38393 41633 38427 41667
rect 43269 41633 43303 41667
rect 15623 41565 15657 41599
rect 16589 41565 16623 41599
rect 18613 41565 18647 41599
rect 20913 41565 20947 41599
rect 22753 41565 22787 41599
rect 24961 41565 24995 41599
rect 26663 41565 26697 41599
rect 27905 41565 27939 41599
rect 29469 41565 29503 41599
rect 29745 41565 29779 41599
rect 35541 41565 35575 41599
rect 36001 41565 36035 41599
rect 39865 41565 39899 41599
rect 41797 41565 41831 41599
rect 43821 41565 43855 41599
rect 15393 41497 15427 41531
rect 28457 41497 28491 41531
rect 40785 41497 40819 41531
rect 15945 41429 15979 41463
rect 25881 41429 25915 41463
rect 27537 41429 27571 41463
rect 32689 41429 32723 41463
rect 33011 41429 33045 41463
rect 35265 41429 35299 41463
rect 37381 41429 37415 41463
rect 16313 41225 16347 41259
rect 17417 41225 17451 41259
rect 18705 41225 18739 41259
rect 21925 41225 21959 41259
rect 23029 41225 23063 41259
rect 23995 41225 24029 41259
rect 28365 41225 28399 41259
rect 28641 41225 28675 41259
rect 29561 41225 29595 41259
rect 33609 41225 33643 41259
rect 33885 41225 33919 41259
rect 34253 41225 34287 41259
rect 34621 41225 34655 41259
rect 37197 41225 37231 41259
rect 40785 41225 40819 41259
rect 41107 41225 41141 41259
rect 43085 41225 43119 41259
rect 21005 41157 21039 41191
rect 25789 41157 25823 41191
rect 26065 41157 26099 41191
rect 31309 41157 31343 41191
rect 35449 41157 35483 41191
rect 38393 41157 38427 41191
rect 42625 41157 42659 41191
rect 16497 41089 16531 41123
rect 19901 41089 19935 41123
rect 22569 41089 22603 41123
rect 24685 41089 24719 41123
rect 24869 41089 24903 41123
rect 29009 41089 29043 41123
rect 32229 41089 32263 41123
rect 32689 41089 32723 41123
rect 35817 41089 35851 41123
rect 36093 41089 36127 41123
rect 37381 41089 37415 41123
rect 37657 41089 37691 41123
rect 39589 41089 39623 41123
rect 40233 41089 40267 41123
rect 42073 41089 42107 41123
rect 43361 41089 43395 41123
rect 23924 41021 23958 41055
rect 24317 41021 24351 41055
rect 27445 41021 27479 41055
rect 29929 41021 29963 41055
rect 30389 41021 30423 41055
rect 38853 41021 38887 41055
rect 39313 41021 39347 41055
rect 41004 41021 41038 41055
rect 41429 41021 41463 41055
rect 15945 40953 15979 40987
rect 16589 40953 16623 40987
rect 17141 40953 17175 40987
rect 19717 40953 19751 40987
rect 19970 40953 20004 40987
rect 20545 40953 20579 40987
rect 22109 40953 22143 40987
rect 22201 40953 22235 40987
rect 25190 40953 25224 40987
rect 27261 40953 27295 40987
rect 27766 40953 27800 40987
rect 30297 40953 30331 40987
rect 30751 40953 30785 40987
rect 32597 40953 32631 40987
rect 33051 40953 33085 40987
rect 35909 40953 35943 40987
rect 37473 40953 37507 40987
rect 42165 40953 42199 40987
rect 15485 40885 15519 40919
rect 18981 40885 19015 40919
rect 21281 40885 21315 40919
rect 23397 40885 23431 40919
rect 26525 40885 26559 40919
rect 31585 40885 31619 40919
rect 35173 40885 35207 40919
rect 38669 40885 38703 40919
rect 39865 40885 39899 40919
rect 41797 40885 41831 40919
rect 16405 40681 16439 40715
rect 17141 40681 17175 40715
rect 21327 40681 21361 40715
rect 21741 40681 21775 40715
rect 22109 40681 22143 40715
rect 24409 40681 24443 40715
rect 24777 40681 24811 40715
rect 27905 40681 27939 40715
rect 28641 40681 28675 40715
rect 29193 40681 29227 40715
rect 30573 40681 30607 40715
rect 33839 40681 33873 40715
rect 35633 40681 35667 40715
rect 36001 40681 36035 40715
rect 36599 40681 36633 40715
rect 38945 40681 38979 40715
rect 41613 40681 41647 40715
rect 15847 40613 15881 40647
rect 17417 40613 17451 40647
rect 19901 40613 19935 40647
rect 22385 40613 22419 40647
rect 22937 40613 22971 40647
rect 25053 40613 25087 40647
rect 25605 40613 25639 40647
rect 35034 40613 35068 40647
rect 37289 40613 37323 40647
rect 41889 40613 41923 40647
rect 42441 40613 42475 40647
rect 18981 40545 19015 40579
rect 21256 40545 21290 40579
rect 23816 40545 23850 40579
rect 26985 40545 27019 40579
rect 27261 40545 27295 40579
rect 30573 40545 30607 40579
rect 31033 40545 31067 40579
rect 32137 40545 32171 40579
rect 32597 40545 32631 40579
rect 33768 40545 33802 40579
rect 36461 40545 36495 40579
rect 39129 40545 39163 40579
rect 39589 40545 39623 40579
rect 43428 40545 43462 40579
rect 15485 40477 15519 40511
rect 17325 40477 17359 40511
rect 17969 40477 18003 40511
rect 22293 40477 22327 40511
rect 23903 40477 23937 40511
rect 24961 40477 24995 40511
rect 27445 40477 27479 40511
rect 28273 40477 28307 40511
rect 32689 40477 32723 40511
rect 34713 40477 34747 40511
rect 39865 40477 39899 40511
rect 41797 40477 41831 40511
rect 16681 40341 16715 40375
rect 19165 40341 19199 40375
rect 38025 40341 38059 40375
rect 40509 40341 40543 40375
rect 43499 40341 43533 40375
rect 17049 40137 17083 40171
rect 17417 40137 17451 40171
rect 18613 40137 18647 40171
rect 19993 40137 20027 40171
rect 21557 40137 21591 40171
rect 23029 40137 23063 40171
rect 25605 40137 25639 40171
rect 26433 40137 26467 40171
rect 28549 40137 28583 40171
rect 28917 40137 28951 40171
rect 32229 40137 32263 40171
rect 33057 40137 33091 40171
rect 34253 40137 34287 40171
rect 35173 40137 35207 40171
rect 37749 40137 37783 40171
rect 39589 40137 39623 40171
rect 41429 40137 41463 40171
rect 42165 40137 42199 40171
rect 17693 40069 17727 40103
rect 22661 40069 22695 40103
rect 23857 40069 23891 40103
rect 26985 40069 27019 40103
rect 32505 40069 32539 40103
rect 36277 40069 36311 40103
rect 21143 40001 21177 40035
rect 22109 40001 22143 40035
rect 23397 40001 23431 40035
rect 33977 40001 34011 40035
rect 34621 40001 34655 40035
rect 36737 40001 36771 40035
rect 38577 40001 38611 40035
rect 40233 40001 40267 40035
rect 41797 40001 41831 40035
rect 42809 40001 42843 40035
rect 43085 40001 43119 40035
rect 16129 39933 16163 39967
rect 19073 39933 19107 39967
rect 21051 39933 21085 39967
rect 23673 39933 23707 39967
rect 24501 39933 24535 39967
rect 24844 39933 24878 39967
rect 25973 39933 26007 39967
rect 26576 39933 26610 39967
rect 27537 39933 27571 39967
rect 27997 39933 28031 39967
rect 30941 39933 30975 39967
rect 31401 39933 31435 39967
rect 33241 39933 33275 39967
rect 33701 39933 33735 39967
rect 35408 39933 35442 39967
rect 35817 39933 35851 39967
rect 37933 39933 37967 39967
rect 38393 39933 38427 39967
rect 40509 39933 40543 39967
rect 15577 39865 15611 39899
rect 16037 39865 16071 39899
rect 16491 39865 16525 39899
rect 18981 39865 19015 39899
rect 19435 39865 19469 39899
rect 22201 39865 22235 39899
rect 25053 39865 25087 39899
rect 26663 39865 26697 39899
rect 35495 39865 35529 39899
rect 36461 39865 36495 39899
rect 36553 39865 36587 39899
rect 40760 39865 40794 39899
rect 42901 39865 42935 39899
rect 15209 39797 15243 39831
rect 21925 39797 21959 39831
rect 24225 39797 24259 39831
rect 25329 39797 25363 39831
rect 27445 39797 27479 39831
rect 27629 39797 27663 39831
rect 30205 39797 30239 39831
rect 30573 39797 30607 39831
rect 30941 39797 30975 39831
rect 39129 39797 39163 39831
rect 42533 39797 42567 39831
rect 43821 39797 43855 39831
rect 17141 39593 17175 39627
rect 22385 39593 22419 39627
rect 22753 39593 22787 39627
rect 24961 39593 24995 39627
rect 26709 39593 26743 39627
rect 27721 39593 27755 39627
rect 28641 39593 28675 39627
rect 30941 39593 30975 39627
rect 32229 39593 32263 39627
rect 33241 39593 33275 39627
rect 36553 39593 36587 39627
rect 36829 39593 36863 39627
rect 37933 39593 37967 39627
rect 39129 39593 39163 39627
rect 39681 39593 39715 39627
rect 41429 39593 41463 39627
rect 42809 39593 42843 39627
rect 16542 39525 16576 39559
rect 18061 39525 18095 39559
rect 18153 39525 18187 39559
rect 18705 39525 18739 39559
rect 21827 39525 21861 39559
rect 30573 39525 30607 39559
rect 34022 39525 34056 39559
rect 35633 39525 35667 39559
rect 40785 39525 40819 39559
rect 41797 39525 41831 39559
rect 43545 39525 43579 39559
rect 44097 39525 44131 39559
rect 19533 39457 19567 39491
rect 23213 39457 23247 39491
rect 24225 39457 24259 39491
rect 25304 39457 25338 39491
rect 26893 39457 26927 39491
rect 27077 39457 27111 39491
rect 31033 39457 31067 39491
rect 32137 39457 32171 39491
rect 32597 39457 32631 39491
rect 34621 39457 34655 39491
rect 37749 39457 37783 39491
rect 40509 39457 40543 39491
rect 42257 39457 42291 39491
rect 16221 39389 16255 39423
rect 21465 39389 21499 39423
rect 28273 39389 28307 39423
rect 33701 39389 33735 39423
rect 35541 39389 35575 39423
rect 38761 39389 38795 39423
rect 42395 39389 42429 39423
rect 43453 39389 43487 39423
rect 24409 39321 24443 39355
rect 25789 39321 25823 39355
rect 31217 39321 31251 39355
rect 36093 39321 36127 39355
rect 19073 39253 19107 39287
rect 19671 39253 19705 39287
rect 23351 39253 23385 39287
rect 25375 39253 25409 39287
rect 29193 39253 29227 39287
rect 29469 39253 29503 39287
rect 16221 39049 16255 39083
rect 17509 39049 17543 39083
rect 20361 39049 20395 39083
rect 22615 39049 22649 39083
rect 26709 39049 26743 39083
rect 28641 39049 28675 39083
rect 29101 39049 29135 39083
rect 30389 39049 30423 39083
rect 32137 39049 32171 39083
rect 32873 39049 32907 39083
rect 34621 39049 34655 39083
rect 36645 39049 36679 39083
rect 36921 39049 36955 39083
rect 38301 39049 38335 39083
rect 40233 39049 40267 39083
rect 41061 39049 41095 39083
rect 41429 39049 41463 39083
rect 42993 39049 43027 39083
rect 43453 39049 43487 39083
rect 22017 38981 22051 39015
rect 23305 38981 23339 39015
rect 25145 38981 25179 39015
rect 32505 38981 32539 39015
rect 37289 38981 37323 39015
rect 13921 38913 13955 38947
rect 15301 38913 15335 38947
rect 19073 38913 19107 38947
rect 21649 38913 21683 38947
rect 22293 38913 22327 38947
rect 29377 38913 29411 38947
rect 29653 38913 29687 38947
rect 33701 38913 33735 38947
rect 39589 38913 39623 38947
rect 13093 38845 13127 38879
rect 13461 38845 13495 38879
rect 13737 38845 13771 38879
rect 14657 38845 14691 38879
rect 14749 38845 14783 38879
rect 15209 38845 15243 38879
rect 16313 38845 16347 38879
rect 16865 38845 16899 38879
rect 18337 38845 18371 38879
rect 18429 38845 18463 38879
rect 18981 38845 19015 38879
rect 19625 38845 19659 38879
rect 21189 38845 21223 38879
rect 21373 38845 21407 38879
rect 22544 38845 22578 38879
rect 22937 38845 22971 38879
rect 24292 38845 24326 38879
rect 24685 38845 24719 38879
rect 25237 38845 25271 38879
rect 27537 38845 27571 38879
rect 27905 38845 27939 38879
rect 28181 38845 28215 38879
rect 30849 38845 30883 38879
rect 33057 38845 33091 38879
rect 33517 38845 33551 38879
rect 35265 38845 35299 38879
rect 35725 38845 35759 38879
rect 37508 38845 37542 38879
rect 38853 38845 38887 38879
rect 39313 38845 39347 38879
rect 40668 38845 40702 38879
rect 41680 38845 41714 38879
rect 43888 38845 43922 38879
rect 17877 38777 17911 38811
rect 20821 38777 20855 38811
rect 24133 38777 24167 38811
rect 25558 38777 25592 38811
rect 27077 38777 27111 38811
rect 28365 38777 28399 38811
rect 29469 38777 29503 38811
rect 30757 38777 30791 38811
rect 31211 38777 31245 38811
rect 36046 38777 36080 38811
rect 38669 38777 38703 38811
rect 15761 38709 15795 38743
rect 16589 38709 16623 38743
rect 24363 38709 24397 38743
rect 26157 38709 26191 38743
rect 31769 38709 31803 38743
rect 34069 38709 34103 38743
rect 35541 38709 35575 38743
rect 37611 38709 37645 38743
rect 38025 38709 38059 38743
rect 40739 38709 40773 38743
rect 41751 38709 41785 38743
rect 42349 38709 42383 38743
rect 43959 38709 43993 38743
rect 44373 38709 44407 38743
rect 16497 38505 16531 38539
rect 16773 38505 16807 38539
rect 17969 38505 18003 38539
rect 19533 38505 19567 38539
rect 21189 38505 21223 38539
rect 25973 38505 26007 38539
rect 28273 38505 28307 38539
rect 31861 38505 31895 38539
rect 32505 38505 32539 38539
rect 35265 38505 35299 38539
rect 36829 38505 36863 38539
rect 38853 38505 38887 38539
rect 14841 38437 14875 38471
rect 16129 38437 16163 38471
rect 18889 38437 18923 38471
rect 23350 38437 23384 38471
rect 24961 38437 24995 38471
rect 25053 38437 25087 38471
rect 26709 38437 26743 38471
rect 28870 38437 28904 38471
rect 30665 38437 30699 38471
rect 38485 38437 38519 38471
rect 39221 38437 39255 38471
rect 41797 38437 41831 38471
rect 41889 38437 41923 38471
rect 44097 38437 44131 38471
rect 15669 38369 15703 38403
rect 15945 38369 15979 38403
rect 18153 38369 18187 38403
rect 18705 38369 18739 38403
rect 19876 38369 19910 38403
rect 20913 38369 20947 38403
rect 21373 38369 21407 38403
rect 32137 38369 32171 38403
rect 33977 38369 34011 38403
rect 35265 38369 35299 38403
rect 35449 38369 35483 38403
rect 36645 38369 36679 38403
rect 37749 38369 37783 38403
rect 38301 38369 38335 38403
rect 40636 38369 40670 38403
rect 13277 38301 13311 38335
rect 23029 38301 23063 38335
rect 26617 38301 26651 38335
rect 27261 38301 27295 38335
rect 28549 38301 28583 38335
rect 30573 38301 30607 38335
rect 39497 38301 39531 38335
rect 44005 38301 44039 38335
rect 44649 38301 44683 38335
rect 25513 38233 25547 38267
rect 31125 38233 31159 38267
rect 34161 38233 34195 38267
rect 41429 38233 41463 38267
rect 42349 38233 42383 38267
rect 17049 38165 17083 38199
rect 17279 38165 17313 38199
rect 19947 38165 19981 38199
rect 22845 38165 22879 38199
rect 23949 38165 23983 38199
rect 27721 38165 27755 38199
rect 29469 38165 29503 38199
rect 31493 38165 31527 38199
rect 33057 38165 33091 38199
rect 33701 38165 33735 38199
rect 36001 38165 36035 38199
rect 39727 38165 39761 38199
rect 40739 38165 40773 38199
rect 41061 38165 41095 38199
rect 15761 37961 15795 37995
rect 17877 37961 17911 37995
rect 18613 37961 18647 37995
rect 21373 37961 21407 37995
rect 26617 37961 26651 37995
rect 26985 37961 27019 37995
rect 27445 37961 27479 37995
rect 28733 37961 28767 37995
rect 30389 37961 30423 37995
rect 32137 37961 32171 37995
rect 33609 37961 33643 37995
rect 33977 37961 34011 37995
rect 35081 37961 35115 37995
rect 35541 37961 35575 37995
rect 36553 37961 36587 37995
rect 39037 37961 39071 37995
rect 40325 37961 40359 37995
rect 46581 37961 46615 37995
rect 15485 37893 15519 37927
rect 16589 37893 16623 37927
rect 20913 37893 20947 37927
rect 29929 37893 29963 37927
rect 42993 37893 43027 37927
rect 44741 37893 44775 37927
rect 19625 37825 19659 37859
rect 19901 37825 19935 37859
rect 22753 37825 22787 37859
rect 28273 37825 28307 37859
rect 31493 37825 31527 37859
rect 32965 37825 32999 37859
rect 35633 37825 35667 37859
rect 40877 37825 40911 37859
rect 44189 37825 44223 37859
rect 45109 37825 45143 37859
rect 15000 37757 15034 37791
rect 18128 37757 18162 37791
rect 22017 37757 22051 37791
rect 22477 37757 22511 37791
rect 23673 37757 23707 37791
rect 27629 37757 27663 37791
rect 28181 37757 28215 37791
rect 30757 37757 30791 37791
rect 31125 37757 31159 37791
rect 31401 37757 31435 37791
rect 37933 37757 37967 37791
rect 38301 37757 38335 37791
rect 38485 37757 38519 37791
rect 46156 37757 46190 37791
rect 14841 37689 14875 37723
rect 16037 37689 16071 37723
rect 16129 37689 16163 37723
rect 18889 37689 18923 37723
rect 19717 37689 19751 37723
rect 23994 37689 24028 37723
rect 25697 37689 25731 37723
rect 25789 37689 25823 37723
rect 26341 37689 26375 37723
rect 29377 37689 29411 37723
rect 29469 37689 29503 37723
rect 32689 37689 32723 37723
rect 32781 37689 32815 37723
rect 35954 37689 35988 37723
rect 37473 37689 37507 37723
rect 38761 37689 38795 37723
rect 40969 37689 41003 37723
rect 41521 37689 41555 37723
rect 42441 37689 42475 37723
rect 42533 37689 42567 37723
rect 43637 37689 43671 37723
rect 43913 37689 43947 37723
rect 44281 37689 44315 37723
rect 15071 37621 15105 37655
rect 17233 37621 17267 37655
rect 18199 37621 18233 37655
rect 19441 37621 19475 37655
rect 20545 37621 20579 37655
rect 21833 37621 21867 37655
rect 23029 37621 23063 37655
rect 23397 37621 23431 37655
rect 24593 37621 24627 37655
rect 24961 37621 24995 37655
rect 25513 37621 25547 37655
rect 29101 37621 29135 37655
rect 34713 37621 34747 37655
rect 36921 37621 36955 37655
rect 39681 37621 39715 37655
rect 41797 37621 41831 37655
rect 42165 37621 42199 37655
rect 46259 37621 46293 37655
rect 15577 37417 15611 37451
rect 18705 37417 18739 37451
rect 23765 37417 23799 37451
rect 24961 37417 24995 37451
rect 27721 37417 27755 37451
rect 29193 37417 29227 37451
rect 30941 37417 30975 37451
rect 32781 37417 32815 37451
rect 39221 37417 39255 37451
rect 39773 37417 39807 37451
rect 41797 37417 41831 37451
rect 42441 37417 42475 37451
rect 44005 37417 44039 37451
rect 16037 37349 16071 37383
rect 16129 37349 16163 37383
rect 16957 37349 16991 37383
rect 17785 37349 17819 37383
rect 17877 37349 17911 37383
rect 19441 37349 19475 37383
rect 21097 37349 21131 37383
rect 23489 37349 23523 37383
rect 28365 37349 28399 37383
rect 33701 37349 33735 37383
rect 35817 37349 35851 37383
rect 40922 37349 40956 37383
rect 44465 37349 44499 37383
rect 46029 37349 46063 37383
rect 14232 37281 14266 37315
rect 22753 37281 22787 37315
rect 23213 37281 23247 37315
rect 24368 37281 24402 37315
rect 25329 37281 25363 37315
rect 26592 37281 26626 37315
rect 29837 37281 29871 37315
rect 31033 37281 31067 37315
rect 35357 37281 35391 37315
rect 35541 37281 35575 37315
rect 36645 37281 36679 37315
rect 37749 37281 37783 37315
rect 19349 37213 19383 37247
rect 19625 37213 19659 37247
rect 21005 37213 21039 37247
rect 21373 37213 21407 37247
rect 24455 37213 24489 37247
rect 25789 37213 25823 37247
rect 28273 37213 28307 37247
rect 28549 37213 28583 37247
rect 32229 37213 32263 37247
rect 33609 37213 33643 37247
rect 34253 37213 34287 37247
rect 38853 37213 38887 37247
rect 40601 37213 40635 37247
rect 44373 37213 44407 37247
rect 44741 37213 44775 37247
rect 45937 37213 45971 37247
rect 46213 37213 46247 37247
rect 16589 37145 16623 37179
rect 18337 37145 18371 37179
rect 26663 37145 26697 37179
rect 33149 37145 33183 37179
rect 41521 37145 41555 37179
rect 14335 37077 14369 37111
rect 22017 37077 22051 37111
rect 24133 37077 24167 37111
rect 25467 37077 25501 37111
rect 29561 37077 29595 37111
rect 30067 37077 30101 37111
rect 30481 37077 30515 37111
rect 31217 37077 31251 37111
rect 36829 37077 36863 37111
rect 37105 37077 37139 37111
rect 37979 37077 38013 37111
rect 38393 37077 38427 37111
rect 15485 36873 15519 36907
rect 16037 36873 16071 36907
rect 19717 36873 19751 36907
rect 20177 36873 20211 36907
rect 22339 36873 22373 36907
rect 23397 36873 23431 36907
rect 24685 36873 24719 36907
rect 25329 36873 25363 36907
rect 26801 36873 26835 36907
rect 28365 36873 28399 36907
rect 30665 36873 30699 36907
rect 32229 36873 32263 36907
rect 35173 36873 35207 36907
rect 35817 36873 35851 36907
rect 36645 36873 36679 36907
rect 37749 36873 37783 36907
rect 42579 36873 42613 36907
rect 43361 36873 43395 36907
rect 43591 36873 43625 36907
rect 16957 36805 16991 36839
rect 19441 36805 19475 36839
rect 23029 36805 23063 36839
rect 34713 36805 34747 36839
rect 38025 36805 38059 36839
rect 39589 36805 39623 36839
rect 40141 36805 40175 36839
rect 40325 36805 40359 36839
rect 41521 36805 41555 36839
rect 45845 36805 45879 36839
rect 16405 36737 16439 36771
rect 18429 36737 18463 36771
rect 19073 36737 19107 36771
rect 20729 36737 20763 36771
rect 23765 36737 23799 36771
rect 24225 36737 24259 36771
rect 25881 36737 25915 36771
rect 26249 36737 26283 36771
rect 30021 36737 30055 36771
rect 32413 36737 32447 36771
rect 32689 36737 32723 36771
rect 36829 36737 36863 36771
rect 40969 36737 41003 36771
rect 41889 36737 41923 36771
rect 44373 36737 44407 36771
rect 44557 36737 44591 36771
rect 46121 36737 46155 36771
rect 14565 36669 14599 36703
rect 22268 36669 22302 36703
rect 27972 36669 28006 36703
rect 31360 36669 31394 36703
rect 34989 36669 35023 36703
rect 38577 36669 38611 36703
rect 39037 36669 39071 36703
rect 40141 36669 40175 36703
rect 40693 36669 40727 36703
rect 42508 36669 42542 36703
rect 42901 36669 42935 36703
rect 43520 36669 43554 36703
rect 14473 36601 14507 36635
rect 14886 36601 14920 36635
rect 16497 36601 16531 36635
rect 17509 36601 17543 36635
rect 17877 36601 17911 36635
rect 18521 36601 18555 36635
rect 20545 36601 20579 36635
rect 20821 36601 20855 36635
rect 21373 36601 21407 36635
rect 21741 36601 21775 36635
rect 23857 36601 23891 36635
rect 25973 36601 26007 36635
rect 29745 36601 29779 36635
rect 29837 36601 29871 36635
rect 31447 36601 31481 36635
rect 32505 36601 32539 36635
rect 33885 36601 33919 36635
rect 37150 36601 37184 36635
rect 39313 36601 39347 36635
rect 41061 36601 41095 36635
rect 44649 36601 44683 36635
rect 45201 36601 45235 36635
rect 14013 36533 14047 36567
rect 22661 36533 22695 36567
rect 27721 36533 27755 36567
rect 28043 36533 28077 36567
rect 28825 36533 28859 36567
rect 29561 36533 29595 36567
rect 31033 36533 31067 36567
rect 31769 36533 31803 36567
rect 33517 36533 33551 36567
rect 35541 36533 35575 36567
rect 36277 36533 36311 36567
rect 38393 36533 38427 36567
rect 43913 36533 43947 36567
rect 45477 36533 45511 36567
rect 46581 36533 46615 36567
rect 15117 36329 15151 36363
rect 15485 36329 15519 36363
rect 16037 36329 16071 36363
rect 17785 36329 17819 36363
rect 19579 36329 19613 36363
rect 20729 36329 20763 36363
rect 24041 36329 24075 36363
rect 25881 36329 25915 36363
rect 27721 36329 27755 36363
rect 29745 36329 29779 36363
rect 32413 36329 32447 36363
rect 38945 36329 38979 36363
rect 40601 36329 40635 36363
rect 43775 36329 43809 36363
rect 14381 36261 14415 36295
rect 14657 36261 14691 36295
rect 16497 36261 16531 36295
rect 23213 36261 23247 36295
rect 26617 36261 26651 36295
rect 26709 36261 26743 36295
rect 28549 36261 28583 36295
rect 30297 36261 30331 36295
rect 30389 36261 30423 36295
rect 33793 36261 33827 36295
rect 34345 36261 34379 36295
rect 36829 36261 36863 36295
rect 41061 36261 41095 36295
rect 41153 36261 41187 36295
rect 44557 36261 44591 36295
rect 45017 36261 45051 36295
rect 13645 36193 13679 36227
rect 14197 36193 14231 36227
rect 15336 36193 15370 36227
rect 17877 36193 17911 36227
rect 18429 36193 18463 36227
rect 19508 36193 19542 36227
rect 21741 36193 21775 36227
rect 21925 36193 21959 36227
rect 23765 36193 23799 36227
rect 24628 36193 24662 36227
rect 36369 36193 36403 36227
rect 36645 36193 36679 36227
rect 37749 36193 37783 36227
rect 38209 36193 38243 36227
rect 39129 36193 39163 36227
rect 39589 36193 39623 36227
rect 43637 36193 43671 36227
rect 46397 36193 46431 36227
rect 16405 36125 16439 36159
rect 17049 36125 17083 36159
rect 18521 36125 18555 36159
rect 22201 36125 22235 36159
rect 23121 36125 23155 36159
rect 24731 36125 24765 36159
rect 26893 36125 26927 36159
rect 28457 36125 28491 36159
rect 30573 36125 30607 36159
rect 32505 36125 32539 36159
rect 32735 36125 32769 36159
rect 33701 36125 33735 36159
rect 35909 36125 35943 36159
rect 39865 36125 39899 36159
rect 41521 36125 41555 36159
rect 41981 36125 42015 36159
rect 44925 36125 44959 36159
rect 45201 36125 45235 36159
rect 29009 36057 29043 36091
rect 37933 36057 37967 36091
rect 19257 35989 19291 36023
rect 21281 35989 21315 36023
rect 26157 35989 26191 36023
rect 33057 35989 33091 36023
rect 37105 35989 37139 36023
rect 38577 35989 38611 36023
rect 44281 35989 44315 36023
rect 46535 35989 46569 36023
rect 14657 35785 14691 35819
rect 15669 35785 15703 35819
rect 16405 35785 16439 35819
rect 16681 35785 16715 35819
rect 18613 35785 18647 35819
rect 20269 35785 20303 35819
rect 23121 35785 23155 35819
rect 23489 35785 23523 35819
rect 23811 35785 23845 35819
rect 24593 35785 24627 35819
rect 24915 35785 24949 35819
rect 26893 35785 26927 35819
rect 28457 35785 28491 35819
rect 29423 35785 29457 35819
rect 30297 35785 30331 35819
rect 32045 35785 32079 35819
rect 34437 35785 34471 35819
rect 36645 35785 36679 35819
rect 39865 35785 39899 35819
rect 40325 35785 40359 35819
rect 41337 35785 41371 35819
rect 45201 35785 45235 35819
rect 45661 35785 45695 35819
rect 17877 35717 17911 35751
rect 21097 35717 21131 35751
rect 24225 35717 24259 35751
rect 27537 35717 27571 35751
rect 13093 35649 13127 35683
rect 14289 35649 14323 35683
rect 17095 35649 17129 35683
rect 19257 35649 19291 35683
rect 19901 35649 19935 35683
rect 21281 35649 21315 35683
rect 27721 35649 27755 35683
rect 13277 35581 13311 35615
rect 13645 35581 13679 35615
rect 13921 35581 13955 35615
rect 14749 35581 14783 35615
rect 17008 35581 17042 35615
rect 18220 35581 18254 35615
rect 22293 35581 22327 35615
rect 22937 35581 22971 35615
rect 23740 35581 23774 35615
rect 24812 35581 24846 35615
rect 25237 35581 25271 35615
rect 15070 35513 15104 35547
rect 19073 35513 19107 35547
rect 19349 35513 19383 35547
rect 20729 35513 20763 35547
rect 21373 35513 21407 35547
rect 21925 35513 21959 35547
rect 28733 35717 28767 35751
rect 31033 35717 31067 35751
rect 32689 35717 32723 35751
rect 34069 35717 34103 35751
rect 36001 35717 36035 35751
rect 38669 35717 38703 35751
rect 46397 35717 46431 35751
rect 36829 35649 36863 35683
rect 41705 35649 41739 35683
rect 44925 35649 44959 35683
rect 29352 35581 29386 35615
rect 29745 35581 29779 35615
rect 30665 35581 30699 35615
rect 31125 35581 31159 35615
rect 32873 35581 32907 35615
rect 33793 35581 33827 35615
rect 35725 35581 35759 35615
rect 35817 35581 35851 35615
rect 38853 35581 38887 35615
rect 39313 35581 39347 35615
rect 40544 35581 40578 35615
rect 40969 35581 41003 35615
rect 43244 35581 43278 35615
rect 44005 35581 44039 35615
rect 25881 35513 25915 35547
rect 25973 35513 26007 35547
rect 26525 35513 26559 35547
rect 27813 35513 27847 35547
rect 28365 35513 28399 35547
rect 28457 35513 28491 35547
rect 31446 35513 31480 35547
rect 33194 35513 33228 35547
rect 37150 35513 37184 35547
rect 39589 35513 39623 35547
rect 41797 35513 41831 35547
rect 42349 35513 42383 35547
rect 44281 35513 44315 35547
rect 44373 35513 44407 35547
rect 15945 35445 15979 35479
rect 17509 35445 17543 35479
rect 18291 35445 18325 35479
rect 22937 35445 22971 35479
rect 25697 35445 25731 35479
rect 29009 35445 29043 35479
rect 32321 35445 32355 35479
rect 36369 35445 36403 35479
rect 37749 35445 37783 35479
rect 38393 35445 38427 35479
rect 40647 35445 40681 35479
rect 43315 35445 43349 35479
rect 43729 35445 43763 35479
rect 14749 35241 14783 35275
rect 15485 35241 15519 35275
rect 16221 35241 16255 35275
rect 18889 35241 18923 35275
rect 21005 35241 21039 35275
rect 22569 35241 22603 35275
rect 23121 35241 23155 35275
rect 26709 35241 26743 35275
rect 30297 35241 30331 35275
rect 30757 35241 30791 35275
rect 32413 35241 32447 35275
rect 33333 35241 33367 35275
rect 33885 35241 33919 35275
rect 39221 35241 39255 35275
rect 41521 35241 41555 35275
rect 44465 35241 44499 35275
rect 46627 35241 46661 35275
rect 16497 35173 16531 35207
rect 24133 35173 24167 35207
rect 28457 35173 28491 35207
rect 29009 35173 29043 35207
rect 34713 35173 34747 35207
rect 36829 35173 36863 35207
rect 38346 35173 38380 35207
rect 40922 35173 40956 35207
rect 43545 35173 43579 35207
rect 45109 35173 45143 35207
rect 15301 35105 15335 35139
rect 18521 35105 18555 35139
rect 22201 35105 22235 35139
rect 27261 35105 27295 35139
rect 30757 35105 30791 35139
rect 31033 35105 31067 35139
rect 34897 35105 34931 35139
rect 36093 35105 36127 35139
rect 36645 35105 36679 35139
rect 40601 35105 40635 35139
rect 46556 35105 46590 35139
rect 16405 35037 16439 35071
rect 17049 35037 17083 35071
rect 24041 35037 24075 35071
rect 24317 35037 24351 35071
rect 28365 35037 28399 35071
rect 32965 35037 32999 35071
rect 35265 35037 35299 35071
rect 38025 35037 38059 35071
rect 43453 35037 43487 35071
rect 43729 35037 43763 35071
rect 45017 35037 45051 35071
rect 45385 35037 45419 35071
rect 38945 34969 38979 35003
rect 41797 34969 41831 35003
rect 13277 34901 13311 34935
rect 13645 34901 13679 34935
rect 17877 34901 17911 34935
rect 19441 34901 19475 34935
rect 25605 34901 25639 34935
rect 25881 34901 25915 34935
rect 27399 34901 27433 34935
rect 35541 34901 35575 34935
rect 37197 34901 37231 34935
rect 14657 34697 14691 34731
rect 15761 34697 15795 34731
rect 16497 34697 16531 34731
rect 16773 34697 16807 34731
rect 17877 34697 17911 34731
rect 20637 34697 20671 34731
rect 21925 34697 21959 34731
rect 23029 34697 23063 34731
rect 24133 34697 24167 34731
rect 27813 34697 27847 34731
rect 28135 34697 28169 34731
rect 29837 34697 29871 34731
rect 31217 34697 31251 34731
rect 36093 34697 36127 34731
rect 38117 34697 38151 34731
rect 38485 34697 38519 34731
rect 39865 34697 39899 34731
rect 40325 34697 40359 34731
rect 43545 34697 43579 34731
rect 45385 34697 45419 34731
rect 16037 34629 16071 34663
rect 18613 34629 18647 34663
rect 21373 34629 21407 34663
rect 22293 34629 22327 34663
rect 23489 34629 23523 34663
rect 29423 34629 29457 34663
rect 33333 34629 33367 34663
rect 36921 34629 36955 34663
rect 39589 34629 39623 34663
rect 45017 34629 45051 34663
rect 19257 34561 19291 34595
rect 19901 34561 19935 34595
rect 27261 34561 27295 34595
rect 28457 34561 28491 34595
rect 28825 34561 28859 34595
rect 30205 34561 30239 34595
rect 31769 34561 31803 34595
rect 33057 34561 33091 34595
rect 33701 34561 33735 34595
rect 37841 34561 37875 34595
rect 40693 34561 40727 34595
rect 41889 34561 41923 34595
rect 42809 34561 42843 34595
rect 44097 34561 44131 34595
rect 13553 34493 13587 34527
rect 13829 34493 13863 34527
rect 14013 34493 14047 34527
rect 14841 34493 14875 34527
rect 17008 34493 17042 34527
rect 17417 34493 17451 34527
rect 18061 34493 18095 34527
rect 22636 34493 22670 34527
rect 23581 34493 23615 34527
rect 24501 34493 24535 34527
rect 28064 34493 28098 34527
rect 29352 34493 29386 34527
rect 30348 34493 30382 34527
rect 31344 34493 31378 34527
rect 32137 34493 32171 34527
rect 32321 34493 32355 34527
rect 32781 34493 32815 34527
rect 34345 34493 34379 34527
rect 35633 34493 35667 34527
rect 37105 34493 37139 34527
rect 37657 34493 37691 34527
rect 38669 34493 38703 34527
rect 41613 34493 41647 34527
rect 42257 34493 42291 34527
rect 46156 34493 46190 34527
rect 46581 34493 46615 34527
rect 13185 34425 13219 34459
rect 15162 34425 15196 34459
rect 17095 34425 17129 34459
rect 19349 34425 19383 34459
rect 20269 34425 20303 34459
rect 20821 34425 20855 34459
rect 20913 34425 20947 34459
rect 23811 34425 23845 34459
rect 25605 34425 25639 34459
rect 25697 34425 25731 34459
rect 26249 34425 26283 34459
rect 30435 34425 30469 34459
rect 34713 34425 34747 34459
rect 38990 34425 39024 34459
rect 41014 34425 41048 34459
rect 42533 34425 42567 34459
rect 42625 34425 42659 34459
rect 43913 34425 43947 34459
rect 44189 34425 44223 34459
rect 44741 34425 44775 34459
rect 18291 34357 18325 34391
rect 19073 34357 19107 34391
rect 22707 34357 22741 34391
rect 25329 34357 25363 34391
rect 30757 34357 30791 34391
rect 31447 34357 31481 34391
rect 35265 34357 35299 34391
rect 36553 34357 36587 34391
rect 46259 34357 46293 34391
rect 46949 34357 46983 34391
rect 13369 34153 13403 34187
rect 14841 34153 14875 34187
rect 15577 34153 15611 34187
rect 16405 34153 16439 34187
rect 16957 34153 16991 34187
rect 19257 34153 19291 34187
rect 19533 34153 19567 34187
rect 21051 34153 21085 34187
rect 24041 34153 24075 34187
rect 31493 34153 31527 34187
rect 34805 34153 34839 34187
rect 36737 34153 36771 34187
rect 38025 34153 38059 34187
rect 42533 34153 42567 34187
rect 44649 34153 44683 34187
rect 17693 34085 17727 34119
rect 17969 34085 18003 34119
rect 18521 34085 18555 34119
rect 19947 34085 19981 34119
rect 24777 34085 24811 34119
rect 26709 34085 26743 34119
rect 28273 34085 28307 34119
rect 29837 34085 29871 34119
rect 32873 34085 32907 34119
rect 34989 34085 35023 34119
rect 38853 34085 38887 34119
rect 39129 34085 39163 34119
rect 40693 34085 40727 34119
rect 41061 34085 41095 34119
rect 41153 34085 41187 34119
rect 43177 34085 43211 34119
rect 43821 34085 43855 34119
rect 19860 34017 19894 34051
rect 20948 34017 20982 34051
rect 22753 34017 22787 34051
rect 23213 34017 23247 34051
rect 32229 34017 32263 34051
rect 32597 34017 32631 34051
rect 33977 34017 34011 34051
rect 35725 34017 35759 34051
rect 36553 34017 36587 34051
rect 37013 34017 37047 34051
rect 38117 34017 38151 34051
rect 38577 34017 38611 34051
rect 39865 34017 39899 34051
rect 45604 34017 45638 34051
rect 16037 33949 16071 33983
rect 17877 33949 17911 33983
rect 23305 33949 23339 33983
rect 24685 33949 24719 33983
rect 24961 33949 24995 33983
rect 26617 33949 26651 33983
rect 26893 33949 26927 33983
rect 28181 33949 28215 33983
rect 29561 33949 29595 33983
rect 29745 33949 29779 33983
rect 33885 33949 33919 33983
rect 35357 33949 35391 33983
rect 41521 33949 41555 33983
rect 43729 33949 43763 33983
rect 28733 33881 28767 33915
rect 30297 33881 30331 33915
rect 33517 33881 33551 33915
rect 35265 33881 35299 33915
rect 36001 33881 36035 33915
rect 36369 33881 36403 33915
rect 44281 33881 44315 33915
rect 21465 33813 21499 33847
rect 27537 33813 27571 33847
rect 31125 33813 31159 33847
rect 31861 33813 31895 33847
rect 34161 33813 34195 33847
rect 35154 33813 35188 33847
rect 40095 33813 40129 33847
rect 45707 33813 45741 33847
rect 16313 33609 16347 33643
rect 17509 33609 17543 33643
rect 19809 33609 19843 33643
rect 22753 33609 22787 33643
rect 23213 33609 23247 33643
rect 25421 33609 25455 33643
rect 25743 33609 25777 33643
rect 28181 33609 28215 33643
rect 31309 33609 31343 33643
rect 31907 33609 31941 33643
rect 32045 33609 32079 33643
rect 35173 33609 35207 33643
rect 35541 33609 35575 33643
rect 36599 33609 36633 33643
rect 36737 33609 36771 33643
rect 36921 33609 36955 33643
rect 38485 33609 38519 33643
rect 39957 33609 39991 33643
rect 42625 33609 42659 33643
rect 43729 33609 43763 33643
rect 44097 33609 44131 33643
rect 45017 33609 45051 33643
rect 45569 33609 45603 33643
rect 15117 33541 15151 33575
rect 30665 33541 30699 33575
rect 32229 33541 32263 33575
rect 35062 33541 35096 33575
rect 37473 33541 37507 33575
rect 37933 33541 37967 33575
rect 41245 33541 41279 33575
rect 41521 33541 41555 33575
rect 16037 33473 16071 33507
rect 16681 33473 16715 33507
rect 19441 33473 19475 33507
rect 24133 33473 24167 33507
rect 24777 33473 24811 33507
rect 26801 33473 26835 33507
rect 32137 33473 32171 33507
rect 35265 33473 35299 33507
rect 36001 33473 36035 33507
rect 36369 33473 36403 33507
rect 36829 33473 36863 33507
rect 40233 33473 40267 33507
rect 14340 33405 14374 33439
rect 14427 33405 14461 33439
rect 15577 33405 15611 33439
rect 15761 33405 15795 33439
rect 17024 33405 17058 33439
rect 18613 33405 18647 33439
rect 18797 33405 18831 33439
rect 21281 33405 21315 33439
rect 21741 33405 21775 33439
rect 21925 33405 21959 33439
rect 25672 33405 25706 33439
rect 26065 33405 26099 33439
rect 29101 33405 29135 33439
rect 29745 33405 29779 33439
rect 32781 33405 32815 33439
rect 33609 33405 33643 33439
rect 34253 33405 34287 33439
rect 38025 33405 38059 33439
rect 38853 33405 38887 33439
rect 39456 33405 39490 33439
rect 40760 33405 40794 33439
rect 41864 33405 41898 33439
rect 42876 33405 42910 33439
rect 43269 33405 43303 33439
rect 44532 33405 44566 33439
rect 14841 33337 14875 33371
rect 17785 33337 17819 33371
rect 19073 33337 19107 33371
rect 19993 33337 20027 33371
rect 20085 33337 20119 33371
rect 20637 33337 20671 33371
rect 23949 33337 23983 33371
rect 24225 33337 24259 33371
rect 26525 33337 26559 33371
rect 26893 33337 26927 33371
rect 27445 33337 27479 33371
rect 29653 33337 29687 33371
rect 30107 33337 30141 33371
rect 31677 33337 31711 33371
rect 31769 33337 31803 33371
rect 33333 33337 33367 33371
rect 33425 33337 33459 33371
rect 33977 33337 34011 33371
rect 34621 33337 34655 33371
rect 34897 33337 34931 33371
rect 36461 33337 36495 33371
rect 39543 33337 39577 33371
rect 42349 33337 42383 33371
rect 17095 33269 17129 33303
rect 20913 33269 20947 33303
rect 21741 33269 21775 33303
rect 25145 33269 25179 33303
rect 27721 33269 27755 33303
rect 28457 33269 28491 33303
rect 38209 33269 38243 33303
rect 40831 33269 40865 33303
rect 41935 33269 41969 33303
rect 42947 33269 42981 33303
rect 44603 33269 44637 33303
rect 17969 33065 18003 33099
rect 23581 33065 23615 33099
rect 24133 33065 24167 33099
rect 26341 33065 26375 33099
rect 29653 33065 29687 33099
rect 30113 33065 30147 33099
rect 35173 33065 35207 33099
rect 36461 33065 36495 33099
rect 36829 33065 36863 33099
rect 15393 32997 15427 33031
rect 15485 32997 15519 33031
rect 19349 32997 19383 33031
rect 21097 32997 21131 33031
rect 26709 32997 26743 33031
rect 28641 32997 28675 33031
rect 32137 32997 32171 33031
rect 13645 32929 13679 32963
rect 14105 32929 14139 32963
rect 17049 32929 17083 32963
rect 17325 32929 17359 32963
rect 19993 32929 20027 32963
rect 23213 32929 23247 32963
rect 25456 32929 25490 32963
rect 30297 32929 30331 32963
rect 30573 32929 30607 32963
rect 33885 32929 33919 32963
rect 34253 32929 34287 32963
rect 34989 32929 35023 32963
rect 14381 32861 14415 32895
rect 15853 32861 15887 32895
rect 17601 32861 17635 32895
rect 18705 32861 18739 32895
rect 19073 32861 19107 32895
rect 21005 32861 21039 32895
rect 26617 32861 26651 32895
rect 27261 32861 27295 32895
rect 28549 32861 28583 32895
rect 32505 32861 32539 32895
rect 32597 32861 32631 32895
rect 21557 32793 21591 32827
rect 29101 32793 29135 32827
rect 31217 32793 31251 32827
rect 31585 32793 31619 32827
rect 32275 32793 32309 32827
rect 41061 32997 41095 33031
rect 44833 32997 44867 33031
rect 35265 32929 35299 32963
rect 37749 32929 37783 32963
rect 38209 32929 38243 32963
rect 39900 32929 39934 32963
rect 43704 32929 43738 32963
rect 46248 32929 46282 32963
rect 35633 32861 35667 32895
rect 38301 32861 38335 32895
rect 40003 32861 40037 32895
rect 40969 32861 41003 32895
rect 41613 32861 41647 32895
rect 44741 32861 44775 32895
rect 45017 32861 45051 32895
rect 35403 32793 35437 32827
rect 37197 32793 37231 32827
rect 18429 32725 18463 32759
rect 20269 32725 20303 32759
rect 25559 32725 25593 32759
rect 27537 32725 27571 32759
rect 31953 32725 31987 32759
rect 32413 32725 32447 32759
rect 33517 32725 33551 32759
rect 33793 32725 33827 32759
rect 35173 32725 35207 32759
rect 35541 32725 35575 32759
rect 35909 32725 35943 32759
rect 38761 32725 38795 32759
rect 43775 32725 43809 32759
rect 44373 32725 44407 32759
rect 46351 32725 46385 32759
rect 13507 32521 13541 32555
rect 13921 32521 13955 32555
rect 14289 32521 14323 32555
rect 15945 32521 15979 32555
rect 16865 32521 16899 32555
rect 17417 32521 17451 32555
rect 19625 32521 19659 32555
rect 22661 32521 22695 32555
rect 23857 32521 23891 32555
rect 24317 32521 24351 32555
rect 26157 32521 26191 32555
rect 26479 32521 26513 32555
rect 27169 32521 27203 32555
rect 31769 32521 31803 32555
rect 32505 32521 32539 32555
rect 33333 32521 33367 32555
rect 34713 32521 34747 32555
rect 35173 32521 35207 32555
rect 35541 32521 35575 32555
rect 37473 32521 37507 32555
rect 39221 32521 39255 32555
rect 40325 32521 40359 32555
rect 40969 32521 41003 32555
rect 41889 32521 41923 32555
rect 15301 32453 15335 32487
rect 15577 32453 15611 32487
rect 17785 32453 17819 32487
rect 25421 32453 25455 32487
rect 30205 32453 30239 32487
rect 31999 32453 32033 32487
rect 32137 32453 32171 32487
rect 32965 32453 32999 32487
rect 34345 32453 34379 32487
rect 35909 32453 35943 32487
rect 38945 32453 38979 32487
rect 12909 32385 12943 32419
rect 14381 32385 14415 32419
rect 18061 32385 18095 32419
rect 24501 32385 24535 32419
rect 24777 32385 24811 32419
rect 32229 32385 32263 32419
rect 33885 32385 33919 32419
rect 35265 32385 35299 32419
rect 37197 32385 37231 32419
rect 38025 32385 38059 32419
rect 41153 32385 41187 32419
rect 43637 32521 43671 32555
rect 44189 32453 44223 32487
rect 42073 32385 42107 32419
rect 43545 32385 43579 32419
rect 43637 32385 43671 32419
rect 44465 32385 44499 32419
rect 46213 32385 46247 32419
rect 47133 32385 47167 32419
rect 13436 32317 13470 32351
rect 16957 32317 16991 32351
rect 20152 32317 20186 32351
rect 20545 32317 20579 32351
rect 21097 32317 21131 32351
rect 26408 32317 26442 32351
rect 29285 32317 29319 32351
rect 31861 32317 31895 32351
rect 33609 32317 33643 32351
rect 35044 32317 35078 32351
rect 36461 32317 36495 32351
rect 37013 32317 37047 32351
rect 41797 32317 41831 32351
rect 41889 32317 41923 32351
rect 45109 32317 45143 32351
rect 14702 32249 14736 32283
rect 18382 32249 18416 32283
rect 19257 32249 19291 32283
rect 20913 32249 20947 32283
rect 21418 32249 21452 32283
rect 23213 32249 23247 32283
rect 24593 32249 24627 32283
rect 27445 32249 27479 32283
rect 27537 32249 27571 32283
rect 28089 32249 28123 32283
rect 29101 32249 29135 32283
rect 29647 32249 29681 32283
rect 33425 32249 33459 32283
rect 34897 32249 34931 32283
rect 36277 32249 36311 32283
rect 37841 32249 37875 32283
rect 38387 32249 38421 32283
rect 41245 32249 41279 32283
rect 42901 32249 42935 32283
rect 42993 32249 43027 32283
rect 44557 32249 44591 32283
rect 46305 32249 46339 32283
rect 46857 32249 46891 32283
rect 13277 32181 13311 32215
rect 16405 32181 16439 32215
rect 17141 32181 17175 32215
rect 18981 32181 19015 32215
rect 20223 32181 20257 32215
rect 22017 32181 22051 32215
rect 22293 32181 22327 32215
rect 26893 32181 26927 32215
rect 28549 32181 28583 32215
rect 30665 32181 30699 32215
rect 31033 32181 31067 32215
rect 31401 32181 31435 32215
rect 39865 32181 39899 32215
rect 42625 32181 42659 32215
rect 43821 32181 43855 32215
rect 45385 32181 45419 32215
rect 45845 32181 45879 32215
rect 14657 31977 14691 32011
rect 19671 31977 19705 32011
rect 21925 31977 21959 32011
rect 27721 31977 27755 32011
rect 28733 31977 28767 32011
rect 29285 31977 29319 32011
rect 30573 31977 30607 32011
rect 31861 31977 31895 32011
rect 33241 31977 33275 32011
rect 34437 31977 34471 32011
rect 35909 31977 35943 32011
rect 37289 31977 37323 32011
rect 40693 31977 40727 32011
rect 41061 31977 41095 32011
rect 42901 31977 42935 32011
rect 44741 31977 44775 32011
rect 46673 31977 46707 32011
rect 13829 31909 13863 31943
rect 15485 31909 15519 31943
rect 18061 31909 18095 31943
rect 21097 31909 21131 31943
rect 21649 31909 21683 31943
rect 25053 31909 25087 31943
rect 27261 31909 27295 31943
rect 28365 31909 28399 31943
rect 30895 31909 30929 31943
rect 32137 31909 32171 31943
rect 33701 31909 33735 31943
rect 36921 31909 36955 31943
rect 38387 31909 38421 31943
rect 40094 31909 40128 31943
rect 41613 31909 41647 31943
rect 41705 31909 41739 31943
rect 43545 31909 43579 31943
rect 44097 31909 44131 31943
rect 45109 31909 45143 31943
rect 46121 31909 46155 31943
rect 16865 31841 16899 31875
rect 19600 31841 19634 31875
rect 23029 31841 23063 31875
rect 23213 31841 23247 31875
rect 29193 31841 29227 31875
rect 29745 31841 29779 31875
rect 30757 31841 30791 31875
rect 34989 31841 35023 31875
rect 36461 31841 36495 31875
rect 38025 31841 38059 31875
rect 46397 31841 46431 31875
rect 13737 31773 13771 31807
rect 14381 31773 14415 31807
rect 15393 31773 15427 31807
rect 17003 31773 17037 31807
rect 17969 31773 18003 31807
rect 18245 31773 18279 31807
rect 21005 31773 21039 31807
rect 23305 31773 23339 31807
rect 24961 31773 24995 31807
rect 25605 31773 25639 31807
rect 32284 31773 32318 31807
rect 32505 31773 32539 31807
rect 35265 31773 35299 31807
rect 39773 31773 39807 31807
rect 41889 31773 41923 31807
rect 43453 31773 43487 31807
rect 45017 31773 45051 31807
rect 15117 31705 15151 31739
rect 15945 31705 15979 31739
rect 31585 31705 31619 31739
rect 32597 31705 32631 31739
rect 36645 31705 36679 31739
rect 38945 31705 38979 31739
rect 45569 31705 45603 31739
rect 16313 31637 16347 31671
rect 24409 31637 24443 31671
rect 29101 31637 29135 31671
rect 30297 31637 30331 31671
rect 32413 31637 32447 31671
rect 35541 31637 35575 31671
rect 36369 31637 36403 31671
rect 13461 31433 13495 31467
rect 13691 31433 13725 31467
rect 14703 31433 14737 31467
rect 15485 31433 15519 31467
rect 17509 31433 17543 31467
rect 17877 31433 17911 31467
rect 20085 31433 20119 31467
rect 20177 31433 20211 31467
rect 21741 31433 21775 31467
rect 22707 31433 22741 31467
rect 25513 31433 25547 31467
rect 27859 31433 27893 31467
rect 31493 31433 31527 31467
rect 34621 31433 34655 31467
rect 35081 31433 35115 31467
rect 35725 31433 35759 31467
rect 36277 31433 36311 31467
rect 39405 31433 39439 31467
rect 40969 31433 41003 31467
rect 42073 31433 42107 31467
rect 42533 31433 42567 31467
rect 45385 31433 45419 31467
rect 45845 31433 45879 31467
rect 14473 31365 14507 31399
rect 16957 31365 16991 31399
rect 15117 31297 15151 31331
rect 15669 31297 15703 31331
rect 18153 31297 18187 31331
rect 19073 31297 19107 31331
rect 13620 31229 13654 31263
rect 14632 31229 14666 31263
rect 18797 31229 18831 31263
rect 15761 31161 15795 31195
rect 16313 31161 16347 31195
rect 18245 31161 18279 31195
rect 24041 31365 24075 31399
rect 27997 31365 28031 31399
rect 28273 31365 28307 31399
rect 31861 31365 31895 31399
rect 42809 31365 42843 31399
rect 22477 31297 22511 31331
rect 24869 31297 24903 31331
rect 29009 31297 29043 31331
rect 31953 31297 31987 31331
rect 39129 31297 39163 31331
rect 40141 31297 40175 31331
rect 41153 31297 41187 31331
rect 22604 31229 22638 31263
rect 23489 31229 23523 31263
rect 27788 31229 27822 31263
rect 27997 31229 28031 31263
rect 29285 31229 29319 31263
rect 29745 31229 29779 31263
rect 31732 31229 31766 31263
rect 33149 31229 33183 31263
rect 33885 31229 33919 31263
rect 34897 31229 34931 31263
rect 36737 31229 36771 31263
rect 37105 31229 37139 31263
rect 37381 31229 37415 31263
rect 38393 31229 38427 31263
rect 38853 31229 38887 31263
rect 44624 31229 44658 31263
rect 45017 31229 45051 31263
rect 46121 31229 46155 31263
rect 46581 31229 46615 31263
rect 20453 31161 20487 31195
rect 20545 31161 20579 31195
rect 21097 31161 21131 31195
rect 23121 31161 23155 31195
rect 24593 31161 24627 31195
rect 24694 31161 24728 31195
rect 25973 31161 26007 31195
rect 26249 31161 26283 31195
rect 26341 31161 26375 31195
rect 26893 31161 26927 31195
rect 31585 31161 31619 31195
rect 33977 31161 34011 31195
rect 37565 31161 37599 31195
rect 41245 31161 41279 31195
rect 41797 31161 41831 31195
rect 43085 31161 43119 31195
rect 43177 31161 43211 31195
rect 43729 31161 43763 31195
rect 46949 31161 46983 31195
rect 14105 31093 14139 31127
rect 19625 31093 19659 31127
rect 20085 31093 20119 31127
rect 21373 31093 21407 31127
rect 24409 31093 24443 31127
rect 28641 31093 28675 31127
rect 29377 31093 29411 31127
rect 30481 31093 30515 31127
rect 30849 31093 30883 31127
rect 32229 31093 32263 31127
rect 32597 31093 32631 31127
rect 35357 31093 35391 31127
rect 38117 31093 38151 31127
rect 39773 31093 39807 31127
rect 44005 31093 44039 31127
rect 44695 31093 44729 31127
rect 46305 31093 46339 31127
rect 15117 30889 15151 30923
rect 16221 30889 16255 30923
rect 17693 30889 17727 30923
rect 23121 30889 23155 30923
rect 23581 30889 23615 30923
rect 24593 30889 24627 30923
rect 25099 30889 25133 30923
rect 30021 30889 30055 30923
rect 31217 30889 31251 30923
rect 31677 30889 31711 30923
rect 34069 30889 34103 30923
rect 35909 30889 35943 30923
rect 41153 30889 41187 30923
rect 42349 30889 42383 30923
rect 43085 30889 43119 30923
rect 43499 30889 43533 30923
rect 15622 30821 15656 30855
rect 18061 30821 18095 30855
rect 21097 30821 21131 30855
rect 26709 30821 26743 30855
rect 27261 30821 27295 30855
rect 29193 30821 29227 30855
rect 32137 30821 32171 30855
rect 33701 30821 33735 30855
rect 41521 30821 41555 30855
rect 44557 30821 44591 30855
rect 45109 30821 45143 30855
rect 12633 30753 12667 30787
rect 13645 30753 13679 30787
rect 14105 30753 14139 30787
rect 19860 30753 19894 30787
rect 23213 30753 23247 30787
rect 24961 30753 24995 30787
rect 31033 30753 31067 30787
rect 32284 30753 32318 30787
rect 34529 30753 34563 30787
rect 34676 30753 34710 30787
rect 36093 30753 36127 30787
rect 37749 30753 37783 30787
rect 39221 30753 39255 30787
rect 39497 30753 39531 30787
rect 43396 30753 43430 30787
rect 45937 30753 45971 30787
rect 14381 30685 14415 30719
rect 15301 30685 15335 30719
rect 17969 30685 18003 30719
rect 19947 30685 19981 30719
rect 21005 30685 21039 30719
rect 21281 30685 21315 30719
rect 26617 30685 26651 30719
rect 28917 30685 28951 30719
rect 29101 30685 29135 30719
rect 30941 30685 30975 30719
rect 32505 30685 32539 30719
rect 34897 30685 34931 30719
rect 38853 30685 38887 30719
rect 39681 30685 39715 30719
rect 41429 30685 41463 30719
rect 42073 30685 42107 30719
rect 44465 30685 44499 30719
rect 46075 30685 46109 30719
rect 12771 30617 12805 30651
rect 18521 30617 18555 30651
rect 29653 30617 29687 30651
rect 32597 30617 32631 30651
rect 34805 30617 34839 30651
rect 36921 30617 36955 30651
rect 37933 30617 37967 30651
rect 20361 30549 20395 30583
rect 24133 30549 24167 30583
rect 26249 30549 26283 30583
rect 32413 30549 32447 30583
rect 33333 30549 33367 30583
rect 34989 30549 35023 30583
rect 35633 30549 35667 30583
rect 36277 30549 36311 30583
rect 38393 30549 38427 30583
rect 40509 30549 40543 30583
rect 46765 30549 46799 30583
rect 13369 30345 13403 30379
rect 15301 30345 15335 30379
rect 16589 30345 16623 30379
rect 17509 30345 17543 30379
rect 19073 30345 19107 30379
rect 20177 30345 20211 30379
rect 21649 30345 21683 30379
rect 22385 30345 22419 30379
rect 23213 30345 23247 30379
rect 24593 30345 24627 30379
rect 25697 30345 25731 30379
rect 27445 30345 27479 30379
rect 28135 30345 28169 30379
rect 30665 30345 30699 30379
rect 31401 30345 31435 30379
rect 31769 30345 31803 30379
rect 33701 30345 33735 30379
rect 34529 30345 34563 30379
rect 35081 30345 35115 30379
rect 36277 30345 36311 30379
rect 37473 30345 37507 30379
rect 37749 30345 37783 30379
rect 38025 30345 38059 30379
rect 38485 30345 38519 30379
rect 42073 30345 42107 30379
rect 43729 30345 43763 30379
rect 45477 30345 45511 30379
rect 47593 30345 47627 30379
rect 13691 30277 13725 30311
rect 20361 30277 20395 30311
rect 21281 30277 21315 30311
rect 31631 30277 31665 30311
rect 33149 30277 33183 30311
rect 33517 30277 33551 30311
rect 35357 30277 35391 30311
rect 35725 30277 35759 30311
rect 46305 30277 46339 30311
rect 14703 30209 14737 30243
rect 13620 30141 13654 30175
rect 14600 30141 14634 30175
rect 19692 30141 19726 30175
rect 20729 30209 20763 30243
rect 22017 30209 22051 30243
rect 29285 30209 29319 30243
rect 31861 30209 31895 30243
rect 33609 30209 33643 30243
rect 34713 30209 34747 30243
rect 36369 30209 36403 30243
rect 41705 30209 41739 30243
rect 42809 30209 42843 30243
rect 43085 30209 43119 30243
rect 45017 30209 45051 30243
rect 22201 30141 22235 30175
rect 22753 30141 22787 30175
rect 23673 30141 23707 30175
rect 26249 30141 26283 30175
rect 28064 30141 28098 30175
rect 30205 30141 30239 30175
rect 31033 30141 31067 30175
rect 33388 30141 33422 30175
rect 36148 30141 36182 30175
rect 37565 30141 37599 30175
rect 38577 30141 38611 30175
rect 39129 30141 39163 30175
rect 40509 30141 40543 30175
rect 46673 30141 46707 30175
rect 46857 30141 46891 30175
rect 15669 30073 15703 30107
rect 15761 30073 15795 30107
rect 16313 30073 16347 30107
rect 18153 30073 18187 30107
rect 18245 30073 18279 30107
rect 18797 30073 18831 30107
rect 20361 30073 20395 30107
rect 20821 30073 20855 30107
rect 24035 30073 24069 30107
rect 26157 30073 26191 30107
rect 26611 30073 26645 30107
rect 28549 30073 28583 30107
rect 29606 30073 29640 30107
rect 31493 30073 31527 30107
rect 33241 30073 33275 30107
rect 36001 30073 36035 30107
rect 39313 30073 39347 30107
rect 40830 30073 40864 30107
rect 42901 30073 42935 30107
rect 44373 30073 44407 30107
rect 44557 30073 44591 30107
rect 44649 30073 44683 30107
rect 12725 30005 12759 30039
rect 13093 30005 13127 30039
rect 14105 30005 14139 30039
rect 14473 30005 14507 30039
rect 16957 30005 16991 30039
rect 17785 30005 17819 30039
rect 19763 30005 19797 30039
rect 20453 30005 20487 30039
rect 24961 30005 24995 30039
rect 27169 30005 27203 30039
rect 29009 30005 29043 30039
rect 32137 30005 32171 30039
rect 32597 30005 32631 30039
rect 36645 30005 36679 30039
rect 37105 30005 37139 30039
rect 39589 30005 39623 30039
rect 40233 30005 40267 30039
rect 41429 30005 41463 30039
rect 42625 30005 42659 30039
rect 46949 30005 46983 30039
rect 15025 29801 15059 29835
rect 16221 29801 16255 29835
rect 17233 29801 17267 29835
rect 18061 29801 18095 29835
rect 20361 29801 20395 29835
rect 23765 29801 23799 29835
rect 28825 29801 28859 29835
rect 30021 29801 30055 29835
rect 30849 29801 30883 29835
rect 31217 29801 31251 29835
rect 31585 29801 31619 29835
rect 32321 29801 32355 29835
rect 34529 29801 34563 29835
rect 35817 29801 35851 29835
rect 36185 29801 36219 29835
rect 36461 29801 36495 29835
rect 36829 29801 36863 29835
rect 38761 29801 38795 29835
rect 39313 29801 39347 29835
rect 40601 29801 40635 29835
rect 42441 29801 42475 29835
rect 43729 29801 43763 29835
rect 44281 29801 44315 29835
rect 44649 29801 44683 29835
rect 44925 29801 44959 29835
rect 15622 29733 15656 29767
rect 18429 29733 18463 29767
rect 20729 29733 20763 29767
rect 21097 29733 21131 29767
rect 23397 29733 23431 29767
rect 24041 29733 24075 29767
rect 24409 29733 24443 29767
rect 26893 29733 26927 29767
rect 29653 29733 29687 29767
rect 30573 29733 30607 29767
rect 34161 29733 34195 29767
rect 37473 29733 37507 29767
rect 41883 29733 41917 29767
rect 45293 29733 45327 29767
rect 13829 29665 13863 29699
rect 14105 29665 14139 29699
rect 19809 29665 19843 29699
rect 22937 29665 22971 29699
rect 23213 29665 23247 29699
rect 31033 29665 31067 29699
rect 31953 29665 31987 29699
rect 33204 29665 33238 29699
rect 34621 29665 34655 29699
rect 36645 29665 36679 29699
rect 40141 29665 40175 29699
rect 41521 29665 41555 29699
rect 42809 29665 42843 29699
rect 43361 29665 43395 29699
rect 46949 29665 46983 29699
rect 47317 29665 47351 29699
rect 14381 29597 14415 29631
rect 15301 29597 15335 29631
rect 18337 29597 18371 29631
rect 21005 29597 21039 29631
rect 21281 29597 21315 29631
rect 24317 29597 24351 29631
rect 26801 29597 26835 29631
rect 28457 29597 28491 29631
rect 33425 29597 33459 29631
rect 34989 29597 35023 29631
rect 38393 29597 38427 29631
rect 45201 29597 45235 29631
rect 45569 29597 45603 29631
rect 18889 29529 18923 29563
rect 24869 29529 24903 29563
rect 27353 29529 27387 29563
rect 33517 29529 33551 29563
rect 35081 29529 35115 29563
rect 40325 29529 40359 29563
rect 19947 29461 19981 29495
rect 26341 29461 26375 29495
rect 29377 29461 29411 29495
rect 32965 29461 32999 29495
rect 33333 29461 33367 29495
rect 34759 29461 34793 29495
rect 34897 29461 34931 29495
rect 37197 29461 37231 29495
rect 38025 29461 38059 29495
rect 39589 29461 39623 29495
rect 46857 29461 46891 29495
rect 13185 29257 13219 29291
rect 14749 29257 14783 29291
rect 16037 29257 16071 29291
rect 17785 29257 17819 29291
rect 18981 29257 19015 29291
rect 20177 29257 20211 29291
rect 20637 29257 20671 29291
rect 21741 29257 21775 29291
rect 22477 29257 22511 29291
rect 24317 29257 24351 29291
rect 24685 29257 24719 29291
rect 25053 29257 25087 29291
rect 26893 29257 26927 29291
rect 28365 29257 28399 29291
rect 29101 29257 29135 29291
rect 36277 29257 36311 29291
rect 37473 29257 37507 29291
rect 43729 29257 43763 29291
rect 44373 29257 44407 29291
rect 45477 29257 45511 29291
rect 47041 29257 47075 29291
rect 17141 29189 17175 29223
rect 19257 29189 19291 29223
rect 21373 29189 21407 29223
rect 33517 29189 33551 29223
rect 35173 29189 35207 29223
rect 39865 29189 39899 29223
rect 41889 29189 41923 29223
rect 46673 29189 46707 29223
rect 14841 29121 14875 29155
rect 20821 29121 20855 29155
rect 26341 29121 26375 29155
rect 27169 29121 27203 29155
rect 29653 29121 29687 29155
rect 33149 29121 33183 29155
rect 33609 29121 33643 29155
rect 34713 29121 34747 29155
rect 35909 29121 35943 29155
rect 36148 29121 36182 29155
rect 36369 29121 36403 29155
rect 37013 29121 37047 29155
rect 40509 29121 40543 29155
rect 13369 29053 13403 29087
rect 13829 29053 13863 29087
rect 14013 29053 14047 29087
rect 16957 29053 16991 29087
rect 18061 29053 18095 29087
rect 22569 29053 22603 29087
rect 23924 29053 23958 29087
rect 25789 29053 25823 29087
rect 26249 29053 26283 29087
rect 28181 29053 28215 29087
rect 31493 29053 31527 29087
rect 31677 29053 31711 29087
rect 32781 29053 32815 29087
rect 33388 29053 33422 29087
rect 34989 29053 35023 29087
rect 37657 29053 37691 29087
rect 38209 29053 38243 29087
rect 38393 29053 38427 29087
rect 39221 29053 39255 29087
rect 41429 29053 41463 29087
rect 18382 28985 18416 29019
rect 19901 28985 19935 29019
rect 20913 28985 20947 29019
rect 23029 28985 23063 29019
rect 29377 28985 29411 29019
rect 29469 28985 29503 29019
rect 30757 28985 30791 29019
rect 31125 28985 31159 29019
rect 32413 28985 32447 29019
rect 33241 28985 33275 29019
rect 35541 28985 35575 29019
rect 36001 28985 36035 29019
rect 36737 28985 36771 29019
rect 39037 28985 39071 29019
rect 40871 28985 40905 29019
rect 42349 29121 42383 29155
rect 42993 29121 43027 29155
rect 44557 29121 44591 29155
rect 44925 29121 44959 29155
rect 42073 29053 42107 29087
rect 45937 29053 45971 29087
rect 47225 29053 47259 29087
rect 42441 28985 42475 29019
rect 44649 28985 44683 29019
rect 14381 28917 14415 28951
rect 15209 28917 15243 28951
rect 15761 28917 15795 28951
rect 17509 28917 17543 28951
rect 22753 28917 22787 28951
rect 23489 28917 23523 28951
rect 23995 28917 24029 28951
rect 25697 28917 25731 28951
rect 28089 28917 28123 28951
rect 28733 28917 28767 28951
rect 31493 28917 31527 28951
rect 33885 28917 33919 28951
rect 34253 28917 34287 28951
rect 38761 28917 38795 28951
rect 39405 28917 39439 28951
rect 40233 28917 40267 28951
rect 41705 28917 41739 28951
rect 41889 28917 41923 28951
rect 43361 28917 43395 28951
rect 13277 28713 13311 28747
rect 13645 28713 13679 28747
rect 14841 28713 14875 28747
rect 15485 28713 15519 28747
rect 18429 28713 18463 28747
rect 19165 28713 19199 28747
rect 21373 28713 21407 28747
rect 25881 28713 25915 28747
rect 26663 28713 26697 28747
rect 28273 28713 28307 28747
rect 29377 28713 29411 28747
rect 30205 28713 30239 28747
rect 32229 28713 32263 28747
rect 33333 28713 33367 28747
rect 34253 28713 34287 28747
rect 35357 28713 35391 28747
rect 36645 28713 36679 28747
rect 37933 28713 37967 28747
rect 38761 28713 38795 28747
rect 41521 28713 41555 28747
rect 42625 28713 42659 28747
rect 44557 28713 44591 28747
rect 45017 28713 45051 28747
rect 15945 28645 15979 28679
rect 18061 28645 18095 28679
rect 18705 28645 18739 28679
rect 24863 28645 24897 28679
rect 33701 28645 33735 28679
rect 39773 28645 39807 28679
rect 41797 28645 41831 28679
rect 14197 28577 14231 28611
rect 17325 28577 17359 28611
rect 17785 28577 17819 28611
rect 19165 28577 19199 28611
rect 19441 28577 19475 28611
rect 20913 28577 20947 28611
rect 22569 28577 22603 28611
rect 22845 28577 22879 28611
rect 26592 28577 26626 28611
rect 28181 28577 28215 28611
rect 28641 28577 28675 28611
rect 29653 28577 29687 28611
rect 30021 28577 30055 28611
rect 31033 28577 31067 28611
rect 32413 28577 32447 28611
rect 32689 28577 32723 28611
rect 34345 28577 34379 28611
rect 34492 28577 34526 28611
rect 36093 28577 36127 28611
rect 36461 28577 36495 28611
rect 37749 28577 37783 28611
rect 39037 28577 39071 28611
rect 39589 28577 39623 28611
rect 40601 28577 40635 28611
rect 42349 28577 42383 28611
rect 43396 28577 43430 28611
rect 45636 28577 45670 28611
rect 46581 28577 46615 28611
rect 15853 28509 15887 28543
rect 16497 28509 16531 28543
rect 22753 28509 22787 28543
rect 24501 28509 24535 28543
rect 30573 28509 30607 28543
rect 31585 28509 31619 28543
rect 34713 28509 34747 28543
rect 41705 28509 41739 28543
rect 31217 28441 31251 28475
rect 34621 28441 34655 28475
rect 14381 28373 14415 28407
rect 19993 28373 20027 28407
rect 21097 28373 21131 28407
rect 21833 28373 21867 28407
rect 25421 28373 25455 28407
rect 34805 28373 34839 28407
rect 38485 28373 38519 28407
rect 40739 28373 40773 28407
rect 41153 28373 41187 28407
rect 43499 28373 43533 28407
rect 45385 28373 45419 28407
rect 45707 28373 45741 28407
rect 46121 28373 46155 28407
rect 46765 28373 46799 28407
rect 47133 28373 47167 28407
rect 14105 28169 14139 28203
rect 15485 28169 15519 28203
rect 15853 28169 15887 28203
rect 17785 28169 17819 28203
rect 18613 28169 18647 28203
rect 19349 28169 19383 28203
rect 20913 28169 20947 28203
rect 22845 28169 22879 28203
rect 29009 28169 29043 28203
rect 30113 28169 30147 28203
rect 31033 28169 31067 28203
rect 31401 28169 31435 28203
rect 33425 28169 33459 28203
rect 34069 28169 34103 28203
rect 34437 28169 34471 28203
rect 35081 28169 35115 28203
rect 36185 28169 36219 28203
rect 37473 28169 37507 28203
rect 39405 28169 39439 28203
rect 39773 28169 39807 28203
rect 40693 28169 40727 28203
rect 42073 28169 42107 28203
rect 43453 28169 43487 28203
rect 44235 28169 44269 28203
rect 18981 28101 19015 28135
rect 30665 28101 30699 28135
rect 33149 28101 33183 28135
rect 36461 28101 36495 28135
rect 42441 28101 42475 28135
rect 19809 28033 19843 28067
rect 24501 28033 24535 28067
rect 25145 28033 25179 28067
rect 28089 28033 28123 28067
rect 31493 28033 31527 28067
rect 39129 28033 39163 28067
rect 46213 28033 46247 28067
rect 46489 28033 46523 28067
rect 13645 27965 13679 27999
rect 14197 27965 14231 27999
rect 14657 27965 14691 27999
rect 16313 27965 16347 27999
rect 16681 27965 16715 27999
rect 16957 27965 16991 27999
rect 18061 27965 18095 27999
rect 20177 27965 20211 27999
rect 20453 27965 20487 27999
rect 21649 27965 21683 27999
rect 21833 27965 21867 27999
rect 22293 27965 22327 27999
rect 23489 27965 23523 27999
rect 24041 27965 24075 27999
rect 24317 27965 24351 27999
rect 25697 27965 25731 27999
rect 28216 27965 28250 27999
rect 28641 27965 28675 27999
rect 29320 27965 29354 27999
rect 29745 27965 29779 27999
rect 30481 27965 30515 27999
rect 33241 27965 33275 27999
rect 35332 27965 35366 27999
rect 36277 27965 36311 27999
rect 36737 27965 36771 27999
rect 37289 27965 37323 27999
rect 38117 27965 38151 27999
rect 38485 27965 38519 27999
rect 38945 27965 38979 27999
rect 42660 27965 42694 27999
rect 43085 27965 43119 27999
rect 44164 27965 44198 27999
rect 13369 27897 13403 27931
rect 17141 27897 17175 27931
rect 24869 27897 24903 27931
rect 25605 27897 25639 27931
rect 26059 27897 26093 27931
rect 28319 27897 28353 27931
rect 31746 27897 31780 27931
rect 41153 27897 41187 27931
rect 41245 27897 41279 27931
rect 41981 27897 42015 27931
rect 46305 27897 46339 27931
rect 14473 27829 14507 27863
rect 17417 27829 17451 27863
rect 18245 27829 18279 27863
rect 19993 27829 20027 27863
rect 21925 27829 21959 27863
rect 26617 27829 26651 27863
rect 26985 27829 27019 27863
rect 29423 27829 29457 27863
rect 32413 27829 32447 27863
rect 32781 27829 32815 27863
rect 35403 27829 35437 27863
rect 35817 27829 35851 27863
rect 37105 27829 37139 27863
rect 37841 27829 37875 27863
rect 42763 27829 42797 27863
rect 44649 27829 44683 27863
rect 45661 27829 45695 27863
rect 47133 27829 47167 27863
rect 15393 27625 15427 27659
rect 22385 27625 22419 27659
rect 23857 27625 23891 27659
rect 26617 27625 26651 27659
rect 29377 27625 29411 27659
rect 31493 27625 31527 27659
rect 31861 27625 31895 27659
rect 32505 27625 32539 27659
rect 33333 27625 33367 27659
rect 34897 27625 34931 27659
rect 38761 27625 38795 27659
rect 39589 27625 39623 27659
rect 41153 27625 41187 27659
rect 19349 27557 19383 27591
rect 22931 27557 22965 27591
rect 25605 27557 25639 27591
rect 25881 27557 25915 27591
rect 28543 27557 28577 27591
rect 30573 27557 30607 27591
rect 35817 27557 35851 27591
rect 41797 27557 41831 27591
rect 41889 27557 41923 27591
rect 44878 27557 44912 27591
rect 46489 27557 46523 27591
rect 47041 27557 47075 27591
rect 14197 27489 14231 27523
rect 15577 27489 15611 27523
rect 15853 27489 15887 27523
rect 17233 27489 17267 27523
rect 17601 27489 17635 27523
rect 19073 27489 19107 27523
rect 21005 27489 21039 27523
rect 21465 27489 21499 27523
rect 22569 27489 22603 27523
rect 24869 27489 24903 27523
rect 25329 27489 25363 27523
rect 26525 27489 26559 27523
rect 26985 27489 27019 27523
rect 32137 27489 32171 27523
rect 34161 27489 34195 27523
rect 34345 27489 34379 27523
rect 38209 27489 38243 27523
rect 43396 27489 43430 27523
rect 44557 27489 44591 27523
rect 16497 27421 16531 27455
rect 17785 27421 17819 27455
rect 18061 27421 18095 27455
rect 21741 27421 21775 27455
rect 24685 27421 24719 27455
rect 28181 27421 28215 27455
rect 30481 27421 30515 27455
rect 34437 27421 34471 27455
rect 35725 27421 35759 27455
rect 36369 27421 36403 27455
rect 39221 27421 39255 27455
rect 42441 27421 42475 27455
rect 46397 27421 46431 27455
rect 31033 27353 31067 27387
rect 14381 27285 14415 27319
rect 19993 27285 20027 27319
rect 23489 27285 23523 27319
rect 29101 27285 29135 27319
rect 33057 27285 33091 27319
rect 35265 27285 35299 27319
rect 36737 27285 36771 27319
rect 38393 27285 38427 27319
rect 40141 27285 40175 27319
rect 40509 27285 40543 27319
rect 43499 27285 43533 27319
rect 45477 27285 45511 27319
rect 46121 27285 46155 27319
rect 13737 27081 13771 27115
rect 17509 27081 17543 27115
rect 21097 27081 21131 27115
rect 23397 27081 23431 27115
rect 26433 27081 26467 27115
rect 26801 27081 26835 27115
rect 28733 27081 28767 27115
rect 30113 27081 30147 27115
rect 30389 27081 30423 27115
rect 38117 27081 38151 27115
rect 42073 27081 42107 27115
rect 44189 27081 44223 27115
rect 45155 27081 45189 27115
rect 47501 27081 47535 27115
rect 24225 27013 24259 27047
rect 24593 27013 24627 27047
rect 29101 27013 29135 27047
rect 14841 26945 14875 26979
rect 17141 26945 17175 26979
rect 18061 26945 18095 26979
rect 19809 26945 19843 26979
rect 21833 26945 21867 26979
rect 24869 26945 24903 26979
rect 25605 26945 25639 26979
rect 29377 26945 29411 26979
rect 29837 26945 29871 26979
rect 14381 26877 14415 26911
rect 14749 26877 14783 26911
rect 15761 26877 15795 26911
rect 16129 26877 16163 26911
rect 16405 26877 16439 26911
rect 24041 26877 24075 26911
rect 25053 26877 25087 26911
rect 25513 26877 25547 26911
rect 26617 26877 26651 26911
rect 27537 26877 27571 26911
rect 27905 26877 27939 26911
rect 28181 26877 28215 26911
rect 18382 26809 18416 26843
rect 19257 26809 19291 26843
rect 19625 26809 19659 26843
rect 20130 26809 20164 26843
rect 21649 26809 21683 26843
rect 22154 26809 22188 26843
rect 23029 26809 23063 26843
rect 26065 26809 26099 26843
rect 28365 26809 28399 26843
rect 29446 26809 29480 26843
rect 34253 27013 34287 27047
rect 37289 27013 37323 27047
rect 46765 27013 46799 27047
rect 30941 26945 30975 26979
rect 31217 26945 31251 26979
rect 33977 26945 34011 26979
rect 34897 26945 34931 26979
rect 36737 26945 36771 26979
rect 38301 26945 38335 26979
rect 38577 26945 38611 26979
rect 42717 26945 42751 26979
rect 43269 26945 43303 26979
rect 43913 26945 43947 26979
rect 33057 26877 33091 26911
rect 33517 26877 33551 26911
rect 33793 26877 33827 26911
rect 40509 26877 40543 26911
rect 45052 26877 45086 26911
rect 30757 26809 30791 26843
rect 31033 26809 31067 26843
rect 32781 26809 32815 26843
rect 35218 26809 35252 26843
rect 36461 26809 36495 26843
rect 36829 26809 36863 26843
rect 37749 26809 37783 26843
rect 38393 26809 38427 26843
rect 39313 26809 39347 26843
rect 40233 26809 40267 26843
rect 40830 26809 40864 26843
rect 43085 26809 43119 26843
rect 43361 26809 43395 26843
rect 46213 26809 46247 26843
rect 46305 26809 46339 26843
rect 14197 26741 14231 26775
rect 15393 26741 15427 26775
rect 15945 26741 15979 26775
rect 17785 26741 17819 26775
rect 18981 26741 19015 26775
rect 20729 26741 20763 26775
rect 22753 26741 22787 26775
rect 27077 26741 27111 26775
rect 30113 26741 30147 26775
rect 32229 26741 32263 26775
rect 34621 26741 34655 26775
rect 35817 26741 35851 26775
rect 36185 26741 36219 26775
rect 39589 26741 39623 26775
rect 41429 26741 41463 26775
rect 41797 26741 41831 26775
rect 44557 26741 44591 26775
rect 45477 26741 45511 26775
rect 45845 26741 45879 26775
rect 47133 26741 47167 26775
rect 15117 26537 15151 26571
rect 16497 26537 16531 26571
rect 18061 26537 18095 26571
rect 19349 26537 19383 26571
rect 19901 26537 19935 26571
rect 21465 26537 21499 26571
rect 21925 26537 21959 26571
rect 27721 26537 27755 26571
rect 28457 26537 28491 26571
rect 29469 26537 29503 26571
rect 30159 26537 30193 26571
rect 30481 26537 30515 26571
rect 30941 26537 30975 26571
rect 32689 26537 32723 26571
rect 33425 26537 33459 26571
rect 33885 26537 33919 26571
rect 34621 26537 34655 26571
rect 38071 26537 38105 26571
rect 44557 26537 44591 26571
rect 46673 26537 46707 26571
rect 15577 26469 15611 26503
rect 18521 26469 18555 26503
rect 22706 26469 22740 26503
rect 36093 26469 36127 26503
rect 36185 26469 36219 26503
rect 39681 26469 39715 26503
rect 41889 26469 41923 26503
rect 42441 26469 42475 26503
rect 43545 26469 43579 26503
rect 45845 26469 45879 26503
rect 15301 26401 15335 26435
rect 17360 26401 17394 26435
rect 20980 26401 21014 26435
rect 22385 26401 22419 26435
rect 24777 26401 24811 26435
rect 25237 26401 25271 26435
rect 25789 26401 25823 26435
rect 26709 26401 26743 26435
rect 27052 26401 27086 26435
rect 29009 26401 29043 26435
rect 30021 26401 30055 26435
rect 31068 26401 31102 26435
rect 32229 26401 32263 26435
rect 33241 26401 33275 26435
rect 34253 26401 34287 26435
rect 37841 26401 37875 26435
rect 38945 26401 38979 26435
rect 39405 26401 39439 26435
rect 40544 26401 40578 26435
rect 47260 26401 47294 26435
rect 18429 26333 18463 26367
rect 18705 26333 18739 26367
rect 25329 26333 25363 26367
rect 27905 26333 27939 26367
rect 36369 26333 36403 26367
rect 41613 26333 41647 26367
rect 41797 26333 41831 26367
rect 43453 26333 43487 26367
rect 43729 26333 43763 26367
rect 45753 26333 45787 26367
rect 47363 26333 47397 26367
rect 32413 26265 32447 26299
rect 35173 26265 35207 26299
rect 46305 26265 46339 26299
rect 14381 26197 14415 26231
rect 16221 26197 16255 26231
rect 17463 26197 17497 26231
rect 21051 26197 21085 26231
rect 22201 26197 22235 26231
rect 23305 26197 23339 26231
rect 27123 26197 27157 26231
rect 28135 26197 28169 26231
rect 29147 26197 29181 26231
rect 31171 26197 31205 26231
rect 35633 26197 35667 26231
rect 38393 26197 38427 26231
rect 40647 26197 40681 26231
rect 40969 26197 41003 26231
rect 16405 25993 16439 26027
rect 16865 25993 16899 26027
rect 19257 25993 19291 26027
rect 21373 25993 21407 26027
rect 22937 25993 22971 26027
rect 24777 25993 24811 26027
rect 28089 25993 28123 26027
rect 32137 25993 32171 26027
rect 33333 25993 33367 26027
rect 33931 25993 33965 26027
rect 36507 25993 36541 26027
rect 39589 25993 39623 26027
rect 40693 25993 40727 26027
rect 41981 25993 42015 26027
rect 42533 25993 42567 26027
rect 42901 25993 42935 26027
rect 43269 25993 43303 26027
rect 44833 25993 44867 26027
rect 45845 25993 45879 26027
rect 46397 25993 46431 26027
rect 24225 25925 24259 25959
rect 29101 25925 29135 25959
rect 30389 25925 30423 25959
rect 45063 25925 45097 25959
rect 14841 25857 14875 25891
rect 18061 25857 18095 25891
rect 20085 25857 20119 25891
rect 20361 25857 20395 25891
rect 21649 25857 21683 25891
rect 22569 25857 22603 25891
rect 22753 25857 22787 25891
rect 25605 25857 25639 25891
rect 29377 25857 29411 25891
rect 31769 25857 31803 25891
rect 34713 25857 34747 25891
rect 37657 25857 37691 25891
rect 38945 25857 38979 25891
rect 41061 25857 41095 25891
rect 41705 25857 41739 25891
rect 43453 25857 43487 25891
rect 17785 25789 17819 25823
rect 15203 25721 15237 25755
rect 16037 25721 16071 25755
rect 17417 25721 17451 25755
rect 18382 25721 18416 25755
rect 19901 25721 19935 25755
rect 20177 25721 20211 25755
rect 21741 25721 21775 25755
rect 22293 25721 22327 25755
rect 23724 25789 23758 25823
rect 27077 25789 27111 25823
rect 28232 25789 28266 25823
rect 28733 25789 28767 25823
rect 31284 25789 31318 25823
rect 32264 25789 32298 25823
rect 32689 25789 32723 25823
rect 33860 25789 33894 25823
rect 34964 25789 34998 25823
rect 36436 25789 36470 25823
rect 38485 25789 38519 25823
rect 38761 25789 38795 25823
rect 44960 25789 44994 25823
rect 45385 25789 45419 25823
rect 46156 25789 46190 25823
rect 46581 25789 46615 25823
rect 47168 25789 47202 25823
rect 47961 25789 47995 25823
rect 23811 25721 23845 25755
rect 25421 25721 25455 25755
rect 25926 25721 25960 25755
rect 28319 25721 28353 25755
rect 29469 25721 29503 25755
rect 30021 25721 30055 25755
rect 41153 25721 41187 25755
rect 43545 25721 43579 25755
rect 44097 25721 44131 25755
rect 44465 25721 44499 25755
rect 47271 25721 47305 25755
rect 14749 25653 14783 25687
rect 15761 25653 15795 25687
rect 16957 25653 16991 25687
rect 18981 25653 19015 25687
rect 21097 25653 21131 25687
rect 22753 25653 22787 25687
rect 26525 25653 26559 25687
rect 31033 25653 31067 25687
rect 31355 25653 31389 25687
rect 32367 25653 32401 25687
rect 34345 25653 34379 25687
rect 35035 25653 35069 25687
rect 35357 25653 35391 25687
rect 36001 25653 36035 25687
rect 36921 25653 36955 25687
rect 38025 25653 38059 25687
rect 39221 25653 39255 25687
rect 47593 25653 47627 25687
rect 14841 25449 14875 25483
rect 16497 25449 16531 25483
rect 20085 25449 20119 25483
rect 21695 25449 21729 25483
rect 23673 25449 23707 25483
rect 24777 25449 24811 25483
rect 25881 25449 25915 25483
rect 26893 25449 26927 25483
rect 29745 25449 29779 25483
rect 31861 25449 31895 25483
rect 34345 25449 34379 25483
rect 34713 25449 34747 25483
rect 36093 25449 36127 25483
rect 36507 25449 36541 25483
rect 41061 25449 41095 25483
rect 15622 25381 15656 25415
rect 17233 25381 17267 25415
rect 18705 25381 18739 25415
rect 18797 25381 18831 25415
rect 22109 25381 22143 25415
rect 22753 25381 22787 25415
rect 25053 25381 25087 25415
rect 28917 25381 28951 25415
rect 30665 25381 30699 25415
rect 32321 25381 32355 25415
rect 34989 25381 35023 25415
rect 41797 25381 41831 25415
rect 43545 25381 43579 25415
rect 45385 25381 45419 25415
rect 15301 25313 15335 25347
rect 17785 25313 17819 25347
rect 21465 25313 21499 25347
rect 26525 25313 26559 25347
rect 33844 25313 33878 25347
rect 36404 25313 36438 25347
rect 37657 25313 37691 25347
rect 39221 25313 39255 25347
rect 39681 25313 39715 25347
rect 17141 25245 17175 25279
rect 18981 25245 19015 25279
rect 22661 25245 22695 25279
rect 23305 25245 23339 25279
rect 24961 25245 24995 25279
rect 25605 25245 25639 25279
rect 28825 25245 28859 25279
rect 29469 25245 29503 25279
rect 30573 25245 30607 25279
rect 30849 25245 30883 25279
rect 32229 25245 32263 25279
rect 32505 25245 32539 25279
rect 33931 25245 33965 25279
rect 34897 25245 34931 25279
rect 38301 25245 38335 25279
rect 39957 25245 39991 25279
rect 41521 25245 41555 25279
rect 41705 25245 41739 25279
rect 41981 25245 42015 25279
rect 43453 25245 43487 25279
rect 43729 25245 43763 25279
rect 45293 25245 45327 25279
rect 45569 25245 45603 25279
rect 46765 25245 46799 25279
rect 16865 25177 16899 25211
rect 35449 25177 35483 25211
rect 37887 25177 37921 25211
rect 38577 25177 38611 25211
rect 16221 25109 16255 25143
rect 18429 25109 18463 25143
rect 20361 25109 20395 25143
rect 27445 25109 27479 25143
rect 36921 25109 36955 25143
rect 44557 25109 44591 25143
rect 46305 25109 46339 25143
rect 14933 24905 14967 24939
rect 17141 24905 17175 24939
rect 17417 24905 17451 24939
rect 19349 24905 19383 24939
rect 19809 24905 19843 24939
rect 23397 24905 23431 24939
rect 25145 24905 25179 24939
rect 28089 24905 28123 24939
rect 28825 24905 28859 24939
rect 31033 24905 31067 24939
rect 31309 24905 31343 24939
rect 31401 24905 31435 24939
rect 32597 24905 32631 24939
rect 32965 24905 32999 24939
rect 34621 24905 34655 24939
rect 37841 24905 37875 24939
rect 39313 24905 39347 24939
rect 39681 24905 39715 24939
rect 43913 24905 43947 24939
rect 16681 24837 16715 24871
rect 24869 24837 24903 24871
rect 26249 24837 26283 24871
rect 15163 24769 15197 24803
rect 17785 24769 17819 24803
rect 18429 24769 18463 24803
rect 18705 24769 18739 24803
rect 22385 24769 22419 24803
rect 23765 24769 23799 24803
rect 24041 24769 24075 24803
rect 25329 24769 25363 24803
rect 27445 24769 27479 24803
rect 30389 24769 30423 24803
rect 15076 24701 15110 24735
rect 32229 24837 32263 24871
rect 36369 24837 36403 24871
rect 40325 24837 40359 24871
rect 46765 24837 46799 24871
rect 31677 24769 31711 24803
rect 33241 24769 33275 24803
rect 33517 24769 33551 24803
rect 34989 24769 35023 24803
rect 35449 24769 35483 24803
rect 37473 24769 37507 24803
rect 38393 24769 38427 24803
rect 38669 24769 38703 24803
rect 40877 24769 40911 24803
rect 41521 24769 41555 24803
rect 44557 24769 44591 24803
rect 44833 24769 44867 24803
rect 45937 24769 45971 24803
rect 46213 24769 46247 24803
rect 42349 24701 42383 24735
rect 16129 24633 16163 24667
rect 16221 24633 16255 24667
rect 18521 24633 18555 24667
rect 19993 24633 20027 24667
rect 20085 24633 20119 24667
rect 20637 24633 20671 24667
rect 21281 24633 21315 24667
rect 22109 24633 22143 24667
rect 22201 24633 22235 24667
rect 23857 24633 23891 24667
rect 25650 24633 25684 24667
rect 27169 24633 27203 24667
rect 27261 24633 27295 24667
rect 29561 24633 29595 24667
rect 30113 24633 30147 24667
rect 30205 24633 30239 24667
rect 31309 24633 31343 24667
rect 31769 24633 31803 24667
rect 33333 24633 33367 24667
rect 34253 24633 34287 24667
rect 35081 24633 35115 24667
rect 36001 24633 36035 24667
rect 36829 24633 36863 24667
rect 36921 24633 36955 24667
rect 38209 24633 38243 24667
rect 38485 24633 38519 24667
rect 40969 24633 41003 24667
rect 42670 24633 42704 24667
rect 44649 24633 44683 24667
rect 45569 24633 45603 24667
rect 46305 24633 46339 24667
rect 15485 24565 15519 24599
rect 15945 24565 15979 24599
rect 21557 24565 21591 24599
rect 23029 24565 23063 24599
rect 26525 24565 26559 24599
rect 26985 24565 27019 24599
rect 29929 24565 29963 24599
rect 41797 24565 41831 24599
rect 42165 24565 42199 24599
rect 43269 24565 43303 24599
rect 43545 24565 43579 24599
rect 44373 24565 44407 24599
rect 14335 24361 14369 24395
rect 18705 24361 18739 24395
rect 22753 24361 22787 24395
rect 25881 24361 25915 24395
rect 27537 24361 27571 24395
rect 28549 24361 28583 24395
rect 29377 24361 29411 24395
rect 30159 24361 30193 24395
rect 30573 24361 30607 24395
rect 31677 24361 31711 24395
rect 33241 24361 33275 24395
rect 35541 24361 35575 24395
rect 40417 24361 40451 24395
rect 42165 24361 42199 24395
rect 45201 24361 45235 24395
rect 45477 24361 45511 24395
rect 16221 24293 16255 24327
rect 16773 24293 16807 24327
rect 19349 24293 19383 24327
rect 21833 24293 21867 24327
rect 21925 24293 21959 24327
rect 23489 24293 23523 24327
rect 25053 24293 25087 24327
rect 26709 24293 26743 24327
rect 27261 24293 27295 24327
rect 32229 24293 32263 24327
rect 32321 24293 32355 24327
rect 32873 24293 32907 24327
rect 34666 24293 34700 24327
rect 36277 24293 36311 24327
rect 39859 24293 39893 24327
rect 41566 24293 41600 24327
rect 44602 24293 44636 24327
rect 46213 24293 46247 24327
rect 18204 24225 18238 24259
rect 30088 24225 30122 24259
rect 31068 24225 31102 24259
rect 37933 24225 37967 24259
rect 38485 24225 38519 24259
rect 14105 24157 14139 24191
rect 15945 24157 15979 24191
rect 16129 24157 16163 24191
rect 18291 24157 18325 24191
rect 19257 24157 19291 24191
rect 19901 24157 19935 24191
rect 22477 24157 22511 24191
rect 23397 24157 23431 24191
rect 24961 24157 24995 24191
rect 25237 24157 25271 24191
rect 26617 24157 26651 24191
rect 28181 24157 28215 24191
rect 34345 24157 34379 24191
rect 36185 24157 36219 24191
rect 37105 24157 37139 24191
rect 38669 24157 38703 24191
rect 39497 24157 39531 24191
rect 41245 24157 41279 24191
rect 44281 24157 44315 24191
rect 46121 24157 46155 24191
rect 46489 24157 46523 24191
rect 23949 24089 23983 24123
rect 24685 24089 24719 24123
rect 31171 24089 31205 24123
rect 35265 24089 35299 24123
rect 36737 24089 36771 24123
rect 18061 24021 18095 24055
rect 20177 24021 20211 24055
rect 29101 24021 29135 24055
rect 34161 24021 34195 24055
rect 35909 24021 35943 24055
rect 40877 24021 40911 24055
rect 42441 24021 42475 24055
rect 14105 23817 14139 23851
rect 15945 23817 15979 23851
rect 17877 23817 17911 23851
rect 19257 23817 19291 23851
rect 20637 23817 20671 23851
rect 21465 23817 21499 23851
rect 22109 23817 22143 23851
rect 22339 23817 22373 23851
rect 22753 23817 22787 23851
rect 23811 23817 23845 23851
rect 24869 23817 24903 23851
rect 25881 23817 25915 23851
rect 26433 23817 26467 23851
rect 26801 23817 26835 23851
rect 28641 23817 28675 23851
rect 29101 23817 29135 23851
rect 30987 23817 31021 23851
rect 31309 23817 31343 23851
rect 32505 23817 32539 23851
rect 32919 23817 32953 23851
rect 36737 23817 36771 23851
rect 37933 23817 37967 23851
rect 38393 23817 38427 23851
rect 42257 23817 42291 23851
rect 43085 23817 43119 23851
rect 44879 23817 44913 23851
rect 45845 23817 45879 23851
rect 17049 23749 17083 23783
rect 18705 23749 18739 23783
rect 25099 23749 25133 23783
rect 25513 23749 25547 23783
rect 31769 23749 31803 23783
rect 36093 23749 36127 23783
rect 41613 23749 41647 23783
rect 46259 23749 46293 23783
rect 14657 23681 14691 23715
rect 16497 23681 16531 23715
rect 18153 23681 18187 23715
rect 19717 23681 19751 23715
rect 21649 23681 21683 23715
rect 23397 23681 23431 23715
rect 28181 23681 28215 23715
rect 29837 23681 29871 23715
rect 30297 23681 30331 23715
rect 32229 23681 32263 23715
rect 33931 23681 33965 23715
rect 34989 23681 35023 23715
rect 35357 23681 35391 23715
rect 37565 23681 37599 23715
rect 40693 23681 40727 23715
rect 42717 23681 42751 23715
rect 43269 23681 43303 23715
rect 43637 23681 43671 23715
rect 15577 23613 15611 23647
rect 16221 23613 16255 23647
rect 21256 23613 21290 23647
rect 22268 23613 22302 23647
rect 23740 23613 23774 23647
rect 25028 23613 25062 23647
rect 26040 23613 26074 23647
rect 27445 23613 27479 23647
rect 27629 23613 27663 23647
rect 28089 23613 28123 23647
rect 30916 23613 30950 23647
rect 32848 23613 32882 23647
rect 33241 23613 33275 23647
rect 33828 23613 33862 23647
rect 38853 23613 38887 23647
rect 39405 23613 39439 23647
rect 39589 23613 39623 23647
rect 44808 23613 44842 23647
rect 45201 23613 45235 23647
rect 46156 23613 46190 23647
rect 46581 23613 46615 23647
rect 14565 23545 14599 23579
rect 14978 23545 15012 23579
rect 16589 23545 16623 23579
rect 17509 23545 17543 23579
rect 18245 23545 18279 23579
rect 19809 23545 19843 23579
rect 20361 23545 20395 23579
rect 24225 23545 24259 23579
rect 29377 23545 29411 23579
rect 29469 23545 29503 23579
rect 33701 23545 33735 23579
rect 35081 23545 35115 23579
rect 36921 23545 36955 23579
rect 37013 23545 37047 23579
rect 41014 23545 41048 23579
rect 41889 23545 41923 23579
rect 43361 23545 43395 23579
rect 26111 23477 26145 23511
rect 34437 23477 34471 23511
rect 38669 23477 38703 23511
rect 39957 23477 39991 23511
rect 40325 23477 40359 23511
rect 44281 23477 44315 23511
rect 14657 23273 14691 23307
rect 19257 23273 19291 23307
rect 21833 23273 21867 23307
rect 23397 23273 23431 23307
rect 24961 23273 24995 23307
rect 28181 23273 28215 23307
rect 33241 23273 33275 23307
rect 34069 23273 34103 23307
rect 34989 23273 35023 23307
rect 36185 23273 36219 23307
rect 36691 23273 36725 23307
rect 37013 23273 37047 23307
rect 40325 23273 40359 23307
rect 40693 23273 40727 23307
rect 44281 23273 44315 23307
rect 44695 23273 44729 23307
rect 46121 23273 46155 23307
rect 15853 23205 15887 23239
rect 16405 23205 16439 23239
rect 18245 23205 18279 23239
rect 18797 23205 18831 23239
rect 22569 23205 22603 23239
rect 26709 23205 26743 23239
rect 27261 23205 27295 23239
rect 29561 23205 29595 23239
rect 29653 23205 29687 23239
rect 32321 23205 32355 23239
rect 32873 23205 32907 23239
rect 40049 23205 40083 23239
rect 41613 23205 41647 23239
rect 14105 23137 14139 23171
rect 19625 23137 19659 23171
rect 21373 23137 21407 23171
rect 23213 23137 23247 23171
rect 24016 23137 24050 23171
rect 25180 23137 25214 23171
rect 34069 23137 34103 23171
rect 34253 23137 34287 23171
rect 35424 23137 35458 23171
rect 36553 23137 36587 23171
rect 37657 23137 37691 23171
rect 39313 23137 39347 23171
rect 39865 23137 39899 23171
rect 40877 23137 40911 23171
rect 41337 23137 41371 23171
rect 43428 23137 43462 23171
rect 44624 23137 44658 23171
rect 15761 23069 15795 23103
rect 18153 23069 18187 23103
rect 19763 23069 19797 23103
rect 22477 23069 22511 23103
rect 22753 23069 22787 23103
rect 26617 23069 26651 23103
rect 28365 23069 28399 23103
rect 30021 23069 30055 23103
rect 31033 23069 31067 23103
rect 32229 23069 32263 23103
rect 38945 23069 38979 23103
rect 23213 23001 23247 23035
rect 25605 23001 25639 23035
rect 14335 22933 14369 22967
rect 16681 22933 16715 22967
rect 20177 22933 20211 22967
rect 21557 22933 21591 22967
rect 23857 22933 23891 22967
rect 24087 22933 24121 22967
rect 25283 22933 25317 22967
rect 27721 22933 27755 22967
rect 28595 22933 28629 22967
rect 29377 22933 29411 22967
rect 35495 22933 35529 22967
rect 37887 22933 37921 22967
rect 43499 22933 43533 22967
rect 14289 22729 14323 22763
rect 15669 22729 15703 22763
rect 17509 22729 17543 22763
rect 17785 22729 17819 22763
rect 21925 22729 21959 22763
rect 23121 22729 23155 22763
rect 25145 22729 25179 22763
rect 26433 22729 26467 22763
rect 30987 22729 31021 22763
rect 31861 22729 31895 22763
rect 32229 22729 32263 22763
rect 33885 22729 33919 22763
rect 36645 22729 36679 22763
rect 38945 22729 38979 22763
rect 39957 22729 39991 22763
rect 44005 22729 44039 22763
rect 20637 22661 20671 22695
rect 21465 22661 21499 22695
rect 29929 22661 29963 22695
rect 35541 22661 35575 22695
rect 38117 22661 38151 22695
rect 42809 22661 42843 22695
rect 14887 22593 14921 22627
rect 16497 22593 16531 22627
rect 18429 22593 18463 22627
rect 22385 22593 22419 22627
rect 23857 22593 23891 22627
rect 24869 22593 24903 22627
rect 25697 22593 25731 22627
rect 26985 22593 27019 22627
rect 27261 22593 27295 22627
rect 29377 22593 29411 22627
rect 30665 22593 30699 22627
rect 32505 22593 32539 22627
rect 32781 22593 32815 22627
rect 34989 22593 35023 22627
rect 37197 22593 37231 22627
rect 37473 22593 37507 22627
rect 43085 22593 43119 22627
rect 46259 22593 46293 22627
rect 14800 22525 14834 22559
rect 30389 22525 30423 22559
rect 30884 22525 30918 22559
rect 39472 22525 39506 22559
rect 41404 22525 41438 22559
rect 41797 22525 41831 22559
rect 44592 22525 44626 22559
rect 45385 22525 45419 22559
rect 46156 22525 46190 22559
rect 46581 22525 46615 22559
rect 15853 22457 15887 22491
rect 15945 22457 15979 22491
rect 18153 22457 18187 22491
rect 18245 22457 18279 22491
rect 20085 22457 20119 22491
rect 20177 22457 20211 22491
rect 22109 22457 22143 22491
rect 22201 22457 22235 22491
rect 23489 22457 23523 22491
rect 23949 22457 23983 22491
rect 24501 22457 24535 22491
rect 25421 22457 25455 22491
rect 25513 22457 25547 22491
rect 27077 22457 27111 22491
rect 29101 22457 29135 22491
rect 29469 22457 29503 22491
rect 31309 22457 31343 22491
rect 32597 22457 32631 22491
rect 34713 22457 34747 22491
rect 35081 22457 35115 22491
rect 37013 22457 37047 22491
rect 37289 22457 37323 22491
rect 40877 22457 40911 22491
rect 43177 22457 43211 22491
rect 43729 22457 43763 22491
rect 15301 22389 15335 22423
rect 16773 22389 16807 22423
rect 19073 22389 19107 22423
rect 19717 22389 19751 22423
rect 26709 22389 26743 22423
rect 28549 22389 28583 22423
rect 33425 22389 33459 22423
rect 34161 22389 34195 22423
rect 36001 22389 36035 22423
rect 39313 22389 39347 22423
rect 39543 22389 39577 22423
rect 41475 22389 41509 22423
rect 44695 22389 44729 22423
rect 45017 22389 45051 22423
rect 15853 22185 15887 22219
rect 16129 22185 16163 22219
rect 18015 22185 18049 22219
rect 18337 22185 18371 22219
rect 21695 22185 21729 22219
rect 22109 22185 22143 22219
rect 22477 22185 22511 22219
rect 23765 22185 23799 22219
rect 25697 22185 25731 22219
rect 26985 22185 27019 22219
rect 27353 22185 27387 22219
rect 29561 22185 29595 22219
rect 32505 22185 32539 22219
rect 33057 22185 33091 22219
rect 34805 22185 34839 22219
rect 35173 22185 35207 22219
rect 37197 22185 37231 22219
rect 40969 22185 41003 22219
rect 43085 22185 43119 22219
rect 15439 22117 15473 22151
rect 19441 22117 19475 22151
rect 19993 22117 20027 22151
rect 22753 22117 22787 22151
rect 24317 22117 24351 22151
rect 27675 22117 27709 22151
rect 28962 22117 28996 22151
rect 30573 22117 30607 22151
rect 34247 22117 34281 22151
rect 35817 22117 35851 22151
rect 36369 22117 36403 22151
rect 37933 22117 37967 22151
rect 38485 22117 38519 22151
rect 41429 22117 41463 22151
rect 43453 22117 43487 22151
rect 43545 22117 43579 22151
rect 45385 22117 45419 22151
rect 15336 22049 15370 22083
rect 16932 22049 16966 22083
rect 17944 22049 17978 22083
rect 21624 22049 21658 22083
rect 26592 22049 26626 22083
rect 27572 22049 27606 22083
rect 29837 22049 29871 22083
rect 31125 22049 31159 22083
rect 40268 22049 40302 22083
rect 46765 22049 46799 22083
rect 19349 21981 19383 22015
rect 22661 21981 22695 22015
rect 22937 21981 22971 22015
rect 24225 21981 24259 22015
rect 24501 21981 24535 22015
rect 25421 21981 25455 22015
rect 28641 21981 28675 22015
rect 30481 21981 30515 22015
rect 32137 21981 32171 22015
rect 33885 21981 33919 22015
rect 35725 21981 35759 22015
rect 37841 21981 37875 22015
rect 40371 21981 40405 22015
rect 41337 21981 41371 22015
rect 41613 21981 41647 22015
rect 45293 21981 45327 22015
rect 45569 21981 45603 22015
rect 17003 21913 17037 21947
rect 20269 21913 20303 21947
rect 44005 21913 44039 21947
rect 26663 21845 26697 21879
rect 31585 21845 31619 21879
rect 36737 21845 36771 21879
rect 37473 21845 37507 21879
rect 44557 21845 44591 21879
rect 46903 21845 46937 21879
rect 17095 21641 17129 21675
rect 18981 21641 19015 21675
rect 19763 21641 19797 21675
rect 20177 21641 20211 21675
rect 21235 21641 21269 21675
rect 23029 21641 23063 21675
rect 24777 21641 24811 21675
rect 25237 21641 25271 21675
rect 26617 21641 26651 21675
rect 27445 21641 27479 21675
rect 28641 21641 28675 21675
rect 29009 21641 29043 21675
rect 30573 21641 30607 21675
rect 32597 21641 32631 21675
rect 34345 21641 34379 21675
rect 35725 21641 35759 21675
rect 36093 21641 36127 21675
rect 38393 21641 38427 21675
rect 39865 21641 39899 21675
rect 41429 21641 41463 21675
rect 41797 21641 41831 21675
rect 43729 21641 43763 21675
rect 45845 21641 45879 21675
rect 47271 21641 47305 21675
rect 16083 21573 16117 21607
rect 30849 21573 30883 21607
rect 46949 21573 46983 21607
rect 16497 21505 16531 21539
rect 19349 21505 19383 21539
rect 22569 21505 22603 21539
rect 24501 21505 24535 21539
rect 25421 21505 25455 21539
rect 25697 21505 25731 21539
rect 31677 21505 31711 21539
rect 33977 21505 34011 21539
rect 34621 21505 34655 21539
rect 34989 21505 35023 21539
rect 42349 21505 42383 21539
rect 42993 21505 43027 21539
rect 43453 21505 43487 21539
rect 44557 21505 44591 21539
rect 46259 21505 46293 21539
rect 16012 21437 16046 21471
rect 17024 21437 17058 21471
rect 19692 21437 19726 21471
rect 21005 21437 21039 21471
rect 21132 21437 21166 21471
rect 22144 21437 22178 21471
rect 27629 21437 27663 21471
rect 28181 21437 28215 21471
rect 29285 21437 29319 21471
rect 33241 21437 33275 21471
rect 33701 21437 33735 21471
rect 36645 21437 36679 21471
rect 38577 21437 38611 21471
rect 39037 21437 39071 21471
rect 39313 21437 39347 21471
rect 40509 21437 40543 21471
rect 46172 21437 46206 21471
rect 47200 21437 47234 21471
rect 47593 21437 47627 21471
rect 17509 21369 17543 21403
rect 22247 21369 22281 21403
rect 23489 21369 23523 21403
rect 23857 21369 23891 21403
rect 23949 21369 23983 21403
rect 25513 21369 25547 21403
rect 27169 21369 27203 21403
rect 28365 21369 28399 21403
rect 29606 21369 29640 21403
rect 31769 21369 31803 21403
rect 32321 21369 32355 21403
rect 33149 21369 33183 21403
rect 36966 21369 37000 21403
rect 40830 21369 40864 21403
rect 42441 21369 42475 21403
rect 44373 21369 44407 21403
rect 44649 21369 44683 21403
rect 45201 21369 45235 21403
rect 15301 21301 15335 21335
rect 16865 21301 16899 21335
rect 18061 21301 18095 21335
rect 18613 21301 18647 21335
rect 21005 21301 21039 21335
rect 21557 21301 21591 21335
rect 22017 21301 22051 21335
rect 30205 21301 30239 21335
rect 31493 21301 31527 21335
rect 36461 21301 36495 21335
rect 37565 21301 37599 21335
rect 38117 21301 38151 21335
rect 40325 21301 40359 21335
rect 42073 21301 42107 21335
rect 45477 21301 45511 21335
rect 46673 21301 46707 21335
rect 17095 21097 17129 21131
rect 22753 21097 22787 21131
rect 23581 21097 23615 21131
rect 24225 21097 24259 21131
rect 27629 21097 27663 21131
rect 28917 21097 28951 21131
rect 31953 21097 31987 21131
rect 32229 21097 32263 21131
rect 37473 21097 37507 21131
rect 40509 21097 40543 21131
rect 41061 21097 41095 21131
rect 42349 21097 42383 21131
rect 44833 21097 44867 21131
rect 18153 21029 18187 21063
rect 22431 21029 22465 21063
rect 28641 21029 28675 21063
rect 29285 21029 29319 21063
rect 29837 21029 29871 21063
rect 30389 21029 30423 21063
rect 36001 21029 36035 21063
rect 37933 21029 37967 21063
rect 41429 21029 41463 21063
rect 44234 21029 44268 21063
rect 45753 21029 45787 21063
rect 45845 21029 45879 21063
rect 17003 20961 17037 20995
rect 19568 20961 19602 20995
rect 19993 20961 20027 20995
rect 22344 20961 22378 20995
rect 25421 20961 25455 20995
rect 26560 20961 26594 20995
rect 28089 20961 28123 20995
rect 28457 20961 28491 20995
rect 32413 20961 32447 20995
rect 32689 20961 32723 20995
rect 34161 20961 34195 20995
rect 34621 20961 34655 20995
rect 39313 20961 39347 20995
rect 39773 20961 39807 20995
rect 42073 20961 42107 20995
rect 18061 20893 18095 20927
rect 18705 20893 18739 20927
rect 21281 20893 21315 20927
rect 29745 20893 29779 20927
rect 34805 20893 34839 20927
rect 35081 20893 35115 20927
rect 35909 20893 35943 20927
rect 37841 20893 37875 20927
rect 38209 20893 38243 20927
rect 40049 20893 40083 20927
rect 41337 20893 41371 20927
rect 43913 20893 43947 20927
rect 46029 20893 46063 20927
rect 25605 20825 25639 20859
rect 36461 20825 36495 20859
rect 41889 20825 41923 20859
rect 42073 20825 42107 20859
rect 19671 20757 19705 20791
rect 26663 20757 26697 20791
rect 31033 20757 31067 20791
rect 33333 20757 33367 20791
rect 38945 20757 38979 20791
rect 17233 20553 17267 20587
rect 17509 20553 17543 20587
rect 17785 20553 17819 20587
rect 18981 20553 19015 20587
rect 19257 20553 19291 20587
rect 21373 20553 21407 20587
rect 22661 20553 22695 20587
rect 25881 20553 25915 20587
rect 27077 20553 27111 20587
rect 27537 20553 27571 20587
rect 30481 20553 30515 20587
rect 30849 20553 30883 20587
rect 31953 20553 31987 20587
rect 32321 20553 32355 20587
rect 32689 20553 32723 20587
rect 32965 20553 32999 20587
rect 34621 20553 34655 20587
rect 37749 20553 37783 20587
rect 38117 20553 38151 20587
rect 38761 20553 38795 20587
rect 39865 20553 39899 20587
rect 42901 20553 42935 20587
rect 44373 20553 44407 20587
rect 44925 20553 44959 20587
rect 45845 20553 45879 20587
rect 16865 20485 16899 20519
rect 28733 20485 28767 20519
rect 33793 20485 33827 20519
rect 44005 20485 44039 20519
rect 45293 20485 45327 20519
rect 45569 20485 45603 20519
rect 21649 20417 21683 20451
rect 31033 20417 31067 20451
rect 34897 20417 34931 20451
rect 36185 20417 36219 20451
rect 43729 20417 43763 20451
rect 16497 20349 16531 20383
rect 16992 20349 17026 20383
rect 18061 20349 18095 20383
rect 19993 20349 20027 20383
rect 20453 20349 20487 20383
rect 23740 20349 23774 20383
rect 24133 20349 24167 20383
rect 25120 20349 25154 20383
rect 25513 20349 25547 20383
rect 26525 20349 26559 20383
rect 27721 20349 27755 20383
rect 29469 20349 29503 20383
rect 32781 20349 32815 20383
rect 33241 20349 33275 20383
rect 36461 20349 36495 20383
rect 36645 20349 36679 20383
rect 37105 20349 37139 20383
rect 38853 20349 38887 20383
rect 39313 20349 39347 20383
rect 39589 20349 39623 20383
rect 40509 20349 40543 20383
rect 45068 20349 45102 20383
rect 45293 20349 45327 20383
rect 18382 20281 18416 20315
rect 19901 20281 19935 20315
rect 20729 20281 20763 20315
rect 21097 20281 21131 20315
rect 21741 20281 21775 20315
rect 22293 20281 22327 20315
rect 26065 20281 26099 20315
rect 27629 20281 27663 20315
rect 29101 20281 29135 20315
rect 29285 20281 29319 20315
rect 29837 20281 29871 20315
rect 31354 20281 31388 20315
rect 35218 20281 35252 20315
rect 40830 20281 40864 20315
rect 42073 20281 42107 20315
rect 43085 20281 43119 20315
rect 43177 20281 43211 20315
rect 45155 20281 45189 20315
rect 46213 20281 46247 20315
rect 46305 20281 46339 20315
rect 46857 20281 46891 20315
rect 23811 20213 23845 20247
rect 25191 20213 25225 20247
rect 30113 20213 30147 20247
rect 34161 20213 34195 20247
rect 35817 20213 35851 20247
rect 36737 20213 36771 20247
rect 40233 20213 40267 20247
rect 41429 20213 41463 20247
rect 41797 20213 41831 20247
rect 18061 20009 18095 20043
rect 18797 20009 18831 20043
rect 19533 20009 19567 20043
rect 21281 20009 21315 20043
rect 21833 20009 21867 20043
rect 26157 20009 26191 20043
rect 27721 20009 27755 20043
rect 29837 20009 29871 20043
rect 32321 20009 32355 20043
rect 33333 20009 33367 20043
rect 34897 20009 34931 20043
rect 36093 20009 36127 20043
rect 36461 20009 36495 20043
rect 36783 20009 36817 20043
rect 38485 20009 38519 20043
rect 40509 20009 40543 20043
rect 43085 20009 43119 20043
rect 45063 20009 45097 20043
rect 45753 20009 45787 20043
rect 46397 20009 46431 20043
rect 18613 19941 18647 19975
rect 23305 19941 23339 19975
rect 26709 19941 26743 19975
rect 29009 19941 29043 19975
rect 41797 19941 41831 19975
rect 41889 19941 41923 19975
rect 42441 19941 42475 19975
rect 43545 19941 43579 19975
rect 16819 19873 16853 19907
rect 17785 19873 17819 19907
rect 18337 19873 18371 19907
rect 19349 19873 19383 19907
rect 24961 19873 24995 19907
rect 29193 19873 29227 19907
rect 30757 19873 30791 19907
rect 30941 19873 30975 19907
rect 32137 19873 32171 19907
rect 33149 19873 33183 19907
rect 34437 19873 34471 19907
rect 35633 19873 35667 19907
rect 36680 19873 36714 19907
rect 38310 19873 38344 19907
rect 39313 19873 39347 19907
rect 39773 19873 39807 19907
rect 44960 19873 44994 19907
rect 45845 19873 45879 19907
rect 17693 19805 17727 19839
rect 18613 19805 18647 19839
rect 20913 19805 20947 19839
rect 23213 19805 23247 19839
rect 23489 19805 23523 19839
rect 25605 19805 25639 19839
rect 26617 19805 26651 19839
rect 26893 19805 26927 19839
rect 31033 19805 31067 19839
rect 40049 19805 40083 19839
rect 43453 19805 43487 19839
rect 43729 19805 43763 19839
rect 16911 19737 16945 19771
rect 22937 19737 22971 19771
rect 35817 19737 35851 19771
rect 39129 19737 39163 19771
rect 46075 19737 46109 19771
rect 20085 19669 20119 19703
rect 29285 19669 29319 19703
rect 34621 19669 34655 19703
rect 35265 19669 35299 19703
rect 41429 19669 41463 19703
rect 19349 19465 19383 19499
rect 22017 19465 22051 19499
rect 22293 19465 22327 19499
rect 23397 19465 23431 19499
rect 24961 19465 24995 19499
rect 25697 19465 25731 19499
rect 26065 19465 26099 19499
rect 27261 19465 27295 19499
rect 30573 19465 30607 19499
rect 30941 19465 30975 19499
rect 36093 19465 36127 19499
rect 38393 19465 38427 19499
rect 38945 19465 38979 19499
rect 39543 19465 39577 19499
rect 42349 19465 42383 19499
rect 45477 19465 45511 19499
rect 46305 19465 46339 19499
rect 16313 19397 16347 19431
rect 20269 19329 20303 19363
rect 20453 19329 20487 19363
rect 16405 19261 16439 19295
rect 16957 19261 16991 19295
rect 18337 19261 18371 19295
rect 18521 19261 18555 19295
rect 26801 19397 26835 19431
rect 39221 19397 39255 19431
rect 28273 19329 28307 19363
rect 34897 19329 34931 19363
rect 37473 19329 37507 19363
rect 39865 19329 39899 19363
rect 43637 19329 43671 19363
rect 22569 19261 22603 19295
rect 23673 19261 23707 19295
rect 24593 19261 24627 19295
rect 27721 19261 27755 19295
rect 27997 19261 28031 19295
rect 28641 19261 28675 19295
rect 29285 19261 29319 19295
rect 29929 19261 29963 19295
rect 31861 19261 31895 19295
rect 33057 19261 33091 19295
rect 36645 19261 36679 19295
rect 39440 19261 39474 19295
rect 17141 19193 17175 19227
rect 17877 19193 17911 19227
rect 20815 19193 20849 19227
rect 21649 19193 21683 19227
rect 22293 19193 22327 19227
rect 22477 19193 22511 19227
rect 26249 19193 26283 19227
rect 26341 19193 26375 19227
rect 27813 19193 27847 19227
rect 29101 19193 29135 19227
rect 31677 19193 31711 19227
rect 32873 19193 32907 19227
rect 35218 19193 35252 19227
rect 37565 19193 37599 19227
rect 38117 19193 38151 19227
rect 41429 19193 41463 19227
rect 41521 19193 41555 19227
rect 42073 19193 42107 19227
rect 42993 19193 43027 19227
rect 43085 19193 43119 19227
rect 44373 19193 44407 19227
rect 17509 19125 17543 19159
rect 18153 19125 18187 19159
rect 21373 19125 21407 19159
rect 22753 19125 22787 19159
rect 23121 19125 23155 19159
rect 24041 19125 24075 19159
rect 31493 19125 31527 19159
rect 31953 19125 31987 19159
rect 32505 19125 32539 19159
rect 33241 19125 33275 19159
rect 33609 19125 33643 19159
rect 33885 19125 33919 19159
rect 34529 19125 34563 19159
rect 35817 19125 35851 19159
rect 37289 19125 37323 19159
rect 41245 19125 41279 19159
rect 42717 19125 42751 19159
rect 43913 19125 43947 19159
rect 45017 19125 45051 19159
rect 16497 18921 16531 18955
rect 16865 18921 16899 18955
rect 17785 18921 17819 18955
rect 18613 18921 18647 18955
rect 23673 18921 23707 18955
rect 29009 18921 29043 18955
rect 34989 18921 35023 18955
rect 35357 18921 35391 18955
rect 38669 18921 38703 18955
rect 41981 18921 42015 18955
rect 42993 18921 43027 18955
rect 43959 18921 43993 18955
rect 21189 18853 21223 18887
rect 21741 18853 21775 18887
rect 23397 18853 23431 18887
rect 25605 18853 25639 18887
rect 26709 18853 26743 18887
rect 27905 18853 27939 18887
rect 29193 18853 29227 18887
rect 30573 18853 30607 18887
rect 34713 18853 34747 18887
rect 35725 18853 35759 18887
rect 37473 18853 37507 18887
rect 38025 18853 38059 18887
rect 41106 18853 41140 18887
rect 45017 18853 45051 18887
rect 45569 18853 45603 18887
rect 46489 18853 46523 18887
rect 46581 18853 46615 18887
rect 17417 18785 17451 18819
rect 19844 18785 19878 18819
rect 23121 18785 23155 18819
rect 25053 18785 25087 18819
rect 28181 18785 28215 18819
rect 29377 18785 29411 18819
rect 30757 18785 30791 18819
rect 32137 18785 32171 18819
rect 32321 18785 32355 18819
rect 34253 18785 34287 18819
rect 34529 18785 34563 18819
rect 36277 18785 36311 18819
rect 39564 18785 39598 18819
rect 40785 18785 40819 18819
rect 43856 18785 43890 18819
rect 19947 18717 19981 18751
rect 21097 18717 21131 18751
rect 26617 18717 26651 18751
rect 27261 18717 27295 18751
rect 31401 18717 31435 18751
rect 35633 18717 35667 18751
rect 37749 18717 37783 18751
rect 44925 18717 44959 18751
rect 46765 18717 46799 18751
rect 22569 18649 22603 18683
rect 28365 18649 28399 18683
rect 41705 18649 41739 18683
rect 18337 18581 18371 18615
rect 20545 18581 20579 18615
rect 26249 18581 26283 18615
rect 29469 18581 29503 18615
rect 30849 18581 30883 18615
rect 32413 18581 32447 18615
rect 36645 18581 36679 18615
rect 39635 18581 39669 18615
rect 40509 18581 40543 18615
rect 43637 18581 43671 18615
rect 17141 18377 17175 18411
rect 17509 18377 17543 18411
rect 21281 18377 21315 18411
rect 21557 18377 21591 18411
rect 22753 18377 22787 18411
rect 23121 18377 23155 18411
rect 24869 18377 24903 18411
rect 25145 18377 25179 18411
rect 25605 18377 25639 18411
rect 26709 18377 26743 18411
rect 29101 18377 29135 18411
rect 30481 18377 30515 18411
rect 31861 18377 31895 18411
rect 36277 18377 36311 18411
rect 37473 18377 37507 18411
rect 38393 18377 38427 18411
rect 41429 18377 41463 18411
rect 41705 18377 41739 18411
rect 43361 18377 43395 18411
rect 45845 18377 45879 18411
rect 18705 18309 18739 18343
rect 24593 18309 24627 18343
rect 39865 18309 39899 18343
rect 40233 18309 40267 18343
rect 45201 18309 45235 18343
rect 18153 18241 18187 18275
rect 20729 18241 20763 18275
rect 27629 18241 27663 18275
rect 29837 18241 29871 18275
rect 32505 18241 32539 18275
rect 37105 18241 37139 18275
rect 42671 18241 42705 18275
rect 43085 18241 43119 18275
rect 43545 18241 43579 18275
rect 46213 18241 46247 18275
rect 46857 18241 46891 18275
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 21741 18173 21775 18207
rect 23740 18173 23774 18207
rect 24685 18173 24719 18207
rect 28733 18173 28767 18207
rect 29285 18173 29319 18207
rect 30757 18173 30791 18207
rect 32137 18173 32171 18207
rect 32781 18173 32815 18207
rect 33517 18173 33551 18207
rect 34897 18173 34931 18207
rect 35081 18173 35115 18207
rect 35817 18173 35851 18207
rect 36461 18173 36495 18207
rect 36829 18173 36863 18207
rect 38761 18173 38795 18207
rect 38853 18173 38887 18207
rect 39313 18173 39347 18207
rect 40509 18173 40543 18207
rect 42568 18173 42602 18207
rect 18245 18105 18279 18139
rect 19717 18105 19751 18139
rect 25789 18105 25823 18139
rect 25881 18105 25915 18139
rect 26433 18105 26467 18139
rect 27353 18105 27387 18139
rect 27445 18105 27479 18139
rect 30573 18105 30607 18139
rect 31125 18105 31159 18139
rect 31953 18105 31987 18139
rect 33241 18105 33275 18139
rect 33333 18105 33367 18139
rect 35449 18105 35483 18139
rect 37841 18105 37875 18139
rect 39589 18105 39623 18139
rect 40871 18105 40905 18139
rect 43866 18105 43900 18139
rect 46305 18105 46339 18139
rect 17877 18037 17911 18071
rect 19349 18037 19383 18071
rect 19993 18037 20027 18071
rect 21925 18037 21959 18071
rect 22293 18037 22327 18071
rect 23811 18037 23845 18071
rect 24225 18037 24259 18071
rect 27077 18037 27111 18071
rect 28365 18037 28399 18071
rect 29469 18037 29503 18071
rect 31493 18037 31527 18071
rect 33609 18037 33643 18071
rect 34253 18037 34287 18071
rect 34621 18037 34655 18071
rect 44465 18037 44499 18071
rect 44925 18037 44959 18071
rect 47133 18037 47167 18071
rect 21005 17833 21039 17867
rect 26341 17833 26375 17867
rect 27537 17833 27571 17867
rect 32413 17833 32447 17867
rect 33333 17833 33367 17867
rect 34069 17833 34103 17867
rect 35633 17833 35667 17867
rect 36185 17833 36219 17867
rect 39957 17833 39991 17867
rect 46213 17833 46247 17867
rect 46489 17833 46523 17867
rect 17319 17765 17353 17799
rect 26709 17765 26743 17799
rect 27261 17765 27295 17799
rect 29193 17765 29227 17799
rect 30573 17765 30607 17799
rect 32137 17765 32171 17799
rect 39681 17765 39715 17799
rect 40850 17765 40884 17799
rect 44925 17765 44959 17799
rect 45477 17765 45511 17799
rect 16957 17697 16991 17731
rect 19533 17697 19567 17731
rect 19809 17697 19843 17731
rect 21097 17697 21131 17731
rect 21465 17697 21499 17731
rect 23397 17697 23431 17731
rect 24409 17697 24443 17731
rect 25421 17697 25455 17731
rect 28089 17697 28123 17731
rect 29377 17697 29411 17731
rect 30665 17697 30699 17731
rect 30849 17697 30883 17731
rect 32321 17697 32355 17731
rect 34529 17697 34563 17731
rect 36001 17697 36035 17731
rect 37749 17697 37783 17731
rect 38945 17697 38979 17731
rect 39405 17697 39439 17731
rect 43269 17697 43303 17731
rect 19901 17629 19935 17663
rect 26617 17629 26651 17663
rect 29653 17629 29687 17663
rect 35173 17629 35207 17663
rect 40601 17629 40635 17663
rect 44833 17629 44867 17663
rect 31585 17561 31619 17595
rect 17877 17493 17911 17527
rect 18153 17493 18187 17527
rect 18521 17493 18555 17527
rect 18889 17493 18923 17527
rect 23305 17493 23339 17527
rect 24593 17493 24627 17527
rect 25559 17493 25593 17527
rect 25881 17493 25915 17527
rect 28319 17493 28353 17527
rect 30113 17493 30147 17527
rect 30941 17493 30975 17527
rect 31953 17493 31987 17527
rect 36553 17493 36587 17527
rect 37933 17493 37967 17527
rect 41521 17493 41555 17527
rect 43499 17493 43533 17527
rect 43821 17493 43855 17527
rect 16865 17289 16899 17323
rect 17095 17289 17129 17323
rect 20361 17289 20395 17323
rect 20637 17289 20671 17323
rect 22753 17289 22787 17323
rect 23397 17289 23431 17323
rect 23949 17289 23983 17323
rect 25053 17289 25087 17323
rect 26525 17289 26559 17323
rect 28733 17289 28767 17323
rect 30665 17289 30699 17323
rect 31125 17289 31159 17323
rect 31493 17289 31527 17323
rect 34529 17289 34563 17323
rect 37749 17289 37783 17323
rect 38301 17289 38335 17323
rect 38669 17289 38703 17323
rect 39865 17289 39899 17323
rect 42625 17289 42659 17323
rect 43269 17289 43303 17323
rect 45155 17289 45189 17323
rect 17509 17221 17543 17255
rect 18705 17221 18739 17255
rect 29929 17221 29963 17255
rect 31769 17221 31803 17255
rect 32045 17221 32079 17255
rect 33701 17221 33735 17255
rect 36369 17221 36403 17255
rect 36553 17221 36587 17255
rect 42993 17221 43027 17255
rect 18153 17153 18187 17187
rect 20821 17153 20855 17187
rect 22017 17153 22051 17187
rect 27353 17153 27387 17187
rect 28365 17153 28399 17187
rect 29377 17153 29411 17187
rect 34069 17153 34103 17187
rect 34989 17153 35023 17187
rect 35909 17153 35943 17187
rect 39589 17153 39623 17187
rect 41705 17153 41739 17187
rect 43821 17153 43855 17187
rect 44833 17153 44867 17187
rect 17024 17085 17058 17119
rect 19625 17085 19659 17119
rect 22569 17085 22603 17119
rect 24133 17085 24167 17119
rect 25640 17085 25674 17119
rect 30941 17085 30975 17119
rect 31953 17085 31987 17119
rect 32229 17085 32263 17119
rect 33517 17085 33551 17119
rect 34897 17085 34931 17119
rect 35173 17085 35207 17119
rect 36461 17085 36495 17119
rect 36737 17085 36771 17119
rect 38853 17085 38887 17119
rect 39405 17085 39439 17119
rect 40544 17085 40578 17119
rect 45084 17085 45118 17119
rect 45477 17085 45511 17119
rect 46156 17085 46190 17119
rect 18245 17017 18279 17051
rect 19257 17017 19291 17051
rect 21142 17017 21176 17051
rect 24777 17017 24811 17051
rect 27066 17017 27100 17051
rect 27162 17017 27196 17051
rect 29469 17017 29503 17051
rect 30389 17017 30423 17051
rect 42026 17017 42060 17051
rect 43545 17017 43579 17051
rect 43637 17017 43671 17051
rect 46581 17017 46615 17051
rect 17877 16949 17911 16983
rect 19809 16949 19843 16983
rect 21741 16949 21775 16983
rect 23121 16949 23155 16983
rect 25513 16949 25547 16983
rect 25743 16949 25777 16983
rect 26065 16949 26099 16983
rect 26801 16949 26835 16983
rect 29009 16949 29043 16983
rect 32413 16949 32447 16983
rect 32965 16949 32999 16983
rect 33425 16949 33459 16983
rect 35357 16949 35391 16983
rect 36921 16949 36955 16983
rect 40233 16949 40267 16983
rect 40647 16949 40681 16983
rect 40969 16949 41003 16983
rect 41521 16949 41555 16983
rect 46259 16949 46293 16983
rect 16819 16745 16853 16779
rect 18797 16745 18831 16779
rect 21189 16745 21223 16779
rect 23075 16745 23109 16779
rect 26341 16745 26375 16779
rect 27721 16745 27755 16779
rect 34345 16745 34379 16779
rect 36829 16745 36863 16779
rect 37289 16745 37323 16779
rect 39129 16745 39163 16779
rect 40969 16745 41003 16779
rect 41705 16745 41739 16779
rect 44189 16745 44223 16779
rect 45109 16745 45143 16779
rect 19165 16677 19199 16711
rect 21557 16677 21591 16711
rect 24961 16677 24995 16711
rect 26893 16677 26927 16711
rect 27445 16677 27479 16711
rect 29330 16677 29364 16711
rect 35909 16677 35943 16711
rect 38162 16677 38196 16711
rect 40325 16677 40359 16711
rect 16748 16609 16782 16643
rect 17969 16609 18003 16643
rect 18153 16609 18187 16643
rect 19257 16609 19291 16643
rect 19809 16609 19843 16643
rect 22937 16609 22971 16643
rect 24593 16609 24627 16643
rect 31033 16609 31067 16643
rect 32413 16609 32447 16643
rect 32689 16609 32723 16643
rect 34161 16609 34195 16643
rect 35817 16609 35851 16643
rect 39589 16609 39623 16643
rect 40049 16609 40083 16643
rect 41188 16609 41222 16643
rect 42232 16609 42266 16643
rect 43428 16609 43462 16643
rect 44649 16609 44683 16643
rect 45753 16609 45787 16643
rect 47225 16609 47259 16643
rect 18245 16541 18279 16575
rect 19993 16541 20027 16575
rect 21465 16541 21499 16575
rect 21741 16541 21775 16575
rect 26801 16541 26835 16575
rect 29009 16541 29043 16575
rect 32505 16541 32539 16575
rect 33149 16541 33183 16575
rect 37841 16541 37875 16575
rect 20361 16473 20395 16507
rect 38761 16473 38795 16507
rect 40693 16473 40727 16507
rect 41291 16473 41325 16507
rect 43913 16473 43947 16507
rect 44833 16473 44867 16507
rect 47409 16473 47443 16507
rect 25237 16405 25271 16439
rect 28273 16405 28307 16439
rect 29929 16405 29963 16439
rect 31217 16405 31251 16439
rect 31585 16405 31619 16439
rect 31953 16405 31987 16439
rect 34989 16405 35023 16439
rect 36461 16405 36495 16439
rect 42303 16405 42337 16439
rect 43499 16405 43533 16439
rect 46121 16405 46155 16439
rect 17509 16201 17543 16235
rect 17877 16201 17911 16235
rect 19257 16201 19291 16235
rect 19717 16201 19751 16235
rect 20361 16201 20395 16235
rect 22017 16201 22051 16235
rect 24225 16201 24259 16235
rect 25605 16201 25639 16235
rect 26157 16201 26191 16235
rect 30389 16201 30423 16235
rect 30849 16201 30883 16235
rect 31677 16201 31711 16235
rect 34345 16201 34379 16235
rect 35541 16201 35575 16235
rect 35909 16201 35943 16235
rect 38853 16201 38887 16235
rect 41981 16201 42015 16235
rect 43453 16201 43487 16235
rect 44649 16201 44683 16235
rect 45569 16201 45603 16235
rect 22937 16133 22971 16167
rect 23305 16133 23339 16167
rect 27721 16133 27755 16167
rect 33425 16133 33459 16167
rect 33609 16133 33643 16167
rect 35173 16133 35207 16167
rect 39313 16133 39347 16167
rect 39589 16133 39623 16167
rect 47225 16133 47259 16167
rect 18613 16065 18647 16099
rect 20453 16065 20487 16099
rect 21741 16065 21775 16099
rect 23673 16065 23707 16099
rect 24685 16065 24719 16099
rect 26801 16065 26835 16099
rect 27077 16065 27111 16099
rect 29469 16065 29503 16099
rect 29745 16065 29779 16099
rect 31079 16065 31113 16099
rect 32873 16065 32907 16099
rect 18337 15997 18371 16031
rect 18521 15997 18555 16031
rect 22477 15997 22511 16031
rect 30976 15997 31010 16031
rect 32137 15997 32171 16031
rect 32229 15997 32263 16031
rect 32413 15997 32447 16031
rect 20774 15929 20808 15963
rect 24501 15929 24535 15963
rect 25006 15929 25040 15963
rect 26617 15929 26651 15963
rect 26893 15929 26927 15963
rect 29561 15929 29595 15963
rect 33241 15929 33275 15963
rect 40601 16065 40635 16099
rect 40877 16065 40911 16099
rect 33793 15997 33827 16031
rect 34989 15997 35023 16031
rect 36369 15997 36403 16031
rect 36921 15997 36955 16031
rect 37933 15997 37967 16031
rect 41613 15997 41647 16031
rect 42165 15997 42199 16031
rect 44281 15997 44315 16031
rect 45937 15997 45971 16031
rect 46397 15997 46431 16031
rect 36185 15929 36219 15963
rect 37105 15929 37139 15963
rect 38254 15929 38288 15963
rect 40325 15929 40359 15963
rect 40693 15929 40727 15963
rect 42073 15929 42107 15963
rect 43637 15929 43671 15963
rect 46121 15929 46155 15963
rect 16773 15861 16807 15895
rect 21373 15861 21407 15895
rect 22661 15861 22695 15895
rect 28365 15861 28399 15895
rect 28641 15861 28675 15895
rect 29101 15861 29135 15895
rect 32045 15861 32079 15895
rect 33425 15861 33459 15895
rect 33977 15861 34011 15895
rect 34713 15861 34747 15895
rect 37473 15861 37507 15895
rect 37749 15861 37783 15895
rect 20453 15657 20487 15691
rect 28917 15657 28951 15691
rect 29837 15657 29871 15691
rect 31217 15657 31251 15691
rect 31953 15657 31987 15691
rect 36921 15657 36955 15691
rect 37565 15657 37599 15691
rect 38025 15657 38059 15691
rect 38761 15657 38795 15691
rect 41153 15657 41187 15691
rect 47501 15657 47535 15691
rect 17785 15589 17819 15623
rect 19717 15589 19751 15623
rect 21189 15589 21223 15623
rect 21741 15589 21775 15623
rect 24961 15589 24995 15623
rect 26617 15589 26651 15623
rect 26709 15589 26743 15623
rect 32137 15589 32171 15623
rect 33701 15589 33735 15623
rect 40049 15589 40083 15623
rect 43545 15589 43579 15623
rect 45937 15589 45971 15623
rect 18153 15521 18187 15555
rect 18429 15521 18463 15555
rect 19844 15521 19878 15555
rect 22753 15521 22787 15555
rect 24225 15521 24259 15555
rect 24777 15521 24811 15555
rect 29101 15521 29135 15555
rect 29377 15521 29411 15555
rect 31033 15521 31067 15555
rect 31585 15521 31619 15555
rect 32781 15521 32815 15555
rect 33885 15521 33919 15555
rect 34897 15521 34931 15555
rect 35127 15521 35161 15555
rect 35633 15521 35667 15555
rect 36461 15521 36495 15555
rect 37749 15521 37783 15555
rect 38209 15521 38243 15555
rect 42257 15521 42291 15555
rect 47317 15521 47351 15555
rect 18613 15453 18647 15487
rect 21097 15453 21131 15487
rect 23397 15453 23431 15487
rect 27077 15453 27111 15487
rect 27537 15453 27571 15487
rect 35265 15453 35299 15487
rect 39957 15453 39991 15487
rect 40601 15453 40635 15487
rect 43453 15453 43487 15487
rect 45845 15453 45879 15487
rect 46489 15453 46523 15487
rect 19947 15385 19981 15419
rect 34069 15385 34103 15419
rect 34713 15385 34747 15419
rect 35062 15385 35096 15419
rect 44005 15385 44039 15419
rect 23765 15317 23799 15351
rect 25237 15317 25271 15351
rect 33241 15317 33275 15351
rect 34345 15317 34379 15351
rect 36645 15317 36679 15351
rect 42073 15317 42107 15351
rect 46765 15317 46799 15351
rect 18245 15113 18279 15147
rect 18613 15113 18647 15147
rect 19027 15113 19061 15147
rect 22753 15113 22787 15147
rect 23397 15113 23431 15147
rect 25881 15113 25915 15147
rect 26157 15113 26191 15147
rect 30205 15113 30239 15147
rect 31585 15113 31619 15147
rect 33406 15113 33440 15147
rect 34621 15113 34655 15147
rect 35173 15113 35207 15147
rect 36645 15113 36679 15147
rect 38301 15113 38335 15147
rect 39589 15113 39623 15147
rect 40233 15113 40267 15147
rect 41705 15113 41739 15147
rect 42901 15113 42935 15147
rect 45845 15113 45879 15147
rect 47317 15113 47351 15147
rect 24685 15045 24719 15079
rect 25375 15045 25409 15079
rect 27261 15045 27295 15079
rect 28733 15045 28767 15079
rect 29101 15045 29135 15079
rect 33517 15045 33551 15079
rect 35035 15045 35069 15079
rect 38669 15045 38703 15079
rect 39037 15045 39071 15079
rect 42211 15045 42245 15079
rect 43269 15045 43303 15079
rect 44005 15045 44039 15079
rect 44925 15045 44959 15079
rect 19901 14977 19935 15011
rect 21281 14977 21315 15011
rect 23765 14977 23799 15011
rect 28089 14977 28123 15011
rect 33609 14977 33643 15011
rect 35265 14977 35299 15011
rect 35909 14977 35943 15011
rect 40601 14977 40635 15011
rect 40877 14977 40911 15011
rect 43453 14977 43487 15011
rect 44373 14977 44407 15011
rect 46213 14977 46247 15011
rect 46489 14977 46523 15011
rect 18956 14909 18990 14943
rect 19349 14909 19383 14943
rect 21649 14909 21683 14943
rect 21925 14909 21959 14943
rect 22201 14909 22235 14943
rect 25272 14909 25306 14943
rect 26341 14909 26375 14943
rect 27537 14909 27571 14943
rect 28181 14909 28215 14943
rect 29285 14909 29319 14943
rect 30941 14909 30975 14943
rect 31100 14909 31134 14943
rect 32137 14909 32171 14943
rect 32229 14909 32263 14943
rect 32781 14909 32815 14943
rect 33149 14909 33183 14943
rect 34897 14909 34931 14943
rect 36277 14909 36311 14943
rect 36921 14909 36955 14943
rect 37473 14909 37507 14943
rect 38485 14909 38519 14943
rect 42108 14909 42142 14943
rect 45068 14909 45102 14943
rect 20263 14841 20297 14875
rect 23857 14841 23891 14875
rect 24409 14841 24443 14875
rect 25145 14841 25179 14875
rect 26662 14841 26696 14875
rect 29606 14841 29640 14875
rect 33241 14841 33275 14875
rect 33977 14841 34011 14875
rect 34345 14841 34379 14875
rect 35633 14841 35667 14875
rect 37657 14841 37691 14875
rect 40693 14841 40727 14875
rect 43545 14841 43579 14875
rect 46305 14841 46339 14875
rect 17601 14773 17635 14807
rect 19809 14773 19843 14807
rect 20821 14773 20855 14807
rect 21833 14773 21867 14807
rect 28319 14773 28353 14807
rect 31171 14773 31205 14807
rect 32413 14773 32447 14807
rect 37933 14773 37967 14807
rect 39957 14773 39991 14807
rect 45155 14773 45189 14807
rect 17417 14569 17451 14603
rect 20729 14569 20763 14603
rect 21925 14569 21959 14603
rect 30573 14569 30607 14603
rect 33793 14569 33827 14603
rect 34069 14569 34103 14603
rect 35541 14569 35575 14603
rect 36461 14569 36495 14603
rect 38761 14569 38795 14603
rect 40601 14569 40635 14603
rect 43177 14569 43211 14603
rect 43729 14569 43763 14603
rect 46213 14569 46247 14603
rect 20177 14501 20211 14535
rect 21097 14501 21131 14535
rect 21649 14501 21683 14535
rect 23397 14501 23431 14535
rect 24961 14501 24995 14535
rect 25513 14501 25547 14535
rect 27077 14501 27111 14535
rect 29469 14501 29503 14535
rect 29745 14501 29779 14535
rect 32873 14501 32907 14535
rect 35173 14501 35207 14535
rect 38162 14501 38196 14535
rect 39773 14501 39807 14535
rect 42625 14501 42659 14535
rect 45201 14501 45235 14535
rect 45293 14501 45327 14535
rect 45845 14501 45879 14535
rect 46489 14501 46523 14535
rect 17969 14433 18003 14467
rect 19441 14433 19475 14467
rect 28733 14433 28767 14467
rect 29193 14433 29227 14467
rect 30573 14433 30607 14467
rect 30849 14433 30883 14467
rect 33057 14433 33091 14467
rect 35081 14433 35115 14467
rect 36001 14433 36035 14467
rect 40325 14433 40359 14467
rect 41220 14433 41254 14467
rect 42200 14433 42234 14467
rect 43729 14433 43763 14467
rect 46708 14433 46742 14467
rect 17601 14365 17635 14399
rect 21005 14365 21039 14399
rect 23305 14365 23339 14399
rect 23949 14365 23983 14399
rect 24869 14365 24903 14399
rect 26709 14365 26743 14399
rect 26985 14365 27019 14399
rect 27353 14365 27387 14399
rect 33425 14365 33459 14399
rect 37841 14365 37875 14399
rect 39681 14365 39715 14399
rect 19901 14297 19935 14331
rect 28273 14229 28307 14263
rect 36185 14229 36219 14263
rect 36921 14229 36955 14263
rect 41291 14229 41325 14263
rect 41613 14229 41647 14263
rect 42303 14229 42337 14263
rect 46811 14229 46845 14263
rect 16497 14025 16531 14059
rect 17693 14025 17727 14059
rect 20913 14025 20947 14059
rect 23213 14025 23247 14059
rect 23857 14025 23891 14059
rect 25789 14025 25823 14059
rect 26341 14025 26375 14059
rect 29469 14025 29503 14059
rect 30113 14025 30147 14059
rect 31493 14025 31527 14059
rect 31769 14025 31803 14059
rect 33517 14025 33551 14059
rect 34345 14025 34379 14059
rect 34621 14025 34655 14059
rect 35357 14025 35391 14059
rect 36277 14025 36311 14059
rect 38577 14025 38611 14059
rect 39957 14025 39991 14059
rect 40647 14025 40681 14059
rect 43177 14025 43211 14059
rect 45477 14025 45511 14059
rect 46857 14025 46891 14059
rect 47225 14025 47259 14059
rect 21649 13957 21683 13991
rect 24317 13957 24351 13991
rect 25329 13957 25363 13991
rect 35035 13957 35069 13991
rect 35173 13957 35207 13991
rect 35909 13957 35943 13991
rect 37933 13957 37967 13991
rect 43453 13957 43487 13991
rect 18061 13889 18095 13923
rect 18429 13889 18463 13923
rect 21373 13889 21407 13923
rect 21833 13889 21867 13923
rect 25145 13889 25179 13923
rect 27353 13889 27387 13923
rect 30573 13889 30607 13923
rect 32873 13889 32907 13923
rect 35265 13889 35299 13923
rect 36921 13889 36955 13923
rect 38209 13889 38243 13923
rect 39681 13889 39715 13923
rect 41705 13889 41739 13923
rect 17877 13821 17911 13855
rect 19901 13821 19935 13855
rect 25329 13821 25363 13855
rect 25421 13821 25455 13855
rect 26617 13821 26651 13855
rect 28457 13821 28491 13855
rect 29285 13821 29319 13855
rect 29929 13821 29963 13855
rect 30481 13821 30515 13855
rect 32229 13821 32263 13855
rect 32321 13821 32355 13855
rect 32505 13821 32539 13855
rect 33149 13821 33183 13855
rect 33701 13821 33735 13855
rect 37013 13821 37047 13855
rect 38761 13821 38795 13855
rect 39221 13821 39255 13855
rect 40544 13821 40578 13855
rect 40969 13821 41003 13855
rect 46397 13821 46431 13855
rect 17141 13753 17175 13787
rect 17509 13753 17543 13787
rect 22195 13753 22229 13787
rect 24501 13753 24535 13787
rect 24593 13753 24627 13787
rect 26893 13753 26927 13787
rect 26985 13753 27019 13787
rect 28733 13753 28767 13787
rect 30914 13753 30948 13787
rect 34897 13753 34931 13787
rect 41797 13753 41831 13787
rect 42349 13753 42383 13787
rect 43729 13753 43763 13787
rect 43821 13753 43855 13787
rect 44373 13753 44407 13787
rect 16865 13685 16899 13719
rect 20361 13685 20395 13719
rect 22753 13685 22787 13719
rect 27813 13685 27847 13719
rect 29929 13685 29963 13719
rect 33885 13685 33919 13719
rect 37375 13685 37409 13719
rect 38945 13685 38979 13719
rect 41521 13685 41555 13719
rect 42625 13685 42659 13719
rect 44649 13685 44683 13719
rect 45201 13685 45235 13719
rect 46581 13685 46615 13719
rect 18429 13481 18463 13515
rect 19073 13481 19107 13515
rect 21051 13481 21085 13515
rect 21373 13481 21407 13515
rect 24501 13481 24535 13515
rect 29561 13481 29595 13515
rect 31217 13481 31251 13515
rect 33793 13481 33827 13515
rect 34529 13481 34563 13515
rect 35449 13481 35483 13515
rect 41705 13481 41739 13515
rect 22522 13413 22556 13447
rect 25053 13413 25087 13447
rect 25605 13413 25639 13447
rect 26709 13413 26743 13447
rect 28686 13413 28720 13447
rect 30389 13413 30423 13447
rect 32597 13413 32631 13447
rect 33149 13413 33183 13447
rect 36737 13413 36771 13447
rect 37013 13413 37047 13447
rect 40871 13413 40905 13447
rect 43821 13413 43855 13447
rect 45385 13413 45419 13447
rect 46765 13413 46799 13447
rect 17969 13345 18003 13379
rect 20821 13345 20855 13379
rect 23121 13345 23155 13379
rect 29285 13345 29319 13379
rect 32781 13345 32815 13379
rect 34621 13345 34655 13379
rect 34805 13345 34839 13379
rect 36001 13345 36035 13379
rect 36553 13345 36587 13379
rect 37933 13345 37967 13379
rect 38393 13345 38427 13379
rect 39497 13345 39531 13379
rect 41429 13345 41463 13379
rect 42324 13345 42358 13379
rect 47133 13345 47167 13379
rect 16129 13277 16163 13311
rect 16497 13277 16531 13311
rect 19349 13277 19383 13311
rect 22201 13277 22235 13311
rect 24961 13277 24995 13311
rect 26617 13277 26651 13311
rect 26893 13277 26927 13311
rect 28365 13277 28399 13311
rect 30297 13277 30331 13311
rect 35173 13277 35207 13311
rect 38669 13277 38703 13311
rect 38945 13277 38979 13311
rect 40509 13277 40543 13311
rect 43729 13277 43763 13311
rect 44373 13277 44407 13311
rect 45293 13277 45327 13311
rect 30849 13209 30883 13243
rect 45845 13209 45879 13243
rect 18705 13141 18739 13175
rect 21925 13141 21959 13175
rect 26341 13141 26375 13175
rect 27721 13141 27755 13175
rect 33517 13141 33551 13175
rect 39681 13141 39715 13175
rect 40417 13141 40451 13175
rect 42165 13141 42199 13175
rect 42395 13141 42429 13175
rect 46305 13141 46339 13175
rect 15853 12937 15887 12971
rect 17785 12937 17819 12971
rect 18245 12937 18279 12971
rect 20913 12937 20947 12971
rect 22845 12937 22879 12971
rect 24593 12937 24627 12971
rect 25145 12937 25179 12971
rect 26985 12937 27019 12971
rect 30665 12937 30699 12971
rect 32229 12937 32263 12971
rect 33609 12937 33643 12971
rect 37289 12937 37323 12971
rect 39589 12937 39623 12971
rect 43177 12937 43211 12971
rect 47133 12937 47167 12971
rect 32505 12869 32539 12903
rect 33149 12869 33183 12903
rect 36277 12869 36311 12903
rect 39865 12869 39899 12903
rect 40325 12869 40359 12903
rect 18797 12801 18831 12835
rect 22385 12801 22419 12835
rect 23811 12801 23845 12835
rect 26525 12801 26559 12835
rect 28365 12801 28399 12835
rect 29377 12801 29411 12835
rect 35909 12801 35943 12835
rect 38669 12801 38703 12835
rect 41521 12801 41555 12835
rect 42165 12801 42199 12835
rect 42809 12801 42843 12835
rect 44005 12801 44039 12835
rect 44649 12801 44683 12835
rect 46489 12801 46523 12835
rect 21741 12733 21775 12767
rect 22109 12733 22143 12767
rect 22293 12733 22327 12767
rect 23724 12733 23758 12767
rect 24133 12733 24167 12767
rect 24685 12733 24719 12767
rect 25881 12733 25915 12767
rect 26249 12733 26283 12767
rect 26433 12733 26467 12767
rect 27537 12733 27571 12767
rect 27905 12733 27939 12767
rect 28089 12733 28123 12767
rect 30916 12733 30950 12767
rect 32321 12733 32355 12767
rect 33333 12733 33367 12767
rect 33517 12733 33551 12767
rect 35081 12733 35115 12767
rect 35265 12733 35299 12767
rect 36461 12733 36495 12767
rect 36921 12733 36955 12767
rect 37473 12733 37507 12767
rect 40509 12733 40543 12767
rect 40969 12733 41003 12767
rect 16589 12665 16623 12699
rect 29469 12665 29503 12699
rect 30021 12665 30055 12699
rect 34161 12665 34195 12699
rect 34713 12665 34747 12699
rect 35633 12665 35667 12699
rect 37933 12665 37967 12699
rect 38990 12665 39024 12699
rect 42257 12665 42291 12699
rect 43453 12665 43487 12699
rect 43729 12665 43763 12699
rect 43821 12665 43855 12699
rect 46213 12665 46247 12699
rect 46305 12665 46339 12699
rect 16221 12597 16255 12631
rect 16957 12597 16991 12631
rect 18705 12597 18739 12631
rect 19165 12597 19199 12631
rect 19717 12597 19751 12631
rect 24869 12597 24903 12631
rect 28641 12597 28675 12631
rect 29009 12597 29043 12631
rect 30297 12597 30331 12631
rect 30987 12597 31021 12631
rect 31309 12597 31343 12631
rect 32781 12597 32815 12631
rect 36645 12597 36679 12631
rect 37657 12597 37691 12631
rect 38485 12597 38519 12631
rect 40601 12597 40635 12631
rect 41981 12597 42015 12631
rect 45293 12597 45327 12631
rect 45937 12597 45971 12631
rect 18429 12393 18463 12427
rect 19349 12393 19383 12427
rect 22201 12393 22235 12427
rect 24777 12393 24811 12427
rect 26065 12393 26099 12427
rect 26709 12393 26743 12427
rect 28365 12393 28399 12427
rect 29377 12393 29411 12427
rect 33333 12393 33367 12427
rect 34713 12393 34747 12427
rect 35173 12393 35207 12427
rect 36185 12393 36219 12427
rect 40325 12393 40359 12427
rect 41337 12393 41371 12427
rect 42303 12393 42337 12427
rect 42625 12393 42659 12427
rect 43821 12393 43855 12427
rect 45201 12393 45235 12427
rect 21097 12325 21131 12359
rect 23121 12325 23155 12359
rect 27261 12325 27295 12359
rect 27813 12325 27847 12359
rect 30113 12325 30147 12359
rect 30665 12325 30699 12359
rect 32505 12325 32539 12359
rect 33885 12325 33919 12359
rect 38162 12325 38196 12359
rect 40779 12325 40813 12359
rect 45477 12325 45511 12359
rect 46029 12325 46063 12359
rect 46857 12325 46891 12359
rect 17141 12257 17175 12291
rect 18981 12257 19015 12291
rect 24593 12257 24627 12291
rect 25053 12257 25087 12291
rect 28676 12257 28710 12291
rect 32689 12257 32723 12291
rect 34069 12257 34103 12291
rect 35633 12257 35667 12291
rect 36645 12257 36679 12291
rect 38761 12257 38795 12291
rect 42200 12257 42234 12291
rect 43396 12257 43430 12291
rect 46949 12257 46983 12291
rect 21005 12189 21039 12223
rect 21281 12189 21315 12223
rect 23029 12189 23063 12223
rect 27169 12189 27203 12223
rect 28779 12189 28813 12223
rect 30021 12189 30055 12223
rect 33057 12189 33091 12223
rect 33793 12189 33827 12223
rect 34437 12189 34471 12223
rect 37841 12189 37875 12223
rect 40417 12189 40451 12223
rect 45385 12189 45419 12223
rect 23581 12121 23615 12155
rect 36829 12121 36863 12155
rect 19901 12053 19935 12087
rect 24409 12053 24443 12087
rect 25513 12053 25547 12087
rect 35541 12053 35575 12087
rect 35817 12053 35851 12087
rect 37565 12053 37599 12087
rect 39129 12053 39163 12087
rect 43499 12053 43533 12087
rect 44189 12053 44223 12087
rect 18521 11849 18555 11883
rect 20177 11849 20211 11883
rect 20545 11849 20579 11883
rect 23029 11849 23063 11883
rect 23397 11849 23431 11883
rect 26249 11849 26283 11883
rect 26709 11849 26743 11883
rect 28181 11849 28215 11883
rect 29101 11849 29135 11883
rect 34161 11849 34195 11883
rect 36093 11849 36127 11883
rect 36645 11849 36679 11883
rect 40325 11849 40359 11883
rect 42073 11849 42107 11883
rect 43269 11849 43303 11883
rect 43545 11849 43579 11883
rect 45385 11849 45419 11883
rect 46857 11849 46891 11883
rect 19901 11781 19935 11815
rect 24961 11781 24995 11815
rect 25053 11781 25087 11815
rect 41705 11781 41739 11815
rect 18613 11713 18647 11747
rect 21189 11713 21223 11747
rect 23765 11713 23799 11747
rect 24409 11713 24443 11747
rect 20428 11645 20462 11679
rect 21557 11645 21591 11679
rect 21833 11645 21867 11679
rect 22109 11645 22143 11679
rect 18934 11577 18968 11611
rect 23857 11577 23891 11611
rect 25973 11713 26007 11747
rect 27169 11713 27203 11747
rect 30297 11713 30331 11747
rect 39957 11713 39991 11747
rect 42257 11713 42291 11747
rect 42533 11713 42567 11747
rect 29745 11645 29779 11679
rect 31493 11645 31527 11679
rect 31769 11645 31803 11679
rect 32597 11645 32631 11679
rect 33149 11645 33183 11679
rect 33793 11645 33827 11679
rect 35265 11645 35299 11679
rect 35541 11645 35575 11679
rect 37105 11645 37139 11679
rect 37473 11645 37507 11679
rect 37749 11645 37783 11679
rect 38853 11645 38887 11679
rect 39405 11645 39439 11679
rect 40509 11645 40543 11679
rect 40969 11645 41003 11679
rect 25329 11577 25363 11611
rect 25421 11577 25455 11611
rect 26893 11577 26927 11611
rect 26985 11577 27019 11611
rect 27813 11577 27847 11611
rect 30021 11577 30055 11611
rect 30113 11577 30147 11611
rect 31585 11577 31619 11611
rect 32137 11577 32171 11611
rect 32965 11577 32999 11611
rect 33517 11577 33551 11611
rect 35725 11577 35759 11611
rect 37933 11577 37967 11611
rect 39589 11577 39623 11611
rect 42349 11577 42383 11611
rect 43821 11577 43855 11611
rect 43913 11577 43947 11611
rect 44465 11577 44499 11611
rect 45661 11577 45695 11611
rect 17233 11509 17267 11543
rect 19533 11509 19567 11543
rect 21741 11509 21775 11543
rect 24685 11509 24719 11543
rect 24961 11509 24995 11543
rect 28641 11509 28675 11543
rect 30941 11509 30975 11543
rect 34713 11509 34747 11543
rect 38209 11509 38243 11543
rect 38669 11509 38703 11543
rect 40601 11509 40635 11543
rect 18613 11305 18647 11339
rect 20453 11305 20487 11339
rect 21465 11305 21499 11339
rect 23029 11305 23063 11339
rect 23535 11305 23569 11339
rect 24961 11305 24995 11339
rect 28733 11305 28767 11339
rect 29929 11305 29963 11339
rect 31585 11305 31619 11339
rect 32505 11305 32539 11339
rect 33885 11305 33919 11339
rect 36737 11305 36771 11339
rect 37289 11305 37323 11339
rect 37933 11305 37967 11339
rect 40233 11305 40267 11339
rect 42165 11305 42199 11339
rect 19257 11237 19291 11271
rect 21970 11237 22004 11271
rect 27261 11237 27295 11271
rect 27813 11237 27847 11271
rect 32873 11237 32907 11271
rect 33425 11237 33459 11271
rect 38761 11237 38795 11271
rect 41014 11237 41048 11271
rect 44005 11237 44039 11271
rect 18096 11169 18130 11203
rect 19809 11169 19843 11203
rect 21097 11169 21131 11203
rect 22569 11169 22603 11203
rect 23432 11169 23466 11203
rect 28641 11169 28675 11203
rect 29193 11169 29227 11203
rect 30481 11169 30515 11203
rect 30665 11169 30699 11203
rect 33057 11169 33091 11203
rect 34989 11169 35023 11203
rect 35541 11169 35575 11203
rect 36553 11169 36587 11203
rect 45512 11169 45546 11203
rect 19165 11101 19199 11135
rect 21649 11101 21683 11135
rect 24593 11101 24627 11135
rect 27169 11101 27203 11135
rect 30941 11101 30975 11135
rect 35725 11101 35759 11135
rect 38669 11101 38703 11135
rect 40693 11101 40727 11135
rect 43913 11101 43947 11135
rect 44557 11101 44591 11135
rect 39221 11033 39255 11067
rect 18199 10965 18233 10999
rect 23857 10965 23891 10999
rect 25513 10965 25547 10999
rect 26801 10965 26835 10999
rect 28089 10965 28123 10999
rect 40509 10965 40543 10999
rect 41613 10965 41647 10999
rect 45615 10965 45649 10999
rect 16221 10761 16255 10795
rect 17095 10761 17129 10795
rect 19165 10761 19199 10795
rect 20821 10761 20855 10795
rect 21281 10761 21315 10795
rect 21557 10761 21591 10795
rect 23397 10761 23431 10795
rect 26479 10761 26513 10795
rect 26893 10761 26927 10795
rect 29101 10761 29135 10795
rect 31309 10761 31343 10795
rect 33425 10761 33459 10795
rect 33793 10761 33827 10795
rect 37289 10761 37323 10795
rect 40325 10761 40359 10795
rect 40785 10761 40819 10795
rect 42441 10761 42475 10795
rect 43453 10761 43487 10795
rect 44925 10761 44959 10795
rect 45477 10761 45511 10795
rect 16773 10693 16807 10727
rect 20085 10693 20119 10727
rect 29561 10693 29595 10727
rect 35081 10693 35115 10727
rect 41797 10693 41831 10727
rect 43821 10693 43855 10727
rect 44557 10693 44591 10727
rect 17877 10625 17911 10659
rect 19533 10625 19567 10659
rect 21741 10625 21775 10659
rect 24593 10625 24627 10659
rect 32137 10625 32171 10659
rect 34621 10625 34655 10659
rect 36093 10625 36127 10659
rect 37841 10625 37875 10659
rect 40877 10625 40911 10659
rect 16405 10557 16439 10591
rect 17024 10557 17058 10591
rect 18464 10557 18498 10591
rect 22937 10557 22971 10591
rect 25513 10557 25547 10591
rect 26157 10557 26191 10591
rect 26376 10557 26410 10591
rect 27445 10557 27479 10591
rect 29377 10557 29411 10591
rect 30389 10557 30423 10591
rect 31677 10557 31711 10591
rect 34897 10557 34931 10591
rect 35357 10557 35391 10591
rect 39129 10557 39163 10591
rect 42660 10557 42694 10591
rect 45937 10557 45971 10591
rect 46765 10557 46799 10591
rect 19625 10489 19659 10523
rect 22062 10489 22096 10523
rect 24041 10489 24075 10523
rect 24409 10489 24443 10523
rect 24914 10489 24948 10523
rect 27261 10489 27295 10523
rect 27766 10489 27800 10523
rect 30297 10489 30331 10523
rect 30710 10489 30744 10523
rect 31953 10489 31987 10523
rect 32458 10489 32492 10523
rect 35909 10489 35943 10523
rect 36414 10489 36448 10523
rect 37657 10489 37691 10523
rect 38162 10489 38196 10523
rect 41198 10489 41232 10523
rect 44005 10489 44039 10523
rect 44097 10489 44131 10523
rect 46121 10489 46155 10523
rect 17509 10421 17543 10455
rect 18245 10421 18279 10455
rect 18567 10421 18601 10455
rect 20453 10421 20487 10455
rect 22661 10421 22695 10455
rect 25789 10421 25823 10455
rect 28365 10421 28399 10455
rect 28641 10421 28675 10455
rect 29929 10421 29963 10455
rect 33057 10421 33091 10455
rect 34345 10421 34379 10455
rect 37013 10421 37047 10455
rect 38761 10421 38795 10455
rect 39497 10421 39531 10455
rect 39957 10421 39991 10455
rect 42763 10421 42797 10455
rect 19809 10217 19843 10251
rect 20085 10217 20119 10251
rect 21649 10217 21683 10251
rect 22569 10217 22603 10251
rect 23259 10217 23293 10251
rect 24409 10217 24443 10251
rect 25145 10217 25179 10251
rect 26663 10217 26697 10251
rect 28457 10217 28491 10251
rect 30021 10217 30055 10251
rect 30481 10217 30515 10251
rect 31217 10217 31251 10251
rect 32321 10217 32355 10251
rect 36093 10217 36127 10251
rect 37933 10217 37967 10251
rect 40233 10217 40267 10251
rect 41153 10217 41187 10251
rect 43729 10217 43763 10251
rect 47685 10217 47719 10251
rect 27858 10149 27892 10183
rect 32873 10149 32907 10183
rect 38761 10149 38795 10183
rect 41797 10149 41831 10183
rect 41889 10149 41923 10183
rect 42441 10149 42475 10183
rect 44005 10149 44039 10183
rect 17509 10081 17543 10115
rect 19349 10081 19383 10115
rect 21557 10081 21591 10115
rect 22109 10081 22143 10115
rect 23156 10081 23190 10115
rect 24133 10081 24167 10115
rect 24593 10081 24627 10115
rect 26560 10081 26594 10115
rect 27537 10081 27571 10115
rect 30389 10081 30423 10115
rect 30757 10081 30791 10115
rect 33057 10081 33091 10115
rect 35173 10081 35207 10115
rect 35449 10081 35483 10115
rect 36461 10081 36495 10115
rect 40141 10081 40175 10115
rect 40693 10081 40727 10115
rect 46029 10081 46063 10115
rect 47501 10081 47535 10115
rect 17877 10013 17911 10047
rect 35633 10013 35667 10047
rect 38669 10013 38703 10047
rect 43913 10013 43947 10047
rect 45937 10013 45971 10047
rect 39221 9945 39255 9979
rect 44465 9945 44499 9979
rect 23857 9877 23891 9911
rect 27169 9877 27203 9911
rect 29285 9877 29319 9911
rect 33149 9877 33183 9911
rect 36645 9877 36679 9911
rect 16773 9673 16807 9707
rect 19395 9673 19429 9707
rect 22017 9673 22051 9707
rect 22477 9673 22511 9707
rect 25697 9673 25731 9707
rect 29101 9673 29135 9707
rect 30389 9673 30423 9707
rect 30665 9673 30699 9707
rect 32413 9673 32447 9707
rect 32689 9673 32723 9707
rect 33333 9673 33367 9707
rect 33701 9673 33735 9707
rect 34713 9673 34747 9707
rect 37013 9673 37047 9707
rect 38485 9673 38519 9707
rect 38715 9673 38749 9707
rect 39037 9673 39071 9707
rect 40647 9673 40681 9707
rect 40969 9673 41003 9707
rect 41797 9673 41831 9707
rect 43545 9673 43579 9707
rect 45937 9673 45971 9707
rect 47501 9673 47535 9707
rect 31033 9605 31067 9639
rect 35173 9605 35207 9639
rect 35725 9605 35759 9639
rect 40141 9605 40175 9639
rect 43085 9605 43119 9639
rect 45569 9605 45603 9639
rect 20269 9537 20303 9571
rect 35817 9537 35851 9571
rect 39405 9537 39439 9571
rect 42533 9537 42567 9571
rect 44373 9537 44407 9571
rect 45017 9537 45051 9571
rect 46213 9537 46247 9571
rect 47133 9537 47167 9571
rect 17509 9469 17543 9503
rect 18312 9469 18346 9503
rect 19324 9469 19358 9503
rect 20177 9469 20211 9503
rect 20361 9469 20395 9503
rect 22636 9469 22670 9503
rect 23489 9469 23523 9503
rect 23765 9469 23799 9503
rect 24225 9469 24259 9503
rect 25789 9469 25823 9503
rect 26249 9469 26283 9503
rect 27905 9469 27939 9503
rect 28181 9469 28215 9503
rect 29285 9469 29319 9503
rect 29745 9469 29779 9503
rect 30849 9469 30883 9503
rect 31309 9469 31343 9503
rect 31861 9469 31895 9503
rect 32873 9469 32907 9503
rect 37565 9469 37599 9503
rect 38025 9469 38059 9503
rect 38612 9469 38646 9503
rect 40544 9469 40578 9503
rect 41337 9469 41371 9503
rect 26525 9401 26559 9435
rect 27169 9401 27203 9435
rect 36138 9401 36172 9435
rect 42625 9401 42659 9435
rect 43821 9401 43855 9435
rect 44097 9401 44131 9435
rect 44189 9401 44223 9435
rect 46305 9401 46339 9435
rect 46857 9401 46891 9435
rect 17141 9333 17175 9367
rect 18383 9333 18417 9367
rect 18797 9333 18831 9367
rect 19809 9333 19843 9367
rect 21557 9333 21591 9367
rect 22707 9333 22741 9367
rect 23121 9333 23155 9367
rect 23857 9333 23891 9367
rect 24869 9333 24903 9367
rect 27445 9333 27479 9367
rect 27721 9333 27755 9367
rect 29561 9333 29595 9367
rect 32045 9333 32079 9367
rect 33057 9333 33091 9367
rect 36737 9333 36771 9367
rect 37749 9333 37783 9367
rect 42257 9333 42291 9367
rect 17601 9129 17635 9163
rect 18843 9129 18877 9163
rect 19901 9129 19935 9163
rect 24225 9129 24259 9163
rect 25789 9129 25823 9163
rect 26249 9129 26283 9163
rect 27813 9129 27847 9163
rect 28181 9129 28215 9163
rect 30619 9129 30653 9163
rect 35541 9129 35575 9163
rect 35817 9129 35851 9163
rect 38117 9129 38151 9163
rect 39865 9129 39899 9163
rect 41613 9129 41647 9163
rect 42717 9129 42751 9163
rect 44465 9129 44499 9163
rect 47363 9129 47397 9163
rect 26887 9061 26921 9095
rect 41889 9061 41923 9095
rect 42441 9061 42475 9095
rect 43545 9061 43579 9095
rect 45845 9061 45879 9095
rect 18705 8993 18739 9027
rect 19717 8993 19751 9027
rect 21005 8993 21039 9027
rect 23213 8993 23247 9027
rect 24720 8993 24754 9027
rect 28917 8993 28951 9027
rect 29377 8993 29411 9027
rect 30548 8993 30582 9027
rect 32597 8993 32631 9027
rect 33057 8993 33091 9027
rect 34437 8993 34471 9027
rect 34989 8993 35023 9027
rect 36093 8993 36127 9027
rect 36553 8993 36587 9027
rect 47225 8993 47259 9027
rect 20913 8925 20947 8959
rect 23857 8925 23891 8959
rect 26525 8925 26559 8959
rect 29653 8925 29687 8959
rect 29929 8925 29963 8959
rect 33333 8925 33367 8959
rect 35173 8925 35207 8959
rect 36829 8925 36863 8959
rect 37749 8925 37783 8959
rect 39497 8925 39531 8959
rect 41797 8925 41831 8959
rect 43453 8925 43487 8959
rect 43729 8925 43763 8959
rect 45753 8925 45787 8959
rect 46029 8925 46063 8959
rect 40417 8857 40451 8891
rect 24823 8789 24857 8823
rect 27445 8789 27479 8823
rect 33701 8789 33735 8823
rect 38669 8789 38703 8823
rect 20085 8585 20119 8619
rect 21649 8585 21683 8619
rect 22477 8585 22511 8619
rect 22753 8585 22787 8619
rect 24685 8585 24719 8619
rect 24961 8585 24995 8619
rect 27353 8585 27387 8619
rect 27675 8585 27709 8619
rect 28733 8585 28767 8619
rect 30849 8585 30883 8619
rect 32597 8585 32631 8619
rect 33057 8585 33091 8619
rect 34437 8585 34471 8619
rect 38117 8585 38151 8619
rect 40969 8585 41003 8619
rect 42441 8585 42475 8619
rect 43637 8585 43671 8619
rect 45385 8585 45419 8619
rect 23029 8517 23063 8551
rect 28273 8517 28307 8551
rect 31217 8517 31251 8551
rect 42257 8517 42291 8551
rect 43085 8517 43119 8551
rect 18613 8449 18647 8483
rect 19809 8449 19843 8483
rect 21005 8449 21039 8483
rect 23765 8449 23799 8483
rect 29561 8449 29595 8483
rect 31401 8449 31435 8483
rect 31677 8449 31711 8483
rect 35633 8449 35667 8483
rect 40233 8449 40267 8483
rect 42165 8449 42199 8483
rect 45753 8449 45787 8483
rect 22569 8381 22603 8415
rect 27604 8381 27638 8415
rect 33241 8381 33275 8415
rect 33793 8381 33827 8415
rect 34897 8381 34931 8415
rect 35449 8381 35483 8415
rect 36737 8381 36771 8415
rect 37197 8381 37231 8415
rect 38669 8381 38703 8415
rect 41245 8381 41279 8415
rect 42257 8381 42291 8415
rect 43212 8381 43246 8415
rect 43315 8381 43349 8415
rect 44281 8381 44315 8415
rect 46213 8381 46247 8415
rect 19165 8313 19199 8347
rect 19257 8313 19291 8347
rect 20729 8313 20763 8347
rect 20821 8313 20855 8347
rect 23397 8313 23431 8347
rect 24086 8313 24120 8347
rect 26065 8313 26099 8347
rect 26157 8313 26191 8347
rect 26709 8313 26743 8347
rect 29101 8313 29135 8347
rect 29923 8313 29957 8347
rect 31493 8313 31527 8347
rect 33977 8313 34011 8347
rect 39031 8313 39065 8347
rect 41521 8313 41555 8347
rect 41613 8313 41647 8347
rect 44005 8313 44039 8347
rect 46121 8313 46155 8347
rect 18981 8245 19015 8279
rect 20545 8245 20579 8279
rect 25881 8245 25915 8279
rect 27077 8245 27111 8279
rect 30481 8245 30515 8279
rect 36093 8245 36127 8279
rect 36553 8245 36587 8279
rect 37013 8245 37047 8279
rect 37841 8245 37875 8279
rect 38577 8245 38611 8279
rect 39589 8245 39623 8279
rect 39865 8245 39899 8279
rect 44465 8245 44499 8279
rect 47225 8245 47259 8279
rect 23673 8041 23707 8075
rect 24225 8041 24259 8075
rect 27629 8041 27663 8075
rect 32873 8041 32907 8075
rect 34897 8041 34931 8075
rect 36369 8041 36403 8075
rect 36829 8041 36863 8075
rect 38761 8041 38795 8075
rect 44281 8041 44315 8075
rect 46535 8041 46569 8075
rect 21097 7973 21131 8007
rect 24961 7973 24995 8007
rect 25053 7973 25087 8007
rect 25605 7973 25639 8007
rect 26709 7973 26743 8007
rect 28273 7973 28307 8007
rect 30015 7973 30049 8007
rect 33695 7973 33729 8007
rect 35443 7973 35477 8007
rect 39767 7973 39801 8007
rect 45017 7973 45051 8007
rect 45569 7973 45603 8007
rect 46213 7973 46247 8007
rect 19476 7905 19510 7939
rect 23857 7905 23891 7939
rect 29653 7905 29687 7939
rect 32388 7905 32422 7939
rect 34253 7905 34287 7939
rect 35081 7905 35115 7939
rect 38368 7905 38402 7939
rect 41705 7905 41739 7939
rect 42349 7905 42383 7939
rect 43821 7905 43855 7939
rect 46432 7905 46466 7939
rect 47409 7905 47443 7939
rect 21005 7837 21039 7871
rect 26617 7837 26651 7871
rect 26893 7837 26927 7871
rect 28181 7837 28215 7871
rect 28457 7837 28491 7871
rect 33333 7837 33367 7871
rect 34621 7837 34655 7871
rect 39405 7837 39439 7871
rect 41521 7837 41555 7871
rect 44925 7837 44959 7871
rect 19165 7769 19199 7803
rect 20729 7769 20763 7803
rect 21557 7769 21591 7803
rect 32459 7769 32493 7803
rect 38439 7769 38473 7803
rect 40325 7769 40359 7803
rect 44005 7769 44039 7803
rect 19579 7701 19613 7735
rect 26065 7701 26099 7735
rect 30573 7701 30607 7735
rect 30849 7701 30883 7735
rect 31309 7701 31343 7735
rect 36001 7701 36035 7735
rect 44649 7701 44683 7735
rect 47547 7701 47581 7735
rect 19441 7497 19475 7531
rect 22661 7497 22695 7531
rect 23305 7497 23339 7531
rect 24133 7497 24167 7531
rect 25237 7497 25271 7531
rect 27859 7497 27893 7531
rect 28181 7497 28215 7531
rect 29653 7497 29687 7531
rect 32229 7497 32263 7531
rect 32597 7497 32631 7531
rect 33793 7497 33827 7531
rect 35173 7497 35207 7531
rect 37013 7497 37047 7531
rect 38485 7497 38519 7531
rect 38761 7497 38795 7531
rect 39129 7497 39163 7531
rect 42533 7497 42567 7531
rect 43223 7497 43257 7531
rect 43821 7497 43855 7531
rect 44373 7497 44407 7531
rect 45569 7497 45603 7531
rect 45937 7497 45971 7531
rect 47133 7497 47167 7531
rect 30297 7429 30331 7463
rect 42901 7429 42935 7463
rect 47501 7429 47535 7463
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 21097 7361 21131 7395
rect 21373 7361 21407 7395
rect 24961 7361 24995 7395
rect 29883 7361 29917 7395
rect 30849 7361 30883 7395
rect 31493 7361 31527 7395
rect 33425 7361 33459 7395
rect 34069 7361 34103 7395
rect 35633 7361 35667 7395
rect 36553 7361 36587 7395
rect 37565 7361 37599 7395
rect 41521 7361 41555 7395
rect 45201 7361 45235 7395
rect 46489 7361 46523 7395
rect 19809 7293 19843 7327
rect 24317 7293 24351 7327
rect 26249 7293 26283 7327
rect 27756 7293 27790 7327
rect 28549 7293 28583 7327
rect 29780 7293 29814 7327
rect 32689 7293 32723 7327
rect 33149 7293 33183 7327
rect 39348 7293 39382 7327
rect 40141 7293 40175 7327
rect 40576 7293 40610 7327
rect 41429 7293 41463 7327
rect 42165 7293 42199 7327
rect 43120 7293 43154 7327
rect 21465 7225 21499 7259
rect 22017 7225 22051 7259
rect 29009 7225 29043 7259
rect 30941 7225 30975 7259
rect 34713 7225 34747 7259
rect 35725 7225 35759 7259
rect 36277 7225 36311 7259
rect 37473 7225 37507 7259
rect 37927 7225 37961 7259
rect 39451 7225 39485 7259
rect 44557 7225 44591 7259
rect 44649 7225 44683 7259
rect 46213 7225 46247 7259
rect 46305 7225 46339 7259
rect 22385 7157 22419 7191
rect 24501 7157 24535 7191
rect 25973 7157 26007 7191
rect 26433 7157 26467 7191
rect 27169 7157 27203 7191
rect 30573 7157 30607 7191
rect 39773 7157 39807 7191
rect 40647 7157 40681 7191
rect 41061 7157 41095 7191
rect 26709 6953 26743 6987
rect 29837 6953 29871 6987
rect 32689 6953 32723 6987
rect 35081 6953 35115 6987
rect 42257 6953 42291 6987
rect 46627 6953 46661 6987
rect 19809 6885 19843 6919
rect 21097 6885 21131 6919
rect 21649 6885 21683 6919
rect 22839 6885 22873 6919
rect 27445 6885 27479 6919
rect 29009 6885 29043 6919
rect 30665 6885 30699 6919
rect 35357 6885 35391 6919
rect 35633 6885 35667 6919
rect 35725 6885 35759 6919
rect 39037 6885 39071 6919
rect 39129 6885 39163 6919
rect 40601 6885 40635 6919
rect 40693 6885 40727 6919
rect 43545 6885 43579 6919
rect 45109 6885 45143 6919
rect 45661 6885 45695 6919
rect 19165 6817 19199 6851
rect 24292 6817 24326 6851
rect 25421 6817 25455 6851
rect 32965 6817 32999 6851
rect 33977 6817 34011 6851
rect 34529 6817 34563 6851
rect 37749 6817 37783 6851
rect 42073 6817 42107 6851
rect 46213 6817 46247 6851
rect 46524 6817 46558 6851
rect 21005 6749 21039 6783
rect 22477 6749 22511 6783
rect 27353 6749 27387 6783
rect 28917 6749 28951 6783
rect 30573 6749 30607 6783
rect 34713 6749 34747 6783
rect 36277 6749 36311 6783
rect 40877 6749 40911 6783
rect 43453 6749 43487 6783
rect 44097 6749 44131 6783
rect 45017 6749 45051 6783
rect 27905 6681 27939 6715
rect 29469 6681 29503 6715
rect 31125 6681 31159 6715
rect 39589 6681 39623 6715
rect 19349 6613 19383 6647
rect 22385 6613 22419 6647
rect 23397 6613 23431 6647
rect 23765 6613 23799 6647
rect 24363 6613 24397 6647
rect 25329 6613 25363 6647
rect 25605 6613 25639 6647
rect 27169 6613 27203 6647
rect 28641 6613 28675 6647
rect 33149 6613 33183 6647
rect 36553 6613 36587 6647
rect 37933 6613 37967 6647
rect 38485 6613 38519 6647
rect 41613 6613 41647 6647
rect 44465 6613 44499 6647
rect 19257 6409 19291 6443
rect 20177 6409 20211 6443
rect 21005 6409 21039 6443
rect 26249 6409 26283 6443
rect 27905 6409 27939 6443
rect 28457 6409 28491 6443
rect 28917 6409 28951 6443
rect 30389 6409 30423 6443
rect 31769 6409 31803 6443
rect 32965 6409 32999 6443
rect 34621 6409 34655 6443
rect 35035 6409 35069 6443
rect 38301 6409 38335 6443
rect 42165 6409 42199 6443
rect 42625 6409 42659 6443
rect 44557 6409 44591 6443
rect 45201 6409 45235 6443
rect 47133 6409 47167 6443
rect 37749 6341 37783 6375
rect 44925 6341 44959 6375
rect 22569 6273 22603 6307
rect 23765 6273 23799 6307
rect 24409 6273 24443 6307
rect 25329 6273 25363 6307
rect 25605 6273 25639 6307
rect 26893 6273 26927 6307
rect 27261 6273 27295 6307
rect 32689 6273 32723 6307
rect 41061 6273 41095 6307
rect 41521 6273 41555 6307
rect 43269 6273 43303 6307
rect 43913 6273 43947 6307
rect 19625 6205 19659 6239
rect 19809 6205 19843 6239
rect 21925 6205 21959 6239
rect 22293 6205 22327 6239
rect 22477 6205 22511 6239
rect 29285 6205 29319 6239
rect 30573 6205 30607 6239
rect 32137 6205 32171 6239
rect 33425 6205 33459 6239
rect 33701 6205 33735 6239
rect 34964 6205 34998 6239
rect 38485 6205 38519 6239
rect 38945 6205 38979 6239
rect 39589 6205 39623 6239
rect 44741 6205 44775 6239
rect 46213 6205 46247 6239
rect 23489 6137 23523 6171
rect 23857 6137 23891 6171
rect 25421 6137 25455 6171
rect 26617 6137 26651 6171
rect 26985 6137 27019 6171
rect 30894 6137 30928 6171
rect 33977 6137 34011 6171
rect 36185 6137 36219 6171
rect 36277 6137 36311 6171
rect 36829 6137 36863 6171
rect 39221 6137 39255 6171
rect 40877 6137 40911 6171
rect 41153 6137 41187 6171
rect 43085 6137 43119 6171
rect 43361 6137 43395 6171
rect 44281 6137 44315 6171
rect 21373 6069 21407 6103
rect 23121 6069 23155 6103
rect 24685 6069 24719 6103
rect 25145 6069 25179 6103
rect 29469 6069 29503 6103
rect 30113 6069 30147 6103
rect 31493 6069 31527 6103
rect 34253 6069 34287 6103
rect 35633 6069 35667 6103
rect 36001 6069 36035 6103
rect 40233 6069 40267 6103
rect 45569 6069 45603 6103
rect 46397 6069 46431 6103
rect 23305 5865 23339 5899
rect 27997 5865 28031 5899
rect 30573 5865 30607 5899
rect 31401 5865 31435 5899
rect 32229 5865 32263 5899
rect 34805 5865 34839 5899
rect 35633 5865 35667 5899
rect 39129 5865 39163 5899
rect 39681 5865 39715 5899
rect 40509 5865 40543 5899
rect 40877 5865 40911 5899
rect 41981 5865 42015 5899
rect 44741 5865 44775 5899
rect 46121 5865 46155 5899
rect 22747 5797 22781 5831
rect 24317 5797 24351 5831
rect 24869 5797 24903 5831
rect 27169 5797 27203 5831
rect 28911 5797 28945 5831
rect 37933 5797 37967 5831
rect 41423 5797 41457 5831
rect 43545 5797 43579 5831
rect 44925 5797 44959 5831
rect 21440 5729 21474 5763
rect 30481 5729 30515 5763
rect 30849 5729 30883 5763
rect 32413 5729 32447 5763
rect 32689 5729 32723 5763
rect 34437 5729 34471 5763
rect 35357 5729 35391 5763
rect 36220 5729 36254 5763
rect 45017 5729 45051 5763
rect 22385 5661 22419 5695
rect 24225 5661 24259 5695
rect 27077 5661 27111 5695
rect 27353 5661 27387 5695
rect 28549 5661 28583 5695
rect 37841 5661 37875 5695
rect 38485 5661 38519 5695
rect 39313 5661 39347 5695
rect 41061 5661 41095 5695
rect 43453 5661 43487 5695
rect 44097 5661 44131 5695
rect 21511 5593 21545 5627
rect 38853 5593 38887 5627
rect 22109 5525 22143 5559
rect 23765 5525 23799 5559
rect 25329 5525 25363 5559
rect 26893 5525 26927 5559
rect 29469 5525 29503 5559
rect 33333 5525 33367 5559
rect 36323 5525 36357 5559
rect 37013 5525 37047 5559
rect 40233 5525 40267 5559
rect 44373 5525 44407 5559
rect 20361 5321 20395 5355
rect 21557 5321 21591 5355
rect 21925 5321 21959 5355
rect 23489 5321 23523 5355
rect 24685 5321 24719 5355
rect 26341 5321 26375 5355
rect 27905 5321 27939 5355
rect 28549 5321 28583 5355
rect 30389 5321 30423 5355
rect 32321 5321 32355 5355
rect 34069 5321 34103 5355
rect 36369 5321 36403 5355
rect 36829 5321 36863 5355
rect 38025 5321 38059 5355
rect 38301 5321 38335 5355
rect 39589 5321 39623 5355
rect 42257 5321 42291 5355
rect 42579 5321 42613 5355
rect 43453 5321 43487 5355
rect 45017 5321 45051 5355
rect 40693 5253 40727 5287
rect 41521 5253 41555 5287
rect 41889 5253 41923 5287
rect 20545 5185 20579 5219
rect 21189 5185 21223 5219
rect 22569 5185 22603 5219
rect 23765 5185 23799 5219
rect 24409 5185 24443 5219
rect 25329 5185 25363 5219
rect 25605 5185 25639 5219
rect 26893 5185 26927 5219
rect 27169 5185 27203 5219
rect 31033 5185 31067 5219
rect 33609 5185 33643 5219
rect 35173 5185 35207 5219
rect 37013 5185 37047 5219
rect 39221 5185 39255 5219
rect 39865 5185 39899 5219
rect 40233 5185 40267 5219
rect 40969 5185 41003 5219
rect 43821 5185 43855 5219
rect 22017 5117 22051 5151
rect 22477 5117 22511 5151
rect 29101 5117 29135 5151
rect 29561 5117 29595 5151
rect 29837 5117 29871 5151
rect 33241 5117 33275 5151
rect 33517 5117 33551 5151
rect 38485 5117 38519 5151
rect 39037 5117 39071 5151
rect 42476 5117 42510 5151
rect 20637 5049 20671 5083
rect 23857 5049 23891 5083
rect 25145 5049 25179 5083
rect 25421 5049 25455 5083
rect 26709 5049 26743 5083
rect 26985 5049 27019 5083
rect 28273 5049 28307 5083
rect 30941 5049 30975 5083
rect 31354 5049 31388 5083
rect 35494 5049 35528 5083
rect 37105 5049 37139 5083
rect 37657 5049 37691 5083
rect 41061 5049 41095 5083
rect 43085 5049 43119 5083
rect 43913 5049 43947 5083
rect 44465 5049 44499 5083
rect 23121 4981 23155 5015
rect 29377 4981 29411 5015
rect 31953 4981 31987 5015
rect 32965 4981 32999 5015
rect 34437 4981 34471 5015
rect 36093 4981 36127 5015
rect 20545 4777 20579 4811
rect 22385 4777 22419 4811
rect 22707 4777 22741 4811
rect 24961 4777 24995 4811
rect 25559 4777 25593 4811
rect 26985 4777 27019 4811
rect 28273 4777 28307 4811
rect 29653 4777 29687 4811
rect 30527 4777 30561 4811
rect 32275 4777 32309 4811
rect 32689 4777 32723 4811
rect 33057 4777 33091 4811
rect 35541 4777 35575 4811
rect 39037 4777 39071 4811
rect 43085 4777 43119 4811
rect 45339 4777 45373 4811
rect 23765 4709 23799 4743
rect 24317 4709 24351 4743
rect 24593 4709 24627 4743
rect 28733 4709 28767 4743
rect 33930 4709 33964 4743
rect 35173 4709 35207 4743
rect 36277 4709 36311 4743
rect 39681 4709 39715 4743
rect 39773 4709 39807 4743
rect 43821 4709 43855 4743
rect 44373 4709 44407 4743
rect 22636 4641 22670 4675
rect 25421 4641 25455 4675
rect 26617 4641 26651 4675
rect 30456 4641 30490 4675
rect 31217 4641 31251 4675
rect 32172 4641 32206 4675
rect 38301 4641 38335 4675
rect 38485 4641 38519 4675
rect 41220 4641 41254 4675
rect 42232 4641 42266 4675
rect 45268 4641 45302 4675
rect 23673 4573 23707 4607
rect 28641 4573 28675 4607
rect 29285 4573 29319 4607
rect 30941 4573 30975 4607
rect 33609 4573 33643 4607
rect 36185 4573 36219 4607
rect 36829 4573 36863 4607
rect 38577 4573 38611 4607
rect 39957 4573 39991 4607
rect 43729 4573 43763 4607
rect 42303 4505 42337 4539
rect 22109 4437 22143 4471
rect 34529 4437 34563 4471
rect 37473 4437 37507 4471
rect 40785 4437 40819 4471
rect 41291 4437 41325 4471
rect 41889 4437 41923 4471
rect 22937 4233 22971 4267
rect 25421 4233 25455 4267
rect 26985 4233 27019 4267
rect 28319 4233 28353 4267
rect 29009 4233 29043 4267
rect 30941 4233 30975 4267
rect 32137 4233 32171 4267
rect 34069 4233 34103 4267
rect 35311 4233 35345 4267
rect 38117 4233 38151 4267
rect 38485 4233 38519 4267
rect 40049 4233 40083 4267
rect 41613 4233 41647 4267
rect 43269 4233 43303 4267
rect 44373 4233 44407 4267
rect 21741 4165 21775 4199
rect 23949 4165 23983 4199
rect 25881 4165 25915 4199
rect 33701 4165 33735 4199
rect 35725 4165 35759 4199
rect 36001 4165 36035 4199
rect 37749 4165 37783 4199
rect 39681 4165 39715 4199
rect 44005 4165 44039 4199
rect 45385 4165 45419 4199
rect 28641 4097 28675 4131
rect 29653 4097 29687 4131
rect 31493 4097 31527 4131
rect 33057 4097 33091 4131
rect 43453 4097 43487 4131
rect 44741 4097 44775 4131
rect 21925 4029 21959 4063
rect 22385 4029 22419 4063
rect 24317 4029 24351 4063
rect 24409 4029 24443 4063
rect 24869 4029 24903 4063
rect 28248 4029 28282 4063
rect 34713 4029 34747 4063
rect 35240 4029 35274 4063
rect 36921 4029 36955 4063
rect 38669 4029 38703 4063
rect 39129 4029 39163 4063
rect 40785 4029 40819 4063
rect 44976 4029 45010 4063
rect 45753 4029 45787 4063
rect 22661 3961 22695 3995
rect 25145 3961 25179 3995
rect 26065 3961 26099 3995
rect 26157 3961 26191 3995
rect 26709 3961 26743 3995
rect 29377 3961 29411 3995
rect 29469 3961 29503 3995
rect 30665 3961 30699 3995
rect 31217 3961 31251 3995
rect 31309 3961 31343 3995
rect 32781 3961 32815 3995
rect 32873 3961 32907 3995
rect 36277 3961 36311 3995
rect 36369 3961 36403 3995
rect 39405 3961 39439 3995
rect 41889 3961 41923 3995
rect 41981 3961 42015 3995
rect 42533 3961 42567 3995
rect 43545 3961 43579 3995
rect 45063 3961 45097 3995
rect 23397 3893 23431 3927
rect 28089 3893 28123 3927
rect 32597 3893 32631 3927
rect 40923 3893 40957 3927
rect 41245 3893 41279 3927
rect 42809 3893 42843 3927
rect 23121 3689 23155 3723
rect 32275 3689 32309 3723
rect 32781 3689 32815 3723
rect 36461 3689 36495 3723
rect 36783 3689 36817 3723
rect 38117 3689 38151 3723
rect 39405 3689 39439 3723
rect 40785 3689 40819 3723
rect 44373 3689 44407 3723
rect 22563 3621 22597 3655
rect 26709 3621 26743 3655
rect 28543 3621 28577 3655
rect 33241 3621 33275 3655
rect 35218 3621 35252 3655
rect 37105 3621 37139 3655
rect 40186 3621 40220 3655
rect 41613 3621 41647 3655
rect 41797 3621 41831 3655
rect 41889 3621 41923 3655
rect 43545 3621 43579 3655
rect 21256 3553 21290 3587
rect 24685 3553 24719 3587
rect 24869 3553 24903 3587
rect 29377 3553 29411 3587
rect 30389 3553 30423 3587
rect 30849 3553 30883 3587
rect 32045 3553 32079 3587
rect 33425 3553 33459 3587
rect 33885 3553 33919 3587
rect 36680 3553 36714 3587
rect 38301 3553 38335 3587
rect 38761 3553 38795 3587
rect 39865 3553 39899 3587
rect 42441 3553 42475 3587
rect 22201 3485 22235 3519
rect 25145 3485 25179 3519
rect 25421 3485 25455 3519
rect 26617 3485 26651 3519
rect 26893 3485 26927 3519
rect 28181 3485 28215 3519
rect 30941 3485 30975 3519
rect 34069 3485 34103 3519
rect 34897 3485 34931 3519
rect 39037 3485 39071 3519
rect 43453 3485 43487 3519
rect 21327 3417 21361 3451
rect 44005 3417 44039 3451
rect 22017 3349 22051 3383
rect 24041 3349 24075 3383
rect 25973 3349 26007 3383
rect 27629 3349 27663 3383
rect 28089 3349 28123 3383
rect 29101 3349 29135 3383
rect 34713 3349 34747 3383
rect 35817 3349 35851 3383
rect 36185 3349 36219 3383
rect 20959 3145 20993 3179
rect 23121 3145 23155 3179
rect 24087 3145 24121 3179
rect 24501 3145 24535 3179
rect 26525 3145 26559 3179
rect 26893 3145 26927 3179
rect 29101 3145 29135 3179
rect 29929 3145 29963 3179
rect 31677 3145 31711 3179
rect 32137 3145 32171 3179
rect 34253 3145 34287 3179
rect 34621 3145 34655 3179
rect 35817 3145 35851 3179
rect 36553 3145 36587 3179
rect 39589 3145 39623 3179
rect 41797 3145 41831 3179
rect 42073 3145 42107 3179
rect 43361 3145 43395 3179
rect 43637 3145 43671 3179
rect 20729 3077 20763 3111
rect 22753 3077 22787 3111
rect 28365 3077 28399 3111
rect 29423 3077 29457 3111
rect 36093 3077 36127 3111
rect 39957 3077 39991 3111
rect 40233 3077 40267 3111
rect 44833 3077 44867 3111
rect 21373 3009 21407 3043
rect 24961 3009 24995 3043
rect 30757 3009 30791 3043
rect 32781 3009 32815 3043
rect 38117 3009 38151 3043
rect 38669 3009 38703 3043
rect 40509 3009 40543 3043
rect 42349 3009 42383 3043
rect 42625 3009 42659 3043
rect 43913 3009 43947 3043
rect 44189 3009 44223 3043
rect 20888 2941 20922 2975
rect 21833 2941 21867 2975
rect 24016 2941 24050 2975
rect 27445 2941 27479 2975
rect 29320 2941 29354 2975
rect 33149 2941 33183 2975
rect 33425 2941 33459 2975
rect 33701 2941 33735 2975
rect 34897 2941 34931 2975
rect 37013 2941 37047 2975
rect 37105 2941 37139 2975
rect 37565 2941 37599 2975
rect 41429 2941 41463 2975
rect 21741 2873 21775 2907
rect 22195 2873 22229 2907
rect 24869 2873 24903 2907
rect 25323 2873 25357 2907
rect 27353 2873 27387 2907
rect 27807 2873 27841 2907
rect 30665 2873 30699 2907
rect 31078 2873 31112 2907
rect 33977 2873 34011 2907
rect 37841 2873 37875 2907
rect 39031 2873 39065 2907
rect 40830 2873 40864 2907
rect 42441 2873 42475 2907
rect 44005 2873 44039 2907
rect 23397 2805 23431 2839
rect 25881 2805 25915 2839
rect 28641 2805 28675 2839
rect 30297 2805 30331 2839
rect 35265 2805 35299 2839
rect 38485 2805 38519 2839
rect 21649 2601 21683 2635
rect 22845 2601 22879 2635
rect 24501 2601 24535 2635
rect 25881 2601 25915 2635
rect 27031 2601 27065 2635
rect 28181 2601 28215 2635
rect 29837 2601 29871 2635
rect 30849 2601 30883 2635
rect 31447 2601 31481 2635
rect 32735 2601 32769 2635
rect 37335 2601 37369 2635
rect 38025 2601 38059 2635
rect 38669 2601 38703 2635
rect 40049 2601 40083 2635
rect 40509 2601 40543 2635
rect 40969 2601 41003 2635
rect 41613 2601 41647 2635
rect 22569 2533 22603 2567
rect 24777 2533 24811 2567
rect 25282 2533 25316 2567
rect 27629 2533 27663 2567
rect 29193 2533 29227 2567
rect 34345 2533 34379 2567
rect 35173 2533 35207 2567
rect 35770 2533 35804 2567
rect 37657 2533 37691 2567
rect 39174 2533 39208 2567
rect 41797 2533 41831 2567
rect 41889 2533 41923 2567
rect 42441 2533 42475 2567
rect 43361 2533 43395 2567
rect 21833 2465 21867 2499
rect 22293 2465 22327 2499
rect 24961 2465 24995 2499
rect 26617 2465 26651 2499
rect 26928 2465 26962 2499
rect 27997 2465 28031 2499
rect 28365 2465 28399 2499
rect 28641 2465 28675 2499
rect 29561 2465 29595 2499
rect 30021 2465 30055 2499
rect 30205 2465 30239 2499
rect 31217 2465 31251 2499
rect 31376 2465 31410 2499
rect 32045 2465 32079 2499
rect 32632 2465 32666 2499
rect 33333 2465 33367 2499
rect 33885 2465 33919 2499
rect 34161 2465 34195 2499
rect 35449 2465 35483 2499
rect 36645 2465 36679 2499
rect 37232 2465 37266 2499
rect 38853 2465 38887 2499
rect 39773 2465 39807 2499
rect 44040 2465 44074 2499
rect 44465 2465 44499 2499
rect 21005 2397 21039 2431
rect 26157 2397 26191 2431
rect 34621 2397 34655 2431
rect 36369 2329 36403 2363
rect 44143 2329 44177 2363
rect 32413 2261 32447 2295
rect 42717 2261 42751 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 48852 47354
rect 1104 47280 48852 47302
rect 41046 47104 41052 47116
rect 41007 47076 41052 47104
rect 41046 47064 41052 47076
rect 41104 47064 41110 47116
rect 41279 46903 41337 46909
rect 41279 46869 41291 46903
rect 41325 46900 41337 46903
rect 41506 46900 41512 46912
rect 41325 46872 41512 46900
rect 41325 46869 41337 46872
rect 41279 46863 41337 46869
rect 41506 46860 41512 46872
rect 41564 46860 41570 46912
rect 1104 46810 48852 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 48852 46810
rect 1104 46736 48852 46758
rect 36078 46588 36084 46640
rect 36136 46628 36142 46640
rect 41046 46628 41052 46640
rect 36136 46600 41052 46628
rect 36136 46588 36142 46600
rect 41046 46588 41052 46600
rect 41104 46628 41110 46640
rect 41141 46631 41199 46637
rect 41141 46628 41153 46631
rect 41104 46600 41153 46628
rect 41104 46588 41110 46600
rect 41141 46597 41153 46600
rect 41187 46597 41199 46631
rect 41141 46591 41199 46597
rect 40865 46563 40923 46569
rect 40865 46529 40877 46563
rect 40911 46560 40923 46563
rect 41506 46560 41512 46572
rect 40911 46532 41512 46560
rect 40911 46529 40923 46532
rect 40865 46523 40923 46529
rect 41506 46520 41512 46532
rect 41564 46520 41570 46572
rect 27960 46495 28018 46501
rect 27960 46461 27972 46495
rect 28006 46492 28018 46495
rect 36056 46495 36114 46501
rect 28006 46464 28488 46492
rect 28006 46461 28018 46464
rect 27960 46455 28018 46461
rect 28460 46368 28488 46464
rect 36056 46461 36068 46495
rect 36102 46492 36114 46495
rect 36262 46492 36268 46504
rect 36102 46464 36268 46492
rect 36102 46461 36114 46464
rect 36056 46455 36114 46461
rect 36262 46452 36268 46464
rect 36320 46492 36326 46504
rect 36449 46495 36507 46501
rect 36449 46492 36461 46495
rect 36320 46464 36461 46492
rect 36320 46452 36326 46464
rect 36449 46461 36461 46464
rect 36495 46461 36507 46495
rect 36449 46455 36507 46461
rect 41601 46427 41659 46433
rect 41601 46393 41613 46427
rect 41647 46424 41659 46427
rect 41690 46424 41696 46436
rect 41647 46396 41696 46424
rect 41647 46393 41659 46396
rect 41601 46387 41659 46393
rect 41690 46384 41696 46396
rect 41748 46384 41754 46436
rect 42153 46427 42211 46433
rect 42153 46393 42165 46427
rect 42199 46424 42211 46427
rect 42334 46424 42340 46436
rect 42199 46396 42340 46424
rect 42199 46393 42211 46396
rect 42153 46387 42211 46393
rect 42334 46384 42340 46396
rect 42392 46384 42398 46436
rect 28031 46359 28089 46365
rect 28031 46325 28043 46359
rect 28077 46356 28089 46359
rect 28166 46356 28172 46368
rect 28077 46328 28172 46356
rect 28077 46325 28089 46328
rect 28031 46319 28089 46325
rect 28166 46316 28172 46328
rect 28224 46316 28230 46368
rect 28442 46356 28448 46368
rect 28403 46328 28448 46356
rect 28442 46316 28448 46328
rect 28500 46316 28506 46368
rect 34698 46316 34704 46368
rect 34756 46356 34762 46368
rect 34885 46359 34943 46365
rect 34885 46356 34897 46359
rect 34756 46328 34897 46356
rect 34756 46316 34762 46328
rect 34885 46325 34897 46328
rect 34931 46325 34943 46359
rect 34885 46319 34943 46325
rect 36127 46359 36185 46365
rect 36127 46325 36139 46359
rect 36173 46356 36185 46359
rect 36354 46356 36360 46368
rect 36173 46328 36360 46356
rect 36173 46325 36185 46328
rect 36127 46319 36185 46325
rect 36354 46316 36360 46328
rect 36412 46316 36418 46368
rect 1104 46266 48852 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 48852 46266
rect 1104 46192 48852 46214
rect 30190 46152 30196 46164
rect 30151 46124 30196 46152
rect 30190 46112 30196 46124
rect 30248 46112 30254 46164
rect 36354 46112 36360 46164
rect 36412 46152 36418 46164
rect 36909 46155 36967 46161
rect 36909 46152 36921 46155
rect 36412 46124 36921 46152
rect 36412 46112 36418 46124
rect 36909 46121 36921 46124
rect 36955 46121 36967 46155
rect 43714 46152 43720 46164
rect 36909 46115 36967 46121
rect 39868 46124 43720 46152
rect 28445 46087 28503 46093
rect 28445 46053 28457 46087
rect 28491 46084 28503 46087
rect 28718 46084 28724 46096
rect 28491 46056 28724 46084
rect 28491 46053 28503 46056
rect 28445 46047 28503 46053
rect 28718 46044 28724 46056
rect 28776 46044 28782 46096
rect 34146 46044 34152 46096
rect 34204 46084 34210 46096
rect 34241 46087 34299 46093
rect 34241 46084 34253 46087
rect 34204 46056 34253 46084
rect 34204 46044 34210 46056
rect 34241 46053 34253 46056
rect 34287 46053 34299 46087
rect 34241 46047 34299 46053
rect 39868 46028 39896 46124
rect 43714 46112 43720 46124
rect 43772 46112 43778 46164
rect 41598 46044 41604 46096
rect 41656 46084 41662 46096
rect 41877 46087 41935 46093
rect 41877 46084 41889 46087
rect 41656 46056 41889 46084
rect 41656 46044 41662 46056
rect 41877 46053 41889 46056
rect 41923 46053 41935 46087
rect 41877 46047 41935 46053
rect 30374 46016 30380 46028
rect 30335 45988 30380 46016
rect 30374 45976 30380 45988
rect 30432 45976 30438 46028
rect 30653 46019 30711 46025
rect 30653 45985 30665 46019
rect 30699 46016 30711 46019
rect 31202 46016 31208 46028
rect 30699 45988 31208 46016
rect 30699 45985 30711 45988
rect 30653 45979 30711 45985
rect 31202 45976 31208 45988
rect 31260 45976 31266 46028
rect 34793 46019 34851 46025
rect 34793 45985 34805 46019
rect 34839 46016 34851 46019
rect 35618 46016 35624 46028
rect 34839 45988 35624 46016
rect 34839 45985 34851 45988
rect 34793 45979 34851 45985
rect 35618 45976 35624 45988
rect 35676 46016 35682 46028
rect 36538 46016 36544 46028
rect 35676 45988 36544 46016
rect 35676 45976 35682 45988
rect 36538 45976 36544 45988
rect 36596 45976 36602 46028
rect 39850 46016 39856 46028
rect 39811 45988 39856 46016
rect 39850 45976 39856 45988
rect 39908 45976 39914 46028
rect 27249 45951 27307 45957
rect 27249 45917 27261 45951
rect 27295 45948 27307 45951
rect 28353 45951 28411 45957
rect 28353 45948 28365 45951
rect 27295 45920 28365 45948
rect 27295 45917 27307 45920
rect 27249 45911 27307 45917
rect 28353 45917 28365 45920
rect 28399 45948 28411 45951
rect 28626 45948 28632 45960
rect 28399 45920 28632 45948
rect 28399 45917 28411 45920
rect 28353 45911 28411 45917
rect 28626 45908 28632 45920
rect 28684 45908 28690 45960
rect 28994 45948 29000 45960
rect 28955 45920 29000 45948
rect 28994 45908 29000 45920
rect 29052 45908 29058 45960
rect 34149 45951 34207 45957
rect 34149 45948 34161 45951
rect 33888 45920 34161 45948
rect 25314 45812 25320 45824
rect 25275 45784 25320 45812
rect 25314 45772 25320 45784
rect 25372 45772 25378 45824
rect 32858 45812 32864 45824
rect 32819 45784 32864 45812
rect 32858 45772 32864 45784
rect 32916 45772 32922 45824
rect 33318 45772 33324 45824
rect 33376 45812 33382 45824
rect 33888 45821 33916 45920
rect 34149 45917 34161 45920
rect 34195 45917 34207 45951
rect 34149 45911 34207 45917
rect 35989 45951 36047 45957
rect 35989 45917 36001 45951
rect 36035 45948 36047 45951
rect 36078 45948 36084 45960
rect 36035 45920 36084 45948
rect 36035 45917 36047 45920
rect 35989 45911 36047 45917
rect 36078 45908 36084 45920
rect 36136 45908 36142 45960
rect 41782 45948 41788 45960
rect 41743 45920 41788 45948
rect 41782 45908 41788 45920
rect 41840 45908 41846 45960
rect 36219 45883 36277 45889
rect 36219 45849 36231 45883
rect 36265 45880 36277 45883
rect 38013 45883 38071 45889
rect 38013 45880 38025 45883
rect 36265 45852 38025 45880
rect 36265 45849 36277 45852
rect 36219 45843 36277 45849
rect 38013 45849 38025 45852
rect 38059 45880 38071 45883
rect 38102 45880 38108 45892
rect 38059 45852 38108 45880
rect 38059 45849 38071 45852
rect 38013 45843 38071 45849
rect 38102 45840 38108 45852
rect 38160 45840 38166 45892
rect 42334 45880 42340 45892
rect 42295 45852 42340 45880
rect 42334 45840 42340 45852
rect 42392 45840 42398 45892
rect 33873 45815 33931 45821
rect 33873 45812 33885 45815
rect 33376 45784 33885 45812
rect 33376 45772 33382 45784
rect 33873 45781 33885 45784
rect 33919 45781 33931 45815
rect 33873 45775 33931 45781
rect 36446 45772 36452 45824
rect 36504 45812 36510 45824
rect 36541 45815 36599 45821
rect 36541 45812 36553 45815
rect 36504 45784 36553 45812
rect 36504 45772 36510 45784
rect 36541 45781 36553 45784
rect 36587 45781 36599 45815
rect 36541 45775 36599 45781
rect 39991 45815 40049 45821
rect 39991 45781 40003 45815
rect 40037 45812 40049 45815
rect 40586 45812 40592 45824
rect 40037 45784 40592 45812
rect 40037 45781 40049 45784
rect 39991 45775 40049 45781
rect 40586 45772 40592 45784
rect 40644 45772 40650 45824
rect 40678 45772 40684 45824
rect 40736 45812 40742 45824
rect 41417 45815 41475 45821
rect 41417 45812 41429 45815
rect 40736 45784 41429 45812
rect 40736 45772 40742 45784
rect 41417 45781 41429 45784
rect 41463 45812 41475 45815
rect 41690 45812 41696 45824
rect 41463 45784 41696 45812
rect 41463 45781 41475 45784
rect 41417 45775 41475 45781
rect 41690 45772 41696 45784
rect 41748 45812 41754 45824
rect 42150 45812 42156 45824
rect 41748 45784 42156 45812
rect 41748 45772 41754 45784
rect 42150 45772 42156 45784
rect 42208 45772 42214 45824
rect 1104 45722 48852 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 48852 45722
rect 1104 45648 48852 45670
rect 18874 45568 18880 45620
rect 18932 45608 18938 45620
rect 21542 45608 21548 45620
rect 18932 45580 21548 45608
rect 18932 45568 18938 45580
rect 21542 45568 21548 45580
rect 21600 45568 21606 45620
rect 28626 45608 28632 45620
rect 28587 45580 28632 45608
rect 28626 45568 28632 45580
rect 28684 45568 28690 45620
rect 28718 45568 28724 45620
rect 28776 45608 28782 45620
rect 30193 45611 30251 45617
rect 30193 45608 30205 45611
rect 28776 45580 30205 45608
rect 28776 45568 28782 45580
rect 25961 45475 26019 45481
rect 25961 45441 25973 45475
rect 26007 45472 26019 45475
rect 27985 45475 28043 45481
rect 27985 45472 27997 45475
rect 26007 45444 27997 45472
rect 26007 45441 26019 45444
rect 25961 45435 26019 45441
rect 27985 45441 27997 45444
rect 28031 45472 28043 45475
rect 28718 45472 28724 45484
rect 28031 45444 28724 45472
rect 28031 45441 28043 45444
rect 27985 45435 28043 45441
rect 28718 45432 28724 45444
rect 28776 45432 28782 45484
rect 25314 45336 25320 45348
rect 25275 45308 25320 45336
rect 25314 45296 25320 45308
rect 25372 45296 25378 45348
rect 25406 45296 25412 45348
rect 25464 45336 25470 45348
rect 27157 45339 27215 45345
rect 25464 45308 25509 45336
rect 25464 45296 25470 45308
rect 27157 45305 27169 45339
rect 27203 45336 27215 45339
rect 27706 45336 27712 45348
rect 27203 45308 27712 45336
rect 27203 45305 27215 45308
rect 27157 45299 27215 45305
rect 27706 45296 27712 45308
rect 27764 45296 27770 45348
rect 27801 45339 27859 45345
rect 27801 45305 27813 45339
rect 27847 45336 27859 45339
rect 28828 45336 28856 45580
rect 30193 45577 30205 45580
rect 30239 45577 30251 45611
rect 30193 45571 30251 45577
rect 30374 45568 30380 45620
rect 30432 45608 30438 45620
rect 30469 45611 30527 45617
rect 30469 45608 30481 45611
rect 30432 45580 30481 45608
rect 30432 45568 30438 45580
rect 30469 45577 30481 45580
rect 30515 45577 30527 45611
rect 34698 45608 34704 45620
rect 34659 45580 34704 45608
rect 30469 45571 30527 45577
rect 34698 45568 34704 45580
rect 34756 45608 34762 45620
rect 34756 45580 35020 45608
rect 34756 45568 34762 45580
rect 29273 45475 29331 45481
rect 29273 45441 29285 45475
rect 29319 45472 29331 45475
rect 29362 45472 29368 45484
rect 29319 45444 29368 45472
rect 29319 45441 29331 45444
rect 29273 45435 29331 45441
rect 29362 45432 29368 45444
rect 29420 45472 29426 45484
rect 30190 45472 30196 45484
rect 29420 45444 30196 45472
rect 29420 45432 29426 45444
rect 30190 45432 30196 45444
rect 30248 45432 30254 45484
rect 34992 45481 35020 45580
rect 36262 45568 36268 45620
rect 36320 45608 36326 45620
rect 39850 45608 39856 45620
rect 36320 45580 39856 45608
rect 36320 45568 36326 45580
rect 39850 45568 39856 45580
rect 39908 45568 39914 45620
rect 42150 45608 42156 45620
rect 42111 45580 42156 45608
rect 42150 45568 42156 45580
rect 42208 45608 42214 45620
rect 42518 45608 42524 45620
rect 42208 45580 42524 45608
rect 42208 45568 42214 45580
rect 42518 45568 42524 45580
rect 42576 45568 42582 45620
rect 35529 45543 35587 45549
rect 35529 45509 35541 45543
rect 35575 45540 35587 45543
rect 35575 45512 36676 45540
rect 35575 45509 35587 45512
rect 35529 45503 35587 45509
rect 34977 45475 35035 45481
rect 34977 45441 34989 45475
rect 35023 45441 35035 45475
rect 34977 45435 35035 45441
rect 36354 45432 36360 45484
rect 36412 45472 36418 45484
rect 36541 45475 36599 45481
rect 36541 45472 36553 45475
rect 36412 45444 36553 45472
rect 36412 45432 36418 45444
rect 36541 45441 36553 45444
rect 36587 45441 36599 45475
rect 36648 45472 36676 45512
rect 41782 45500 41788 45552
rect 41840 45540 41846 45552
rect 43349 45543 43407 45549
rect 43349 45540 43361 45543
rect 41840 45512 43361 45540
rect 41840 45500 41846 45512
rect 43349 45509 43361 45512
rect 43395 45509 43407 45543
rect 43349 45503 43407 45509
rect 36814 45472 36820 45484
rect 36648 45444 36820 45472
rect 36541 45435 36599 45441
rect 36814 45432 36820 45444
rect 36872 45432 36878 45484
rect 38102 45472 38108 45484
rect 38063 45444 38108 45472
rect 38102 45432 38108 45444
rect 38160 45432 38166 45484
rect 38378 45472 38384 45484
rect 38339 45444 38384 45472
rect 38378 45432 38384 45444
rect 38436 45432 38442 45484
rect 40586 45472 40592 45484
rect 40547 45444 40592 45472
rect 40586 45432 40592 45444
rect 40644 45432 40650 45484
rect 42426 45472 42432 45484
rect 42339 45444 42432 45472
rect 42426 45432 42432 45444
rect 42484 45472 42490 45484
rect 44039 45475 44097 45481
rect 44039 45472 44051 45475
rect 42484 45444 44051 45472
rect 42484 45432 42490 45444
rect 44039 45441 44051 45444
rect 44085 45441 44097 45475
rect 44039 45435 44097 45441
rect 32769 45407 32827 45413
rect 32769 45373 32781 45407
rect 32815 45404 32827 45407
rect 32858 45404 32864 45416
rect 32815 45376 32864 45404
rect 32815 45373 32827 45376
rect 32769 45367 32827 45373
rect 32858 45364 32864 45376
rect 32916 45364 32922 45416
rect 43952 45407 44010 45413
rect 43952 45373 43964 45407
rect 43998 45404 44010 45407
rect 43998 45376 44496 45404
rect 43998 45373 44010 45376
rect 43952 45367 44010 45373
rect 27847 45308 28856 45336
rect 29089 45339 29147 45345
rect 27847 45305 27859 45308
rect 27801 45299 27859 45305
rect 29089 45305 29101 45339
rect 29135 45336 29147 45339
rect 29635 45339 29693 45345
rect 29635 45336 29647 45339
rect 29135 45308 29647 45336
rect 29135 45305 29147 45308
rect 29089 45299 29147 45305
rect 29635 45305 29647 45308
rect 29681 45336 29693 45339
rect 30190 45336 30196 45348
rect 29681 45308 30196 45336
rect 29681 45305 29693 45308
rect 29635 45299 29693 45305
rect 25130 45268 25136 45280
rect 25091 45240 25136 45268
rect 25130 45228 25136 45240
rect 25188 45228 25194 45280
rect 27525 45271 27583 45277
rect 27525 45237 27537 45271
rect 27571 45268 27583 45271
rect 27614 45268 27620 45280
rect 27571 45240 27620 45268
rect 27571 45237 27583 45240
rect 27525 45231 27583 45237
rect 27614 45228 27620 45240
rect 27672 45268 27678 45280
rect 27816 45268 27844 45299
rect 30190 45296 30196 45308
rect 30248 45296 30254 45348
rect 33091 45339 33149 45345
rect 33091 45305 33103 45339
rect 33137 45305 33149 45339
rect 34146 45336 34152 45348
rect 34059 45308 34152 45336
rect 33091 45299 33149 45305
rect 27672 45240 27844 45268
rect 30929 45271 30987 45277
rect 27672 45228 27678 45240
rect 30929 45237 30941 45271
rect 30975 45268 30987 45271
rect 31202 45268 31208 45280
rect 30975 45240 31208 45268
rect 30975 45237 30987 45240
rect 30929 45231 30987 45237
rect 31202 45228 31208 45240
rect 31260 45228 31266 45280
rect 31294 45228 31300 45280
rect 31352 45268 31358 45280
rect 32214 45268 32220 45280
rect 31352 45240 32220 45268
rect 31352 45228 31358 45240
rect 32214 45228 32220 45240
rect 32272 45228 32278 45280
rect 32677 45271 32735 45277
rect 32677 45237 32689 45271
rect 32723 45268 32735 45271
rect 33106 45268 33134 45299
rect 34146 45296 34152 45308
rect 34204 45336 34210 45348
rect 35069 45339 35127 45345
rect 35069 45336 35081 45339
rect 34204 45308 35081 45336
rect 34204 45296 34210 45308
rect 35069 45305 35081 45308
rect 35115 45336 35127 45339
rect 35250 45336 35256 45348
rect 35115 45308 35256 45336
rect 35115 45305 35127 45308
rect 35069 45299 35127 45305
rect 35250 45296 35256 45308
rect 35308 45296 35314 45348
rect 36633 45339 36691 45345
rect 36633 45305 36645 45339
rect 36679 45305 36691 45339
rect 36633 45299 36691 45305
rect 38197 45339 38255 45345
rect 38197 45305 38209 45339
rect 38243 45305 38255 45339
rect 40678 45336 40684 45348
rect 40591 45308 40684 45336
rect 38197 45299 38255 45305
rect 33410 45268 33416 45280
rect 32723 45240 33416 45268
rect 32723 45237 32735 45240
rect 32677 45231 32735 45237
rect 33410 45228 33416 45240
rect 33468 45228 33474 45280
rect 33689 45271 33747 45277
rect 33689 45237 33701 45271
rect 33735 45268 33747 45271
rect 34164 45268 34192 45296
rect 36078 45268 36084 45280
rect 33735 45240 34192 45268
rect 36039 45240 36084 45268
rect 33735 45237 33747 45240
rect 33689 45231 33747 45237
rect 36078 45228 36084 45240
rect 36136 45228 36142 45280
rect 36446 45228 36452 45280
rect 36504 45268 36510 45280
rect 36648 45268 36676 45299
rect 37829 45271 37887 45277
rect 37829 45268 37841 45271
rect 36504 45240 37841 45268
rect 36504 45228 36510 45240
rect 37829 45237 37841 45240
rect 37875 45268 37887 45271
rect 38212 45268 38240 45299
rect 40678 45296 40684 45308
rect 40736 45296 40742 45348
rect 41233 45339 41291 45345
rect 41233 45305 41245 45339
rect 41279 45336 41291 45339
rect 41506 45336 41512 45348
rect 41279 45308 41512 45336
rect 41279 45305 41291 45308
rect 41233 45299 41291 45305
rect 41506 45296 41512 45308
rect 41564 45296 41570 45348
rect 42518 45336 42524 45348
rect 41708 45308 42288 45336
rect 42479 45308 42524 45336
rect 37875 45240 38240 45268
rect 37875 45237 37887 45240
rect 37829 45231 37887 45237
rect 39574 45228 39580 45280
rect 39632 45268 39638 45280
rect 40221 45271 40279 45277
rect 40221 45268 40233 45271
rect 39632 45240 40233 45268
rect 39632 45228 39638 45240
rect 40221 45237 40233 45240
rect 40267 45268 40279 45271
rect 40696 45268 40724 45296
rect 40267 45240 40724 45268
rect 40267 45237 40279 45240
rect 40221 45231 40279 45237
rect 41598 45228 41604 45280
rect 41656 45268 41662 45280
rect 41708 45277 41736 45308
rect 41693 45271 41751 45277
rect 41693 45268 41705 45271
rect 41656 45240 41705 45268
rect 41656 45228 41662 45240
rect 41693 45237 41705 45240
rect 41739 45237 41751 45271
rect 42260 45268 42288 45308
rect 42518 45296 42524 45308
rect 42576 45296 42582 45348
rect 43073 45339 43131 45345
rect 43073 45305 43085 45339
rect 43119 45336 43131 45339
rect 43714 45336 43720 45348
rect 43119 45308 43720 45336
rect 43119 45305 43131 45308
rect 43073 45299 43131 45305
rect 43714 45296 43720 45308
rect 43772 45296 43778 45348
rect 43806 45268 43812 45280
rect 42260 45240 43812 45268
rect 41693 45231 41751 45237
rect 43806 45228 43812 45240
rect 43864 45228 43870 45280
rect 44468 45277 44496 45376
rect 44453 45271 44511 45277
rect 44453 45237 44465 45271
rect 44499 45268 44511 45271
rect 44818 45268 44824 45280
rect 44499 45240 44824 45268
rect 44499 45237 44511 45240
rect 44453 45231 44511 45237
rect 44818 45228 44824 45240
rect 44876 45228 44882 45280
rect 1104 45178 48852 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 48852 45178
rect 1104 45104 48852 45126
rect 27614 45064 27620 45076
rect 27575 45036 27620 45064
rect 27614 45024 27620 45036
rect 27672 45024 27678 45076
rect 29362 45064 29368 45076
rect 29323 45036 29368 45064
rect 29362 45024 29368 45036
rect 29420 45024 29426 45076
rect 30374 45024 30380 45076
rect 30432 45064 30438 45076
rect 30432 45036 32168 45064
rect 30432 45024 30438 45036
rect 25041 44999 25099 45005
rect 25041 44965 25053 44999
rect 25087 44996 25099 44999
rect 25130 44996 25136 45008
rect 25087 44968 25136 44996
rect 25087 44965 25099 44968
rect 25041 44959 25099 44965
rect 25130 44956 25136 44968
rect 25188 44996 25194 45008
rect 25406 44996 25412 45008
rect 25188 44968 25412 44996
rect 25188 44956 25194 44968
rect 25406 44956 25412 44968
rect 25464 44956 25470 45008
rect 28166 44956 28172 45008
rect 28224 44996 28230 45008
rect 28353 44999 28411 45005
rect 28353 44996 28365 44999
rect 28224 44968 28365 44996
rect 28224 44956 28230 44968
rect 28353 44965 28365 44968
rect 28399 44965 28411 44999
rect 28353 44959 28411 44965
rect 28442 44956 28448 45008
rect 28500 44996 28506 45008
rect 28994 44996 29000 45008
rect 28500 44968 28545 44996
rect 28955 44968 29000 44996
rect 28500 44956 28506 44968
rect 28994 44956 29000 44968
rect 29052 44956 29058 45008
rect 32140 44940 32168 45036
rect 32214 45024 32220 45076
rect 32272 45064 32278 45076
rect 36078 45064 36084 45076
rect 32272 45036 36084 45064
rect 32272 45024 32278 45036
rect 36078 45024 36084 45036
rect 36136 45024 36142 45076
rect 38378 45064 38384 45076
rect 36188 45036 38384 45064
rect 32858 44996 32864 45008
rect 32819 44968 32864 44996
rect 32858 44956 32864 44968
rect 32916 44956 32922 45008
rect 34146 44996 34152 45008
rect 34107 44968 34152 44996
rect 34146 44956 34152 44968
rect 34204 44956 34210 45008
rect 34701 44999 34759 45005
rect 34701 44965 34713 44999
rect 34747 44996 34759 44999
rect 34790 44996 34796 45008
rect 34747 44968 34796 44996
rect 34747 44965 34759 44968
rect 34701 44959 34759 44965
rect 34790 44956 34796 44968
rect 34848 44996 34854 45008
rect 36188 44996 36216 45036
rect 38378 45024 38384 45036
rect 38436 45024 38442 45076
rect 40586 45064 40592 45076
rect 40547 45036 40592 45064
rect 40586 45024 40592 45036
rect 40644 45024 40650 45076
rect 42426 45064 42432 45076
rect 42387 45036 42432 45064
rect 42426 45024 42432 45036
rect 42484 45024 42490 45076
rect 34848 44968 36216 44996
rect 36265 44999 36323 45005
rect 34848 44956 34854 44968
rect 36265 44965 36277 44999
rect 36311 44996 36323 44999
rect 36446 44996 36452 45008
rect 36311 44968 36452 44996
rect 36311 44965 36323 44968
rect 36265 44959 36323 44965
rect 36446 44956 36452 44968
rect 36504 44956 36510 45008
rect 36538 44956 36544 45008
rect 36596 44996 36602 45008
rect 36817 44999 36875 45005
rect 36817 44996 36829 44999
rect 36596 44968 36829 44996
rect 36596 44956 36602 44968
rect 36817 44965 36829 44968
rect 36863 44965 36875 44999
rect 36817 44959 36875 44965
rect 39663 44999 39721 45005
rect 39663 44965 39675 44999
rect 39709 44996 39721 44999
rect 39942 44996 39948 45008
rect 39709 44968 39948 44996
rect 39709 44965 39721 44968
rect 39663 44959 39721 44965
rect 39942 44956 39948 44968
rect 40000 44956 40006 45008
rect 40218 44956 40224 45008
rect 40276 44996 40282 45008
rect 41233 44999 41291 45005
rect 41233 44996 41245 44999
rect 40276 44968 41245 44996
rect 40276 44956 40282 44968
rect 41233 44965 41245 44968
rect 41279 44996 41291 44999
rect 41598 44996 41604 45008
rect 41279 44968 41604 44996
rect 41279 44965 41291 44968
rect 41233 44959 41291 44965
rect 41598 44956 41604 44968
rect 41656 44956 41662 45008
rect 43533 44999 43591 45005
rect 43533 44965 43545 44999
rect 43579 44996 43591 44999
rect 43806 44996 43812 45008
rect 43579 44968 43812 44996
rect 43579 44965 43591 44968
rect 43533 44959 43591 44965
rect 43806 44956 43812 44968
rect 43864 44956 43870 45008
rect 23842 44928 23848 44940
rect 23803 44900 23848 44928
rect 23842 44888 23848 44900
rect 23900 44888 23906 44940
rect 26881 44931 26939 44937
rect 26881 44897 26893 44931
rect 26927 44928 26939 44931
rect 27062 44928 27068 44940
rect 26927 44900 27068 44928
rect 26927 44897 26939 44900
rect 26881 44891 26939 44897
rect 27062 44888 27068 44900
rect 27120 44888 27126 44940
rect 30374 44928 30380 44940
rect 30335 44900 30380 44928
rect 30374 44888 30380 44900
rect 30432 44888 30438 44940
rect 30837 44931 30895 44937
rect 30837 44897 30849 44931
rect 30883 44928 30895 44931
rect 31202 44928 31208 44940
rect 30883 44900 31208 44928
rect 30883 44897 30895 44900
rect 30837 44891 30895 44897
rect 31202 44888 31208 44900
rect 31260 44888 31266 44940
rect 32122 44928 32128 44940
rect 32035 44900 32128 44928
rect 32122 44888 32128 44900
rect 32180 44888 32186 44940
rect 32214 44888 32220 44940
rect 32272 44928 32278 44940
rect 32585 44931 32643 44937
rect 32585 44928 32597 44931
rect 32272 44900 32597 44928
rect 32272 44888 32278 44900
rect 32585 44897 32597 44900
rect 32631 44897 32643 44931
rect 32585 44891 32643 44897
rect 37645 44931 37703 44937
rect 37645 44897 37657 44931
rect 37691 44928 37703 44931
rect 37734 44928 37740 44940
rect 37691 44900 37740 44928
rect 37691 44897 37703 44900
rect 37645 44891 37703 44897
rect 37734 44888 37740 44900
rect 37792 44888 37798 44940
rect 24946 44860 24952 44872
rect 24907 44832 24952 44860
rect 24946 44820 24952 44832
rect 25004 44820 25010 44872
rect 25593 44863 25651 44869
rect 25593 44829 25605 44863
rect 25639 44860 25651 44863
rect 25866 44860 25872 44872
rect 25639 44832 25872 44860
rect 25639 44829 25651 44832
rect 25593 44823 25651 44829
rect 25866 44820 25872 44832
rect 25924 44860 25930 44872
rect 27798 44860 27804 44872
rect 25924 44832 27804 44860
rect 25924 44820 25930 44832
rect 27798 44820 27804 44832
rect 27856 44820 27862 44872
rect 30742 44820 30748 44872
rect 30800 44860 30806 44872
rect 30929 44863 30987 44869
rect 30929 44860 30941 44863
rect 30800 44832 30941 44860
rect 30800 44820 30806 44832
rect 30929 44829 30941 44832
rect 30975 44829 30987 44863
rect 34054 44860 34060 44872
rect 34015 44832 34060 44860
rect 30929 44823 30987 44829
rect 34054 44820 34060 44832
rect 34112 44820 34118 44872
rect 36170 44860 36176 44872
rect 36083 44832 36176 44860
rect 36170 44820 36176 44832
rect 36228 44860 36234 44872
rect 37875 44863 37933 44869
rect 37875 44860 37887 44863
rect 36228 44832 37887 44860
rect 36228 44820 36234 44832
rect 37875 44829 37887 44832
rect 37921 44829 37933 44863
rect 39298 44860 39304 44872
rect 39259 44832 39304 44860
rect 37875 44823 37933 44829
rect 39298 44820 39304 44832
rect 39356 44820 39362 44872
rect 41141 44863 41199 44869
rect 41141 44829 41153 44863
rect 41187 44829 41199 44863
rect 41506 44860 41512 44872
rect 41467 44832 41512 44860
rect 41141 44823 41199 44829
rect 23983 44795 24041 44801
rect 23983 44761 23995 44795
rect 24029 44792 24041 44795
rect 24964 44792 24992 44820
rect 24029 44764 24992 44792
rect 35069 44795 35127 44801
rect 24029 44761 24041 44764
rect 23983 44755 24041 44761
rect 35069 44761 35081 44795
rect 35115 44792 35127 44795
rect 35250 44792 35256 44804
rect 35115 44764 35256 44792
rect 35115 44761 35127 44764
rect 35069 44755 35127 44761
rect 35250 44752 35256 44764
rect 35308 44752 35314 44804
rect 41156 44792 41184 44823
rect 41506 44820 41512 44832
rect 41564 44820 41570 44872
rect 43438 44860 43444 44872
rect 43399 44832 43444 44860
rect 43438 44820 43444 44832
rect 43496 44820 43502 44872
rect 43714 44860 43720 44872
rect 43675 44832 43720 44860
rect 43714 44820 43720 44832
rect 43772 44820 43778 44872
rect 41322 44792 41328 44804
rect 41156 44764 41328 44792
rect 41322 44752 41328 44764
rect 41380 44752 41386 44804
rect 27111 44727 27169 44733
rect 27111 44693 27123 44727
rect 27157 44724 27169 44727
rect 27430 44724 27436 44736
rect 27157 44696 27436 44724
rect 27157 44693 27169 44696
rect 27111 44687 27169 44693
rect 27430 44684 27436 44696
rect 27488 44684 27494 44736
rect 31386 44724 31392 44736
rect 31347 44696 31392 44724
rect 31386 44684 31392 44696
rect 31444 44684 31450 44736
rect 35342 44724 35348 44736
rect 35303 44696 35348 44724
rect 35342 44684 35348 44696
rect 35400 44684 35406 44736
rect 38562 44684 38568 44736
rect 38620 44724 38626 44736
rect 38657 44727 38715 44733
rect 38657 44724 38669 44727
rect 38620 44696 38669 44724
rect 38620 44684 38626 44696
rect 38657 44693 38669 44696
rect 38703 44693 38715 44727
rect 40218 44724 40224 44736
rect 40179 44696 40224 44724
rect 38657 44687 38715 44693
rect 40218 44684 40224 44696
rect 40276 44684 40282 44736
rect 1104 44634 48852 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 48852 44634
rect 1104 44560 48852 44582
rect 22278 44520 22284 44532
rect 22239 44492 22284 44520
rect 22278 44480 22284 44492
rect 22336 44480 22342 44532
rect 24946 44480 24952 44532
rect 25004 44520 25010 44532
rect 26145 44523 26203 44529
rect 26145 44520 26157 44523
rect 25004 44492 26157 44520
rect 25004 44480 25010 44492
rect 26145 44489 26157 44492
rect 26191 44489 26203 44523
rect 26145 44483 26203 44489
rect 28166 44480 28172 44532
rect 28224 44520 28230 44532
rect 28721 44523 28779 44529
rect 28721 44520 28733 44523
rect 28224 44492 28733 44520
rect 28224 44480 28230 44492
rect 28721 44489 28733 44492
rect 28767 44489 28779 44523
rect 28721 44483 28779 44489
rect 30285 44523 30343 44529
rect 30285 44489 30297 44523
rect 30331 44520 30343 44523
rect 30374 44520 30380 44532
rect 30331 44492 30380 44520
rect 30331 44489 30343 44492
rect 30285 44483 30343 44489
rect 30374 44480 30380 44492
rect 30432 44480 30438 44532
rect 32214 44520 32220 44532
rect 32175 44492 32220 44520
rect 32214 44480 32220 44492
rect 32272 44480 32278 44532
rect 32631 44523 32689 44529
rect 32631 44489 32643 44523
rect 32677 44520 32689 44523
rect 33318 44520 33324 44532
rect 32677 44492 33324 44520
rect 32677 44489 32689 44492
rect 32631 44483 32689 44489
rect 33318 44480 33324 44492
rect 33376 44480 33382 44532
rect 33413 44523 33471 44529
rect 33413 44489 33425 44523
rect 33459 44520 33471 44523
rect 33643 44523 33701 44529
rect 33643 44520 33655 44523
rect 33459 44492 33655 44520
rect 33459 44489 33471 44492
rect 33413 44483 33471 44489
rect 33643 44489 33655 44492
rect 33689 44520 33701 44523
rect 34054 44520 34060 44532
rect 33689 44492 34060 44520
rect 33689 44489 33701 44492
rect 33643 44483 33701 44489
rect 34054 44480 34060 44492
rect 34112 44480 34118 44532
rect 39574 44520 39580 44532
rect 39535 44492 39580 44520
rect 39574 44480 39580 44492
rect 39632 44480 39638 44532
rect 40218 44520 40224 44532
rect 40179 44492 40224 44520
rect 40218 44480 40224 44492
rect 40276 44480 40282 44532
rect 40635 44523 40693 44529
rect 40635 44489 40647 44523
rect 40681 44520 40693 44523
rect 41782 44520 41788 44532
rect 40681 44492 41788 44520
rect 40681 44489 40693 44492
rect 40635 44483 40693 44489
rect 41782 44480 41788 44492
rect 41840 44480 41846 44532
rect 42150 44480 42156 44532
rect 42208 44520 42214 44532
rect 42245 44523 42303 44529
rect 42245 44520 42257 44523
rect 42208 44492 42257 44520
rect 42208 44480 42214 44492
rect 42245 44489 42257 44492
rect 42291 44520 42303 44523
rect 42337 44523 42395 44529
rect 42337 44520 42349 44523
rect 42291 44492 42349 44520
rect 42291 44489 42303 44492
rect 42245 44483 42303 44489
rect 42337 44489 42349 44492
rect 42383 44489 42395 44523
rect 42337 44483 42395 44489
rect 27706 44412 27712 44464
rect 27764 44452 27770 44464
rect 29411 44455 29469 44461
rect 29411 44452 29423 44455
rect 27764 44424 29423 44452
rect 27764 44412 27770 44424
rect 29411 44421 29423 44424
rect 29457 44421 29469 44455
rect 29411 44415 29469 44421
rect 29825 44455 29883 44461
rect 29825 44421 29837 44455
rect 29871 44452 29883 44455
rect 33965 44455 34023 44461
rect 33965 44452 33977 44455
rect 29871 44424 33977 44452
rect 29871 44421 29883 44424
rect 29825 44415 29883 44421
rect 33965 44421 33977 44424
rect 34011 44452 34023 44455
rect 38565 44455 38623 44461
rect 34011 44424 37228 44452
rect 34011 44421 34023 44424
rect 33965 44415 34023 44421
rect 21542 44344 21548 44396
rect 21600 44384 21606 44396
rect 25682 44384 25688 44396
rect 21600 44356 23474 44384
rect 25643 44356 25688 44384
rect 21600 44344 21606 44356
rect 18744 44319 18802 44325
rect 18744 44285 18756 44319
rect 18790 44316 18802 44319
rect 18831 44319 18889 44325
rect 18790 44285 18803 44316
rect 18744 44279 18803 44285
rect 18831 44285 18843 44319
rect 18877 44316 18889 44319
rect 19150 44316 19156 44328
rect 18877 44288 19156 44316
rect 18877 44285 18889 44288
rect 18831 44279 18889 44285
rect 18775 44248 18803 44279
rect 19150 44276 19156 44288
rect 19208 44276 19214 44328
rect 21796 44319 21854 44325
rect 21796 44285 21808 44319
rect 21842 44316 21854 44319
rect 22278 44316 22284 44328
rect 21842 44288 22284 44316
rect 21842 44285 21854 44288
rect 21796 44279 21854 44285
rect 22278 44276 22284 44288
rect 22336 44276 22342 44328
rect 23446 44316 23474 44356
rect 25682 44344 25688 44356
rect 25740 44344 25746 44396
rect 27430 44384 27436 44396
rect 27391 44356 27436 44384
rect 27430 44344 27436 44356
rect 27488 44344 27494 44396
rect 27798 44384 27804 44396
rect 27759 44356 27804 44384
rect 27798 44344 27804 44356
rect 27856 44344 27862 44396
rect 24188 44319 24246 44325
rect 24188 44316 24200 44319
rect 23446 44288 24200 44316
rect 24188 44285 24200 44288
rect 24234 44316 24246 44319
rect 24581 44319 24639 44325
rect 24581 44316 24593 44319
rect 24234 44288 24593 44316
rect 24234 44285 24246 44288
rect 24188 44279 24246 44285
rect 24581 44285 24593 44288
rect 24627 44285 24639 44319
rect 24581 44279 24639 44285
rect 29340 44319 29398 44325
rect 29340 44285 29352 44319
rect 29386 44316 29398 44319
rect 29840 44316 29868 44415
rect 30745 44387 30803 44393
rect 30745 44353 30757 44387
rect 30791 44384 30803 44387
rect 30834 44384 30840 44396
rect 30791 44356 30840 44384
rect 30791 44353 30803 44356
rect 30745 44347 30803 44353
rect 30834 44344 30840 44356
rect 30892 44384 30898 44396
rect 31386 44384 31392 44396
rect 30892 44356 31392 44384
rect 30892 44344 30898 44356
rect 31386 44344 31392 44356
rect 31444 44344 31450 44396
rect 29386 44288 29868 44316
rect 32560 44319 32618 44325
rect 29386 44285 29398 44288
rect 29340 44279 29398 44285
rect 32560 44285 32572 44319
rect 32606 44316 32618 44319
rect 32950 44316 32956 44328
rect 32606 44288 32956 44316
rect 32606 44285 32618 44288
rect 32560 44279 32618 44285
rect 32950 44276 32956 44288
rect 33008 44276 33014 44328
rect 33572 44319 33630 44325
rect 33572 44285 33584 44319
rect 33618 44316 33630 44319
rect 33980 44316 34008 44415
rect 34977 44387 35035 44393
rect 34977 44353 34989 44387
rect 35023 44384 35035 44387
rect 35342 44384 35348 44396
rect 35023 44356 35348 44384
rect 35023 44353 35035 44356
rect 34977 44347 35035 44353
rect 35342 44344 35348 44356
rect 35400 44344 35406 44396
rect 35621 44387 35679 44393
rect 35621 44353 35633 44387
rect 35667 44384 35679 44387
rect 35986 44384 35992 44396
rect 35667 44356 35992 44384
rect 35667 44353 35679 44356
rect 35621 44347 35679 44353
rect 35986 44344 35992 44356
rect 36044 44384 36050 44396
rect 36817 44387 36875 44393
rect 36817 44384 36829 44387
rect 36044 44356 36829 44384
rect 36044 44344 36050 44356
rect 36817 44353 36829 44356
rect 36863 44353 36875 44387
rect 36817 44347 36875 44353
rect 33618 44288 34008 44316
rect 33618 44285 33630 44288
rect 33572 44279 33630 44285
rect 18775 44220 19288 44248
rect 19260 44192 19288 44220
rect 21358 44208 21364 44260
rect 21416 44248 21422 44260
rect 23842 44248 23848 44260
rect 21416 44220 23848 44248
rect 21416 44208 21422 44220
rect 23842 44208 23848 44220
rect 23900 44208 23906 44260
rect 24397 44251 24455 44257
rect 24397 44217 24409 44251
rect 24443 44248 24455 44251
rect 25222 44248 25228 44260
rect 24443 44220 25228 44248
rect 24443 44217 24455 44220
rect 24397 44211 24455 44217
rect 25222 44208 25228 44220
rect 25280 44208 25286 44260
rect 25317 44251 25375 44257
rect 25317 44217 25329 44251
rect 25363 44248 25375 44251
rect 25406 44248 25412 44260
rect 25363 44220 25412 44248
rect 25363 44217 25375 44220
rect 25317 44211 25375 44217
rect 19242 44180 19248 44192
rect 19203 44152 19248 44180
rect 19242 44140 19248 44152
rect 19300 44140 19306 44192
rect 21867 44183 21925 44189
rect 21867 44149 21879 44183
rect 21913 44180 21925 44183
rect 22002 44180 22008 44192
rect 21913 44152 22008 44180
rect 21913 44149 21925 44152
rect 21867 44143 21925 44149
rect 22002 44140 22008 44152
rect 22060 44140 22066 44192
rect 25041 44183 25099 44189
rect 25041 44149 25053 44183
rect 25087 44180 25099 44183
rect 25332 44180 25360 44211
rect 25406 44208 25412 44220
rect 25464 44208 25470 44260
rect 26697 44251 26755 44257
rect 26697 44217 26709 44251
rect 26743 44248 26755 44251
rect 27525 44251 27583 44257
rect 27525 44248 27537 44251
rect 26743 44220 27537 44248
rect 26743 44217 26755 44220
rect 26697 44211 26755 44217
rect 27525 44217 27537 44220
rect 27571 44248 27583 44251
rect 27614 44248 27620 44260
rect 27571 44220 27620 44248
rect 27571 44217 27583 44220
rect 27525 44211 27583 44217
rect 27614 44208 27620 44220
rect 27672 44208 27678 44260
rect 30190 44208 30196 44260
rect 30248 44248 30254 44260
rect 30561 44251 30619 44257
rect 30561 44248 30573 44251
rect 30248 44220 30573 44248
rect 30248 44208 30254 44220
rect 30561 44217 30573 44220
rect 30607 44248 30619 44251
rect 31066 44251 31124 44257
rect 31066 44248 31078 44251
rect 30607 44220 31078 44248
rect 30607 44217 30619 44220
rect 30561 44211 30619 44217
rect 31066 44217 31078 44220
rect 31112 44217 31124 44251
rect 31066 44211 31124 44217
rect 34425 44251 34483 44257
rect 34425 44217 34437 44251
rect 34471 44248 34483 44251
rect 35069 44251 35127 44257
rect 35069 44248 35081 44251
rect 34471 44220 35081 44248
rect 34471 44217 34483 44220
rect 34425 44211 34483 44217
rect 35069 44217 35081 44220
rect 35115 44248 35127 44251
rect 35250 44248 35256 44260
rect 35115 44220 35256 44248
rect 35115 44217 35127 44220
rect 35069 44211 35127 44217
rect 35250 44208 35256 44220
rect 35308 44208 35314 44260
rect 36538 44248 36544 44260
rect 36499 44220 36544 44248
rect 36538 44208 36544 44220
rect 36596 44208 36602 44260
rect 36633 44251 36691 44257
rect 36633 44217 36645 44251
rect 36679 44217 36691 44251
rect 37200 44248 37228 44424
rect 38565 44421 38577 44455
rect 38611 44452 38623 44455
rect 39942 44452 39948 44464
rect 38611 44424 39948 44452
rect 38611 44421 38623 44424
rect 38565 44415 38623 44421
rect 37826 44384 37832 44396
rect 37787 44356 37832 44384
rect 37826 44344 37832 44356
rect 37884 44344 37890 44396
rect 38562 44276 38568 44328
rect 38620 44316 38626 44328
rect 38657 44319 38715 44325
rect 38657 44316 38669 44319
rect 38620 44288 38669 44316
rect 38620 44276 38626 44288
rect 38657 44285 38669 44288
rect 38703 44285 38715 44319
rect 38657 44279 38715 44285
rect 39034 44257 39062 44424
rect 39942 44412 39948 44424
rect 40000 44452 40006 44464
rect 49510 44452 49516 44464
rect 40000 44424 49516 44452
rect 40000 44412 40006 44424
rect 49510 44412 49516 44424
rect 49568 44412 49574 44464
rect 41647 44387 41705 44393
rect 41647 44353 41659 44387
rect 41693 44384 41705 44387
rect 42613 44387 42671 44393
rect 42613 44384 42625 44387
rect 41693 44356 42625 44384
rect 41693 44353 41705 44356
rect 41647 44347 41705 44353
rect 42613 44353 42625 44356
rect 42659 44384 42671 44387
rect 42702 44384 42708 44396
rect 42659 44356 42708 44384
rect 42659 44353 42671 44356
rect 42613 44347 42671 44353
rect 42702 44344 42708 44356
rect 42760 44344 42766 44396
rect 43625 44387 43683 44393
rect 43625 44353 43637 44387
rect 43671 44384 43683 44387
rect 43806 44384 43812 44396
rect 43671 44356 43812 44384
rect 43671 44353 43683 44356
rect 43625 44347 43683 44353
rect 43806 44344 43812 44356
rect 43864 44344 43870 44396
rect 40564 44319 40622 44325
rect 40564 44316 40576 44319
rect 39132 44288 40576 44316
rect 39019 44251 39077 44257
rect 37200 44220 37872 44248
rect 36633 44211 36691 44217
rect 27062 44180 27068 44192
rect 25087 44152 25360 44180
rect 27023 44152 27068 44180
rect 25087 44149 25099 44152
rect 25041 44143 25099 44149
rect 27062 44140 27068 44152
rect 27120 44140 27126 44192
rect 27154 44140 27160 44192
rect 27212 44180 27218 44192
rect 28442 44180 28448 44192
rect 27212 44152 28448 44180
rect 27212 44140 27218 44152
rect 28442 44140 28448 44152
rect 28500 44180 28506 44192
rect 31665 44183 31723 44189
rect 31665 44180 31677 44183
rect 28500 44152 31677 44180
rect 28500 44140 28506 44152
rect 31665 44149 31677 44152
rect 31711 44149 31723 44183
rect 31665 44143 31723 44149
rect 35989 44183 36047 44189
rect 35989 44149 36001 44183
rect 36035 44180 36047 44183
rect 36357 44183 36415 44189
rect 36357 44180 36369 44183
rect 36035 44152 36369 44180
rect 36035 44149 36047 44152
rect 35989 44143 36047 44149
rect 36357 44149 36369 44152
rect 36403 44180 36415 44183
rect 36446 44180 36452 44192
rect 36403 44152 36452 44180
rect 36403 44149 36415 44152
rect 36357 44143 36415 44149
rect 36446 44140 36452 44152
rect 36504 44180 36510 44192
rect 36648 44180 36676 44211
rect 37844 44192 37872 44220
rect 39019 44217 39031 44251
rect 39065 44217 39077 44251
rect 39019 44211 39077 44217
rect 36504 44152 36676 44180
rect 36504 44140 36510 44152
rect 37826 44140 37832 44192
rect 37884 44180 37890 44192
rect 39132 44180 39160 44288
rect 40564 44285 40576 44288
rect 40610 44316 40622 44319
rect 40957 44319 41015 44325
rect 40957 44316 40969 44319
rect 40610 44288 40969 44316
rect 40610 44285 40622 44288
rect 40564 44279 40622 44285
rect 40957 44285 40969 44288
rect 41003 44285 41015 44319
rect 40957 44279 41015 44285
rect 41560 44319 41618 44325
rect 41560 44285 41572 44319
rect 41606 44285 41618 44319
rect 41560 44279 41618 44285
rect 43257 44319 43315 44325
rect 43257 44285 43269 44319
rect 43303 44316 43315 44319
rect 43714 44316 43720 44328
rect 43303 44288 43720 44316
rect 43303 44285 43315 44288
rect 43257 44279 43315 44285
rect 41322 44180 41328 44192
rect 37884 44152 39160 44180
rect 41283 44152 41328 44180
rect 37884 44140 37890 44152
rect 41322 44140 41328 44152
rect 41380 44140 41386 44192
rect 41575 44180 41603 44279
rect 43714 44276 43720 44288
rect 43772 44276 43778 44328
rect 44152 44319 44210 44325
rect 44152 44285 44164 44319
rect 44198 44316 44210 44319
rect 44266 44316 44272 44328
rect 44198 44288 44272 44316
rect 44198 44285 44210 44288
rect 44152 44279 44210 44285
rect 44266 44276 44272 44288
rect 44324 44316 44330 44328
rect 44545 44319 44603 44325
rect 44545 44316 44557 44319
rect 44324 44288 44557 44316
rect 44324 44276 44330 44288
rect 44545 44285 44557 44288
rect 44591 44285 44603 44319
rect 44545 44279 44603 44285
rect 42245 44251 42303 44257
rect 42245 44217 42257 44251
rect 42291 44248 42303 44251
rect 42682 44251 42740 44257
rect 42682 44248 42694 44251
rect 42291 44220 42694 44248
rect 42291 44217 42303 44220
rect 42245 44211 42303 44217
rect 42682 44217 42694 44220
rect 42728 44217 42740 44251
rect 42682 44211 42740 44217
rect 43438 44208 43444 44260
rect 43496 44248 43502 44260
rect 43901 44251 43959 44257
rect 43901 44248 43913 44251
rect 43496 44220 43913 44248
rect 43496 44208 43502 44220
rect 43901 44217 43913 44220
rect 43947 44217 43959 44251
rect 43901 44211 43959 44217
rect 42061 44183 42119 44189
rect 42061 44180 42073 44183
rect 41575 44152 42073 44180
rect 42061 44149 42073 44152
rect 42107 44180 42119 44183
rect 42150 44180 42156 44192
rect 42107 44152 42156 44180
rect 42107 44149 42119 44152
rect 42061 44143 42119 44149
rect 42150 44140 42156 44152
rect 42208 44140 42214 44192
rect 43622 44140 43628 44192
rect 43680 44180 43686 44192
rect 44223 44183 44281 44189
rect 44223 44180 44235 44183
rect 43680 44152 44235 44180
rect 43680 44140 43686 44152
rect 44223 44149 44235 44152
rect 44269 44149 44281 44183
rect 44223 44143 44281 44149
rect 1104 44090 48852 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 48852 44090
rect 1104 44016 48852 44038
rect 24995 43979 25053 43985
rect 24995 43945 25007 43979
rect 25041 43976 25053 43979
rect 25314 43976 25320 43988
rect 25041 43948 25320 43976
rect 25041 43945 25053 43948
rect 24995 43939 25053 43945
rect 25314 43936 25320 43948
rect 25372 43936 25378 43988
rect 25406 43936 25412 43988
rect 25464 43976 25470 43988
rect 27154 43976 27160 43988
rect 25464 43948 27160 43976
rect 25464 43936 25470 43948
rect 27154 43936 27160 43948
rect 27212 43936 27218 43988
rect 27430 43936 27436 43988
rect 27488 43976 27494 43988
rect 27709 43979 27767 43985
rect 27709 43976 27721 43979
rect 27488 43948 27721 43976
rect 27488 43936 27494 43948
rect 27709 43945 27721 43948
rect 27755 43945 27767 43979
rect 31294 43976 31300 43988
rect 27709 43939 27767 43945
rect 27816 43948 31300 43976
rect 19245 43911 19303 43917
rect 19245 43877 19257 43911
rect 19291 43908 19303 43911
rect 19334 43908 19340 43920
rect 19291 43880 19340 43908
rect 19291 43877 19303 43880
rect 19245 43871 19303 43877
rect 19334 43868 19340 43880
rect 19392 43868 19398 43920
rect 22005 43911 22063 43917
rect 22005 43877 22017 43911
rect 22051 43908 22063 43911
rect 22094 43908 22100 43920
rect 22051 43880 22100 43908
rect 22051 43877 22063 43880
rect 22005 43871 22063 43877
rect 22094 43868 22100 43880
rect 22152 43868 22158 43920
rect 25222 43868 25228 43920
rect 25280 43908 25286 43920
rect 25685 43911 25743 43917
rect 25685 43908 25697 43911
rect 25280 43880 25697 43908
rect 25280 43868 25286 43880
rect 25685 43877 25697 43880
rect 25731 43877 25743 43911
rect 27816 43908 27844 43948
rect 31294 43936 31300 43948
rect 31352 43936 31358 43988
rect 32122 43936 32128 43988
rect 32180 43976 32186 43988
rect 32309 43979 32367 43985
rect 32309 43976 32321 43979
rect 32180 43948 32321 43976
rect 32180 43936 32186 43948
rect 32309 43945 32321 43948
rect 32355 43945 32367 43979
rect 33410 43976 33416 43988
rect 33371 43948 33416 43976
rect 32309 43939 32367 43945
rect 28442 43908 28448 43920
rect 25685 43871 25743 43877
rect 26436 43880 27844 43908
rect 28403 43880 28448 43908
rect 24762 43800 24768 43852
rect 24820 43840 24826 43852
rect 24924 43843 24982 43849
rect 24924 43840 24936 43843
rect 24820 43812 24936 43840
rect 24820 43800 24826 43812
rect 24924 43809 24936 43812
rect 24970 43840 24982 43843
rect 25314 43840 25320 43852
rect 24970 43812 25320 43840
rect 24970 43809 24982 43812
rect 24924 43803 24982 43809
rect 25314 43800 25320 43812
rect 25372 43840 25378 43852
rect 26436 43840 26464 43880
rect 28442 43868 28448 43880
rect 28500 43868 28506 43920
rect 28994 43908 29000 43920
rect 28955 43880 29000 43908
rect 28994 43868 29000 43880
rect 29052 43908 29058 43920
rect 29273 43911 29331 43917
rect 29273 43908 29285 43911
rect 29052 43880 29285 43908
rect 29052 43868 29058 43880
rect 29273 43877 29285 43880
rect 29319 43877 29331 43911
rect 29273 43871 29331 43877
rect 30190 43868 30196 43920
rect 30248 43908 30254 43920
rect 30330 43911 30388 43917
rect 30330 43908 30342 43911
rect 30248 43880 30342 43908
rect 30248 43868 30254 43880
rect 30330 43877 30342 43880
rect 30376 43877 30388 43911
rect 30330 43871 30388 43877
rect 25372 43812 26464 43840
rect 25372 43800 25378 43812
rect 26786 43800 26792 43852
rect 26844 43840 26850 43852
rect 26916 43843 26974 43849
rect 26916 43840 26928 43843
rect 26844 43812 26928 43840
rect 26844 43800 26850 43812
rect 26916 43809 26928 43812
rect 26962 43809 26974 43843
rect 27430 43840 27436 43852
rect 27343 43812 27436 43840
rect 26916 43803 26974 43809
rect 27430 43800 27436 43812
rect 27488 43840 27494 43852
rect 27614 43840 27620 43852
rect 27488 43812 27620 43840
rect 27488 43800 27494 43812
rect 27614 43800 27620 43812
rect 27672 43800 27678 43852
rect 30009 43843 30067 43849
rect 30009 43809 30021 43843
rect 30055 43840 30067 43843
rect 30742 43840 30748 43852
rect 30055 43812 30748 43840
rect 30055 43809 30067 43812
rect 30009 43803 30067 43809
rect 30742 43800 30748 43812
rect 30800 43800 30806 43852
rect 19150 43772 19156 43784
rect 19111 43744 19156 43772
rect 19150 43732 19156 43744
rect 19208 43732 19214 43784
rect 21910 43772 21916 43784
rect 21871 43744 21916 43772
rect 21910 43732 21916 43744
rect 21968 43732 21974 43784
rect 22557 43775 22615 43781
rect 22557 43741 22569 43775
rect 22603 43772 22615 43775
rect 23382 43772 23388 43784
rect 22603 43744 23388 43772
rect 22603 43741 22615 43744
rect 22557 43735 22615 43741
rect 18046 43664 18052 43716
rect 18104 43704 18110 43716
rect 19705 43707 19763 43713
rect 19705 43704 19717 43707
rect 18104 43676 19717 43704
rect 18104 43664 18110 43676
rect 19705 43673 19717 43676
rect 19751 43704 19763 43707
rect 22572 43704 22600 43735
rect 23382 43732 23388 43744
rect 23440 43732 23446 43784
rect 28350 43772 28356 43784
rect 28311 43744 28356 43772
rect 28350 43732 28356 43744
rect 28408 43732 28414 43784
rect 19751 43676 22600 43704
rect 32324 43704 32352 43939
rect 33410 43936 33416 43948
rect 33468 43936 33474 43988
rect 34931 43979 34989 43985
rect 34931 43945 34943 43979
rect 34977 43976 34989 43979
rect 35342 43976 35348 43988
rect 34977 43948 35348 43976
rect 34977 43945 34989 43948
rect 34931 43939 34989 43945
rect 35342 43936 35348 43948
rect 35400 43936 35406 43988
rect 36081 43979 36139 43985
rect 36081 43945 36093 43979
rect 36127 43976 36139 43979
rect 36170 43976 36176 43988
rect 36127 43948 36176 43976
rect 36127 43945 36139 43948
rect 36081 43939 36139 43945
rect 36170 43936 36176 43948
rect 36228 43936 36234 43988
rect 40037 43979 40095 43985
rect 40037 43945 40049 43979
rect 40083 43976 40095 43979
rect 41322 43976 41328 43988
rect 40083 43948 41328 43976
rect 40083 43945 40095 43948
rect 40037 43939 40095 43945
rect 41322 43936 41328 43948
rect 41380 43936 41386 43988
rect 42702 43976 42708 43988
rect 42663 43948 42708 43976
rect 42702 43936 42708 43948
rect 42760 43936 42766 43988
rect 35250 43908 35256 43920
rect 35211 43880 35256 43908
rect 35250 43868 35256 43880
rect 35308 43868 35314 43920
rect 39209 43911 39267 43917
rect 39209 43877 39221 43911
rect 39255 43908 39267 43911
rect 39298 43908 39304 43920
rect 39255 43880 39304 43908
rect 39255 43877 39267 43880
rect 39209 43871 39267 43877
rect 39298 43868 39304 43880
rect 39356 43908 39362 43920
rect 39485 43911 39543 43917
rect 39485 43908 39497 43911
rect 39356 43880 39497 43908
rect 39356 43868 39362 43880
rect 39485 43877 39497 43880
rect 39531 43877 39543 43911
rect 39485 43871 39543 43877
rect 42383 43911 42441 43917
rect 42383 43877 42395 43911
rect 42429 43908 42441 43911
rect 43438 43908 43444 43920
rect 42429 43880 43444 43908
rect 42429 43877 42441 43880
rect 42383 43871 42441 43877
rect 43438 43868 43444 43880
rect 43496 43868 43502 43920
rect 43533 43911 43591 43917
rect 43533 43877 43545 43911
rect 43579 43908 43591 43911
rect 43806 43908 43812 43920
rect 43579 43880 43812 43908
rect 43579 43877 43591 43880
rect 43533 43871 43591 43877
rect 43806 43868 43812 43880
rect 43864 43908 43870 43920
rect 44082 43908 44088 43920
rect 43864 43880 44088 43908
rect 43864 43868 43870 43880
rect 44082 43868 44088 43880
rect 44140 43868 44146 43920
rect 34698 43800 34704 43852
rect 34756 43840 34762 43852
rect 34828 43843 34886 43849
rect 34828 43840 34840 43843
rect 34756 43812 34840 43840
rect 34756 43800 34762 43812
rect 34828 43809 34840 43812
rect 34874 43809 34886 43843
rect 36170 43840 36176 43852
rect 36131 43812 36176 43840
rect 34828 43803 34886 43809
rect 36170 43800 36176 43812
rect 36228 43800 36234 43852
rect 36311 43843 36369 43849
rect 36311 43809 36323 43843
rect 36357 43840 36369 43843
rect 36538 43840 36544 43852
rect 36357 43812 36544 43840
rect 36357 43809 36369 43812
rect 36311 43803 36369 43809
rect 36538 43800 36544 43812
rect 36596 43840 36602 43852
rect 37001 43843 37059 43849
rect 37001 43840 37013 43843
rect 36596 43812 37013 43840
rect 36596 43800 36602 43812
rect 37001 43809 37013 43812
rect 37047 43809 37059 43843
rect 37001 43803 37059 43809
rect 38473 43843 38531 43849
rect 38473 43809 38485 43843
rect 38519 43809 38531 43843
rect 38930 43840 38936 43852
rect 38891 43812 38936 43840
rect 38473 43803 38531 43809
rect 33042 43772 33048 43784
rect 33003 43744 33048 43772
rect 33042 43732 33048 43744
rect 33100 43732 33106 43784
rect 38378 43704 38384 43716
rect 32324 43676 38384 43704
rect 19751 43673 19763 43676
rect 19705 43667 19763 43673
rect 38378 43664 38384 43676
rect 38436 43704 38442 43716
rect 38488 43704 38516 43803
rect 38930 43800 38936 43812
rect 38988 43800 38994 43852
rect 41046 43840 41052 43852
rect 41007 43812 41052 43840
rect 41046 43800 41052 43812
rect 41104 43800 41110 43852
rect 42280 43843 42338 43849
rect 42280 43840 42292 43843
rect 41892 43812 42292 43840
rect 41892 43784 41920 43812
rect 42280 43809 42292 43812
rect 42326 43840 42338 43843
rect 42518 43840 42524 43852
rect 42326 43812 42524 43840
rect 42326 43809 42338 43812
rect 42280 43803 42338 43809
rect 42518 43800 42524 43812
rect 42576 43800 42582 43852
rect 41874 43732 41880 43784
rect 41932 43732 41938 43784
rect 43441 43775 43499 43781
rect 43441 43741 43453 43775
rect 43487 43772 43499 43775
rect 43622 43772 43628 43784
rect 43487 43744 43628 43772
rect 43487 43741 43499 43744
rect 43441 43735 43499 43741
rect 43622 43732 43628 43744
rect 43680 43732 43686 43784
rect 43714 43732 43720 43784
rect 43772 43772 43778 43784
rect 43772 43744 43817 43772
rect 43772 43732 43778 43744
rect 38436 43676 38516 43704
rect 38436 43664 38442 43676
rect 42150 43664 42156 43716
rect 42208 43704 42214 43716
rect 42702 43704 42708 43716
rect 42208 43676 42708 43704
rect 42208 43664 42214 43676
rect 42702 43664 42708 43676
rect 42760 43664 42766 43716
rect 16482 43636 16488 43648
rect 16443 43608 16488 43636
rect 16482 43596 16488 43608
rect 16540 43596 16546 43648
rect 26602 43596 26608 43648
rect 26660 43636 26666 43648
rect 27019 43639 27077 43645
rect 27019 43636 27031 43639
rect 26660 43608 27031 43636
rect 26660 43596 26666 43608
rect 27019 43605 27031 43608
rect 27065 43605 27077 43639
rect 30926 43636 30932 43648
rect 30887 43608 30932 43636
rect 27019 43599 27077 43605
rect 30926 43596 30932 43608
rect 30984 43596 30990 43648
rect 31202 43636 31208 43648
rect 31163 43608 31208 43636
rect 31202 43596 31208 43608
rect 31260 43596 31266 43648
rect 33965 43639 34023 43645
rect 33965 43605 33977 43639
rect 34011 43636 34023 43639
rect 34238 43636 34244 43648
rect 34011 43608 34244 43636
rect 34011 43605 34023 43608
rect 33965 43599 34023 43605
rect 34238 43596 34244 43608
rect 34296 43596 34302 43648
rect 36630 43636 36636 43648
rect 36591 43608 36636 43636
rect 36630 43596 36636 43608
rect 36688 43596 36694 43648
rect 41187 43639 41245 43645
rect 41187 43605 41199 43639
rect 41233 43636 41245 43639
rect 41693 43639 41751 43645
rect 41693 43636 41705 43639
rect 41233 43608 41705 43636
rect 41233 43605 41245 43608
rect 41187 43599 41245 43605
rect 41693 43605 41705 43608
rect 41739 43636 41751 43639
rect 41782 43636 41788 43648
rect 41739 43608 41788 43636
rect 41739 43605 41751 43608
rect 41693 43599 41751 43605
rect 41782 43596 41788 43608
rect 41840 43596 41846 43648
rect 1104 43546 48852 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 48852 43546
rect 1104 43472 48852 43494
rect 19150 43392 19156 43444
rect 19208 43432 19214 43444
rect 20441 43435 20499 43441
rect 20441 43432 20453 43435
rect 19208 43404 20453 43432
rect 19208 43392 19214 43404
rect 20441 43401 20453 43404
rect 20487 43401 20499 43435
rect 20441 43395 20499 43401
rect 21361 43435 21419 43441
rect 21361 43401 21373 43435
rect 21407 43432 21419 43435
rect 24762 43432 24768 43444
rect 21407 43404 24768 43432
rect 21407 43401 21419 43404
rect 21361 43395 21419 43401
rect 17037 43367 17095 43373
rect 17037 43333 17049 43367
rect 17083 43364 17095 43367
rect 18046 43364 18052 43376
rect 17083 43336 18052 43364
rect 17083 43333 17095 43336
rect 17037 43327 17095 43333
rect 18046 43324 18052 43336
rect 18104 43324 18110 43376
rect 16482 43296 16488 43308
rect 16443 43268 16488 43296
rect 16482 43256 16488 43268
rect 16540 43256 16546 43308
rect 17218 43256 17224 43308
rect 17276 43296 17282 43308
rect 19429 43299 19487 43305
rect 19429 43296 19441 43299
rect 17276 43268 19441 43296
rect 17276 43256 17282 43268
rect 19429 43265 19441 43268
rect 19475 43296 19487 43299
rect 19475 43268 20576 43296
rect 19475 43265 19487 43268
rect 19429 43259 19487 43265
rect 18116 43231 18174 43237
rect 18116 43197 18128 43231
rect 18162 43228 18174 43231
rect 18162 43200 18644 43228
rect 18162 43197 18174 43200
rect 18116 43191 18174 43197
rect 16301 43163 16359 43169
rect 16301 43129 16313 43163
rect 16347 43160 16359 43163
rect 16574 43160 16580 43172
rect 16347 43132 16580 43160
rect 16347 43129 16359 43132
rect 16301 43123 16359 43129
rect 16574 43120 16580 43132
rect 16632 43120 16638 43172
rect 18616 43104 18644 43200
rect 18966 43120 18972 43172
rect 19024 43160 19030 43172
rect 19142 43163 19200 43169
rect 19142 43160 19154 43163
rect 19024 43132 19154 43160
rect 19024 43120 19030 43132
rect 19142 43129 19154 43132
rect 19188 43129 19200 43163
rect 19142 43123 19200 43129
rect 19245 43163 19303 43169
rect 19245 43129 19257 43163
rect 19291 43129 19303 43163
rect 20548 43160 20576 43268
rect 20876 43231 20934 43237
rect 20876 43197 20888 43231
rect 20922 43228 20934 43231
rect 21376 43228 21404 43395
rect 24762 43392 24768 43404
rect 24820 43392 24826 43444
rect 26602 43432 26608 43444
rect 26563 43404 26608 43432
rect 26602 43392 26608 43404
rect 26660 43392 26666 43444
rect 28350 43392 28356 43444
rect 28408 43432 28414 43444
rect 28626 43432 28632 43444
rect 28408 43404 28632 43432
rect 28408 43392 28414 43404
rect 28626 43392 28632 43404
rect 28684 43392 28690 43444
rect 30742 43432 30748 43444
rect 30703 43404 30748 43432
rect 30742 43392 30748 43404
rect 30800 43392 30806 43444
rect 34238 43432 34244 43444
rect 34199 43404 34244 43432
rect 34238 43392 34244 43404
rect 34296 43392 34302 43444
rect 34698 43432 34704 43444
rect 34659 43404 34704 43432
rect 34698 43392 34704 43404
rect 34756 43392 34762 43444
rect 36170 43392 36176 43444
rect 36228 43432 36234 43444
rect 36265 43435 36323 43441
rect 36265 43432 36277 43435
rect 36228 43404 36277 43432
rect 36228 43392 36234 43404
rect 36265 43401 36277 43404
rect 36311 43432 36323 43435
rect 42150 43432 42156 43444
rect 36311 43404 42156 43432
rect 36311 43401 36323 43404
rect 36265 43395 36323 43401
rect 42150 43392 42156 43404
rect 42208 43392 42214 43444
rect 43165 43435 43223 43441
rect 43165 43401 43177 43435
rect 43211 43432 43223 43435
rect 43622 43432 43628 43444
rect 43211 43404 43628 43432
rect 43211 43401 43223 43404
rect 43165 43395 43223 43401
rect 43622 43392 43628 43404
rect 43680 43392 43686 43444
rect 44082 43432 44088 43444
rect 44043 43404 44088 43432
rect 44082 43392 44088 43404
rect 44140 43392 44146 43444
rect 21910 43324 21916 43376
rect 21968 43364 21974 43376
rect 23201 43367 23259 43373
rect 23201 43364 23213 43367
rect 21968 43336 23213 43364
rect 21968 43324 21974 43336
rect 23201 43333 23213 43336
rect 23247 43333 23259 43367
rect 23201 43327 23259 43333
rect 22189 43299 22247 43305
rect 22189 43296 22201 43299
rect 20922 43200 21404 43228
rect 21468 43268 22201 43296
rect 20922 43197 20934 43200
rect 20876 43191 20934 43197
rect 21468 43160 21496 43268
rect 22189 43265 22201 43268
rect 22235 43296 22247 43299
rect 22370 43296 22376 43308
rect 22235 43268 22376 43296
rect 22235 43265 22247 43268
rect 22189 43259 22247 43265
rect 22370 43256 22376 43268
rect 22428 43256 22434 43308
rect 26620 43296 26648 43392
rect 30374 43324 30380 43376
rect 30432 43364 30438 43376
rect 32125 43367 32183 43373
rect 32125 43364 32137 43367
rect 30432 43336 32137 43364
rect 30432 43324 30438 43336
rect 32125 43333 32137 43336
rect 32171 43364 32183 43367
rect 37458 43364 37464 43376
rect 32171 43336 37464 43364
rect 32171 43333 32183 43336
rect 32125 43327 32183 43333
rect 27341 43299 27399 43305
rect 27341 43296 27353 43299
rect 26620 43268 27353 43296
rect 27341 43265 27353 43268
rect 27387 43265 27399 43299
rect 27614 43296 27620 43308
rect 27575 43268 27620 43296
rect 27341 43259 27399 43265
rect 27614 43256 27620 43268
rect 27672 43256 27678 43308
rect 28353 43299 28411 43305
rect 28353 43265 28365 43299
rect 28399 43296 28411 43299
rect 28442 43296 28448 43308
rect 28399 43268 28448 43296
rect 28399 43265 28411 43268
rect 28353 43259 28411 43265
rect 28442 43256 28448 43268
rect 28500 43256 28506 43308
rect 28994 43256 29000 43308
rect 29052 43296 29058 43308
rect 29365 43299 29423 43305
rect 29365 43296 29377 43299
rect 29052 43268 29377 43296
rect 29052 43256 29058 43268
rect 29365 43265 29377 43268
rect 29411 43265 29423 43299
rect 29638 43296 29644 43308
rect 29599 43268 29644 43296
rect 29365 43259 29423 43265
rect 29638 43256 29644 43268
rect 29696 43256 29702 43308
rect 23912 43231 23970 43237
rect 23912 43197 23924 43231
rect 23958 43228 23970 43231
rect 23958 43200 24440 43228
rect 23958 43197 23970 43200
rect 23912 43191 23970 43197
rect 20548 43132 21496 43160
rect 19245 43123 19303 43129
rect 18187 43095 18245 43101
rect 18187 43061 18199 43095
rect 18233 43092 18245 43095
rect 18414 43092 18420 43104
rect 18233 43064 18420 43092
rect 18233 43061 18245 43064
rect 18187 43055 18245 43061
rect 18414 43052 18420 43064
rect 18472 43052 18478 43104
rect 18598 43092 18604 43104
rect 18559 43064 18604 43092
rect 18598 43052 18604 43064
rect 18656 43052 18662 43104
rect 18874 43092 18880 43104
rect 18835 43064 18880 43092
rect 18874 43052 18880 43064
rect 18932 43092 18938 43104
rect 19260 43092 19288 43123
rect 21726 43120 21732 43172
rect 21784 43160 21790 43172
rect 21913 43163 21971 43169
rect 21913 43160 21925 43163
rect 21784 43132 21925 43160
rect 21784 43120 21790 43132
rect 21913 43129 21925 43132
rect 21959 43129 21971 43163
rect 21913 43123 21971 43129
rect 22005 43163 22063 43169
rect 22005 43129 22017 43163
rect 22051 43160 22063 43163
rect 22094 43160 22100 43172
rect 22051 43132 22100 43160
rect 22051 43129 22063 43132
rect 22005 43123 22063 43129
rect 20073 43095 20131 43101
rect 20073 43092 20085 43095
rect 18932 43064 20085 43092
rect 18932 43052 18938 43064
rect 20073 43061 20085 43064
rect 20119 43061 20131 43095
rect 20073 43055 20131 43061
rect 20947 43095 21005 43101
rect 20947 43061 20959 43095
rect 20993 43092 21005 43095
rect 21174 43092 21180 43104
rect 20993 43064 21180 43092
rect 20993 43061 21005 43064
rect 20947 43055 21005 43061
rect 21174 43052 21180 43064
rect 21232 43052 21238 43104
rect 21637 43095 21695 43101
rect 21637 43061 21649 43095
rect 21683 43092 21695 43095
rect 22020 43092 22048 43123
rect 22094 43120 22100 43132
rect 22152 43120 22158 43172
rect 22922 43092 22928 43104
rect 21683 43064 22048 43092
rect 22883 43064 22928 43092
rect 21683 43061 21695 43064
rect 21637 43055 21695 43061
rect 22922 43052 22928 43064
rect 22980 43052 22986 43104
rect 23983 43095 24041 43101
rect 23983 43061 23995 43095
rect 24029 43092 24041 43095
rect 24210 43092 24216 43104
rect 24029 43064 24216 43092
rect 24029 43061 24041 43064
rect 23983 43055 24041 43061
rect 24210 43052 24216 43064
rect 24268 43052 24274 43104
rect 24412 43101 24440 43200
rect 32030 43188 32036 43240
rect 32088 43228 32094 43240
rect 32140 43228 32168 43327
rect 37458 43324 37464 43336
rect 37516 43364 37522 43376
rect 38197 43367 38255 43373
rect 38197 43364 38209 43367
rect 37516 43336 38209 43364
rect 37516 43324 37522 43336
rect 38197 43333 38209 43336
rect 38243 43333 38255 43367
rect 38197 43327 38255 43333
rect 32214 43256 32220 43308
rect 32272 43296 32278 43308
rect 33042 43296 33048 43308
rect 32272 43268 32812 43296
rect 32955 43268 33048 43296
rect 32272 43256 32278 43268
rect 32784 43237 32812 43268
rect 33042 43256 33048 43268
rect 33100 43296 33106 43308
rect 33689 43299 33747 43305
rect 33689 43296 33701 43299
rect 33100 43268 33701 43296
rect 33100 43256 33106 43268
rect 33689 43265 33701 43268
rect 33735 43265 33747 43299
rect 35342 43296 35348 43308
rect 35303 43268 35348 43296
rect 33689 43259 33747 43265
rect 35342 43256 35348 43268
rect 35400 43256 35406 43308
rect 36814 43296 36820 43308
rect 36775 43268 36820 43296
rect 36814 43256 36820 43268
rect 36872 43256 36878 43308
rect 32309 43231 32367 43237
rect 32309 43228 32321 43231
rect 32088 43200 32321 43228
rect 32088 43188 32094 43200
rect 32309 43197 32321 43200
rect 32355 43197 32367 43231
rect 32309 43191 32367 43197
rect 32769 43231 32827 43237
rect 32769 43197 32781 43231
rect 32815 43197 32827 43231
rect 38212 43228 38240 43327
rect 39758 43256 39764 43308
rect 39816 43296 39822 43308
rect 41046 43296 41052 43308
rect 39816 43268 41052 43296
rect 39816 43256 39822 43268
rect 41046 43256 41052 43268
rect 41104 43256 41110 43308
rect 41782 43296 41788 43308
rect 41743 43268 41788 43296
rect 41782 43256 41788 43268
rect 41840 43256 41846 43308
rect 38381 43231 38439 43237
rect 38381 43228 38393 43231
rect 38212 43200 38393 43228
rect 32769 43191 32827 43197
rect 38381 43197 38393 43200
rect 38427 43197 38439 43231
rect 38930 43228 38936 43240
rect 38891 43200 38936 43228
rect 38381 43191 38439 43197
rect 38930 43188 38936 43200
rect 38988 43188 38994 43240
rect 40532 43231 40590 43237
rect 40532 43228 40544 43231
rect 40236 43200 40544 43228
rect 24762 43120 24768 43172
rect 24820 43160 24826 43172
rect 24949 43163 25007 43169
rect 24949 43160 24961 43163
rect 24820 43132 24961 43160
rect 24820 43120 24826 43132
rect 24949 43129 24961 43132
rect 24995 43129 25007 43163
rect 24949 43123 25007 43129
rect 25041 43163 25099 43169
rect 25041 43129 25053 43163
rect 25087 43129 25099 43163
rect 25590 43160 25596 43172
rect 25551 43132 25596 43160
rect 25041 43123 25099 43129
rect 24397 43095 24455 43101
rect 24397 43061 24409 43095
rect 24443 43092 24455 43095
rect 24486 43092 24492 43104
rect 24443 43064 24492 43092
rect 24443 43061 24455 43064
rect 24397 43055 24455 43061
rect 24486 43052 24492 43064
rect 24544 43052 24550 43104
rect 25056 43092 25084 43123
rect 25590 43120 25596 43132
rect 25648 43120 25654 43172
rect 27430 43160 27436 43172
rect 27391 43132 27436 43160
rect 27430 43120 27436 43132
rect 27488 43120 27494 43172
rect 29457 43163 29515 43169
rect 29457 43129 29469 43163
rect 29503 43160 29515 43163
rect 30926 43160 30932 43172
rect 29503 43132 30932 43160
rect 29503 43129 29515 43132
rect 29457 43123 29515 43129
rect 25958 43092 25964 43104
rect 25056 43064 25964 43092
rect 25958 43052 25964 43064
rect 26016 43052 26022 43104
rect 26786 43052 26792 43104
rect 26844 43092 26850 43104
rect 26881 43095 26939 43101
rect 26881 43092 26893 43095
rect 26844 43064 26893 43092
rect 26844 43052 26850 43064
rect 26881 43061 26893 43064
rect 26927 43061 26939 43095
rect 26881 43055 26939 43061
rect 29089 43095 29147 43101
rect 29089 43061 29101 43095
rect 29135 43092 29147 43095
rect 29472 43092 29500 43123
rect 30926 43120 30932 43132
rect 30984 43120 30990 43172
rect 34974 43160 34980 43172
rect 34935 43132 34980 43160
rect 34974 43120 34980 43132
rect 35032 43120 35038 43172
rect 35069 43163 35127 43169
rect 35069 43129 35081 43163
rect 35115 43129 35127 43163
rect 36538 43160 36544 43172
rect 36499 43132 36544 43160
rect 35069 43123 35127 43129
rect 29135 43064 29500 43092
rect 29135 43061 29147 43064
rect 29089 43055 29147 43061
rect 30190 43052 30196 43104
rect 30248 43092 30254 43104
rect 30285 43095 30343 43101
rect 30285 43092 30297 43095
rect 30248 43064 30297 43092
rect 30248 43052 30254 43064
rect 30285 43061 30297 43064
rect 30331 43061 30343 43095
rect 30285 43055 30343 43061
rect 33042 43052 33048 43104
rect 33100 43092 33106 43104
rect 33321 43095 33379 43101
rect 33321 43092 33333 43095
rect 33100 43064 33333 43092
rect 33100 43052 33106 43064
rect 33321 43061 33333 43064
rect 33367 43092 33379 43095
rect 33410 43092 33416 43104
rect 33367 43064 33416 43092
rect 33367 43061 33379 43064
rect 33321 43055 33379 43061
rect 33410 43052 33416 43064
rect 33468 43052 33474 43104
rect 34238 43052 34244 43104
rect 34296 43092 34302 43104
rect 35084 43092 35112 43123
rect 36538 43120 36544 43132
rect 36596 43120 36602 43172
rect 36630 43120 36636 43172
rect 36688 43160 36694 43172
rect 36688 43132 36733 43160
rect 36688 43120 36694 43132
rect 34296 43064 35112 43092
rect 37553 43095 37611 43101
rect 34296 43052 34302 43064
rect 37553 43061 37565 43095
rect 37599 43092 37611 43095
rect 37829 43095 37887 43101
rect 37829 43092 37841 43095
rect 37599 43064 37841 43092
rect 37599 43061 37611 43064
rect 37553 43055 37611 43061
rect 37829 43061 37841 43064
rect 37875 43092 37887 43095
rect 38102 43092 38108 43104
rect 37875 43064 38108 43092
rect 37875 43061 37887 43064
rect 37829 43055 37887 43061
rect 38102 43052 38108 43064
rect 38160 43052 38166 43104
rect 38470 43092 38476 43104
rect 38431 43064 38476 43092
rect 38470 43052 38476 43064
rect 38528 43052 38534 43104
rect 39482 43052 39488 43104
rect 39540 43092 39546 43104
rect 40236 43101 40264 43200
rect 40532 43197 40544 43200
rect 40578 43197 40590 43231
rect 40532 43191 40590 43197
rect 42610 43188 42616 43240
rect 42668 43228 42674 43240
rect 43324 43231 43382 43237
rect 43324 43228 43336 43231
rect 42668 43200 43336 43228
rect 42668 43188 42674 43200
rect 43324 43197 43336 43200
rect 43370 43228 43382 43231
rect 43717 43231 43775 43237
rect 43717 43228 43729 43231
rect 43370 43200 43729 43228
rect 43370 43197 43382 43200
rect 43324 43191 43382 43197
rect 43717 43197 43729 43200
rect 43763 43197 43775 43231
rect 43717 43191 43775 43197
rect 41601 43163 41659 43169
rect 41601 43129 41613 43163
rect 41647 43160 41659 43163
rect 41877 43163 41935 43169
rect 41877 43160 41889 43163
rect 41647 43132 41889 43160
rect 41647 43129 41659 43132
rect 41601 43123 41659 43129
rect 41877 43129 41889 43132
rect 41923 43160 41935 43163
rect 42058 43160 42064 43172
rect 41923 43132 42064 43160
rect 41923 43129 41935 43132
rect 41877 43123 41935 43129
rect 42058 43120 42064 43132
rect 42116 43120 42122 43172
rect 42429 43163 42487 43169
rect 42429 43129 42441 43163
rect 42475 43129 42487 43163
rect 42429 43123 42487 43129
rect 40221 43095 40279 43101
rect 40221 43092 40233 43095
rect 39540 43064 40233 43092
rect 39540 43052 39546 43064
rect 40221 43061 40233 43064
rect 40267 43061 40279 43095
rect 40221 43055 40279 43061
rect 40635 43095 40693 43101
rect 40635 43061 40647 43095
rect 40681 43092 40693 43095
rect 40862 43092 40868 43104
rect 40681 43064 40868 43092
rect 40681 43061 40693 43064
rect 40635 43055 40693 43061
rect 40862 43052 40868 43064
rect 40920 43052 40926 43104
rect 41782 43052 41788 43104
rect 41840 43092 41846 43104
rect 42334 43092 42340 43104
rect 41840 43064 42340 43092
rect 41840 43052 41846 43064
rect 42334 43052 42340 43064
rect 42392 43092 42398 43104
rect 42444 43092 42472 43123
rect 42518 43120 42524 43172
rect 42576 43160 42582 43172
rect 42797 43163 42855 43169
rect 42797 43160 42809 43163
rect 42576 43132 42809 43160
rect 42576 43120 42582 43132
rect 42797 43129 42809 43132
rect 42843 43160 42855 43163
rect 43990 43160 43996 43172
rect 42843 43132 43996 43160
rect 42843 43129 42855 43132
rect 42797 43123 42855 43129
rect 43990 43120 43996 43132
rect 44048 43120 44054 43172
rect 42392 43064 42472 43092
rect 43395 43095 43453 43101
rect 42392 43052 42398 43064
rect 43395 43061 43407 43095
rect 43441 43092 43453 43095
rect 43530 43092 43536 43104
rect 43441 43064 43536 43092
rect 43441 43061 43453 43064
rect 43395 43055 43453 43061
rect 43530 43052 43536 43064
rect 43588 43052 43594 43104
rect 1104 43002 48852 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 48852 43002
rect 1104 42928 48852 42950
rect 15519 42891 15577 42897
rect 15519 42857 15531 42891
rect 15565 42888 15577 42891
rect 16482 42888 16488 42900
rect 15565 42860 16488 42888
rect 15565 42857 15577 42860
rect 15519 42851 15577 42857
rect 16482 42848 16488 42860
rect 16540 42848 16546 42900
rect 18414 42848 18420 42900
rect 18472 42888 18478 42900
rect 18966 42888 18972 42900
rect 18472 42860 18972 42888
rect 18472 42848 18478 42860
rect 18966 42848 18972 42860
rect 19024 42848 19030 42900
rect 21039 42891 21097 42897
rect 21039 42857 21051 42891
rect 21085 42888 21097 42891
rect 21910 42888 21916 42900
rect 21085 42860 21916 42888
rect 21085 42857 21097 42860
rect 21039 42851 21097 42857
rect 21910 42848 21916 42860
rect 21968 42848 21974 42900
rect 23983 42891 24041 42897
rect 23983 42857 23995 42891
rect 24029 42888 24041 42891
rect 24762 42888 24768 42900
rect 24029 42860 24768 42888
rect 24029 42857 24041 42860
rect 23983 42851 24041 42857
rect 24762 42848 24768 42860
rect 24820 42848 24826 42900
rect 26878 42888 26884 42900
rect 26839 42860 26884 42888
rect 26878 42848 26884 42860
rect 26936 42848 26942 42900
rect 32214 42848 32220 42900
rect 32272 42888 32278 42900
rect 32309 42891 32367 42897
rect 32309 42888 32321 42891
rect 32272 42860 32321 42888
rect 32272 42848 32278 42860
rect 32309 42857 32321 42860
rect 32355 42857 32367 42891
rect 33042 42888 33048 42900
rect 33003 42860 33048 42888
rect 32309 42851 32367 42857
rect 33042 42848 33048 42860
rect 33100 42848 33106 42900
rect 33597 42891 33655 42897
rect 33597 42857 33609 42891
rect 33643 42888 33655 42891
rect 33643 42860 34836 42888
rect 33643 42857 33655 42860
rect 33597 42851 33655 42857
rect 34808 42832 34836 42860
rect 36538 42848 36544 42900
rect 36596 42888 36602 42900
rect 36817 42891 36875 42897
rect 36817 42888 36829 42891
rect 36596 42860 36829 42888
rect 36596 42848 36602 42860
rect 36817 42857 36829 42860
rect 36863 42888 36875 42891
rect 37875 42891 37933 42897
rect 37875 42888 37887 42891
rect 36863 42860 37887 42888
rect 36863 42857 36875 42860
rect 36817 42851 36875 42857
rect 37875 42857 37887 42860
rect 37921 42857 37933 42891
rect 37875 42851 37933 42857
rect 38194 42848 38200 42900
rect 38252 42888 38258 42900
rect 40770 42888 40776 42900
rect 38252 42860 39614 42888
rect 40683 42860 40776 42888
rect 38252 42848 38258 42860
rect 16298 42780 16304 42832
rect 16356 42820 16362 42832
rect 16574 42820 16580 42832
rect 16356 42792 16580 42820
rect 16356 42780 16362 42792
rect 16574 42780 16580 42792
rect 16632 42780 16638 42832
rect 18874 42780 18880 42832
rect 18932 42820 18938 42832
rect 19242 42820 19248 42832
rect 18932 42792 19248 42820
rect 18932 42780 18938 42792
rect 19242 42780 19248 42792
rect 19300 42780 19306 42832
rect 19426 42780 19432 42832
rect 19484 42820 19490 42832
rect 19484 42792 20979 42820
rect 19484 42780 19490 42792
rect 15448 42755 15506 42761
rect 15448 42721 15460 42755
rect 15494 42752 15506 42755
rect 15930 42752 15936 42764
rect 15494 42724 15936 42752
rect 15494 42721 15506 42724
rect 15448 42715 15506 42721
rect 15930 42712 15936 42724
rect 15988 42712 15994 42764
rect 18100 42755 18158 42761
rect 18100 42721 18112 42755
rect 18146 42752 18158 42755
rect 18966 42752 18972 42764
rect 18146 42724 18972 42752
rect 18146 42721 18158 42724
rect 18100 42715 18158 42721
rect 18966 42712 18972 42724
rect 19024 42712 19030 42764
rect 20951 42761 20979 42792
rect 21174 42780 21180 42832
rect 21232 42820 21238 42832
rect 21818 42820 21824 42832
rect 21232 42792 21824 42820
rect 21232 42780 21238 42792
rect 21818 42780 21824 42792
rect 21876 42820 21882 42832
rect 22005 42823 22063 42829
rect 22005 42820 22017 42823
rect 21876 42792 22017 42820
rect 21876 42780 21882 42792
rect 22005 42789 22017 42792
rect 22051 42789 22063 42823
rect 22005 42783 22063 42789
rect 22094 42780 22100 42832
rect 22152 42820 22158 42832
rect 22922 42820 22928 42832
rect 22152 42792 22928 42820
rect 22152 42780 22158 42792
rect 22922 42780 22928 42792
rect 22980 42780 22986 42832
rect 24946 42780 24952 42832
rect 25004 42820 25010 42832
rect 25041 42823 25099 42829
rect 25041 42820 25053 42823
rect 25004 42792 25053 42820
rect 25004 42780 25010 42792
rect 25041 42789 25053 42792
rect 25087 42789 25099 42823
rect 25041 42783 25099 42789
rect 25958 42780 25964 42832
rect 26016 42820 26022 42832
rect 28442 42820 28448 42832
rect 26016 42792 28448 42820
rect 26016 42780 26022 42792
rect 28442 42780 28448 42792
rect 28500 42780 28506 42832
rect 28810 42820 28816 42832
rect 28771 42792 28816 42820
rect 28810 42780 28816 42792
rect 28868 42780 28874 42832
rect 29365 42823 29423 42829
rect 29365 42789 29377 42823
rect 29411 42820 29423 42823
rect 29638 42820 29644 42832
rect 29411 42792 29644 42820
rect 29411 42789 29423 42792
rect 29365 42783 29423 42789
rect 29638 42780 29644 42792
rect 29696 42780 29702 42832
rect 30190 42780 30196 42832
rect 30248 42820 30254 42832
rect 30514 42823 30572 42829
rect 30514 42820 30526 42823
rect 30248 42792 30526 42820
rect 30248 42780 30254 42792
rect 30514 42789 30526 42792
rect 30560 42789 30572 42823
rect 34790 42820 34796 42832
rect 34703 42792 34796 42820
rect 30514 42783 30572 42789
rect 34790 42780 34796 42792
rect 34848 42780 34854 42832
rect 34974 42780 34980 42832
rect 35032 42820 35038 42832
rect 35713 42823 35771 42829
rect 35713 42820 35725 42823
rect 35032 42792 35725 42820
rect 35032 42780 35038 42792
rect 35713 42789 35725 42792
rect 35759 42820 35771 42823
rect 36722 42820 36728 42832
rect 35759 42792 36728 42820
rect 35759 42789 35771 42792
rect 35713 42783 35771 42789
rect 36722 42780 36728 42792
rect 36780 42780 36786 42832
rect 39586 42829 39614 42860
rect 40770 42848 40776 42860
rect 40828 42888 40834 42900
rect 41506 42888 41512 42900
rect 40828 42860 41512 42888
rect 40828 42848 40834 42860
rect 41506 42848 41512 42860
rect 41564 42848 41570 42900
rect 39571 42823 39629 42829
rect 39571 42789 39583 42823
rect 39617 42789 39629 42823
rect 39571 42783 39629 42789
rect 40862 42780 40868 42832
rect 40920 42820 40926 42832
rect 41049 42823 41107 42829
rect 41049 42820 41061 42823
rect 40920 42792 41061 42820
rect 40920 42780 40926 42792
rect 41049 42789 41061 42792
rect 41095 42789 41107 42823
rect 41049 42783 41107 42789
rect 41138 42780 41144 42832
rect 41196 42820 41202 42832
rect 41524 42820 41552 42848
rect 41693 42823 41751 42829
rect 41693 42820 41705 42823
rect 41196 42792 41241 42820
rect 41524 42792 41705 42820
rect 41196 42780 41202 42792
rect 41693 42789 41705 42792
rect 41739 42789 41751 42823
rect 43530 42820 43536 42832
rect 43491 42792 43536 42820
rect 41693 42783 41751 42789
rect 43530 42780 43536 42792
rect 43588 42780 43594 42832
rect 20936 42755 20994 42761
rect 20936 42721 20948 42755
rect 20982 42752 20994 42755
rect 21358 42752 21364 42764
rect 20982 42724 21364 42752
rect 20982 42721 20994 42724
rect 20936 42715 20994 42721
rect 21358 42712 21364 42724
rect 21416 42712 21422 42764
rect 23842 42752 23848 42764
rect 23803 42724 23848 42752
rect 23842 42712 23848 42724
rect 23900 42712 23906 42764
rect 25590 42712 25596 42764
rect 25648 42752 25654 42764
rect 27065 42755 27123 42761
rect 25648 42724 25693 42752
rect 25648 42712 25654 42724
rect 27065 42721 27077 42755
rect 27111 42752 27123 42755
rect 27154 42752 27160 42764
rect 27111 42724 27160 42752
rect 27111 42721 27123 42724
rect 27065 42715 27123 42721
rect 27154 42712 27160 42724
rect 27212 42712 27218 42764
rect 27338 42752 27344 42764
rect 27251 42724 27344 42752
rect 27338 42712 27344 42724
rect 27396 42752 27402 42764
rect 28350 42752 28356 42764
rect 27396 42724 28356 42752
rect 27396 42712 27402 42724
rect 28350 42712 28356 42724
rect 28408 42712 28414 42764
rect 35342 42712 35348 42764
rect 35400 42752 35406 42764
rect 36078 42752 36084 42764
rect 35400 42724 36084 42752
rect 35400 42712 35406 42724
rect 36078 42712 36084 42724
rect 36136 42712 36142 42764
rect 36170 42712 36176 42764
rect 36228 42752 36234 42764
rect 37804 42755 37862 42761
rect 36228 42724 36273 42752
rect 36228 42712 36234 42724
rect 37804 42721 37816 42755
rect 37850 42752 37862 42755
rect 38010 42752 38016 42764
rect 37850 42724 38016 42752
rect 37850 42721 37862 42724
rect 37804 42715 37862 42721
rect 38010 42712 38016 42724
rect 38068 42712 38074 42764
rect 38102 42712 38108 42764
rect 38160 42752 38166 42764
rect 38838 42752 38844 42764
rect 38160 42724 38844 42752
rect 38160 42712 38166 42724
rect 38838 42712 38844 42724
rect 38896 42712 38902 42764
rect 16206 42644 16212 42696
rect 16264 42684 16270 42696
rect 16485 42687 16543 42693
rect 16485 42684 16497 42687
rect 16264 42656 16497 42684
rect 16264 42644 16270 42656
rect 16485 42653 16497 42656
rect 16531 42653 16543 42687
rect 16485 42647 16543 42653
rect 18187 42687 18245 42693
rect 18187 42653 18199 42687
rect 18233 42684 18245 42687
rect 19150 42684 19156 42696
rect 18233 42656 19156 42684
rect 18233 42653 18245 42656
rect 18187 42647 18245 42653
rect 19150 42644 19156 42656
rect 19208 42644 19214 42696
rect 24210 42644 24216 42696
rect 24268 42684 24274 42696
rect 24670 42684 24676 42696
rect 24268 42656 24676 42684
rect 24268 42644 24274 42656
rect 24670 42644 24676 42656
rect 24728 42684 24734 42696
rect 24949 42687 25007 42693
rect 24949 42684 24961 42687
rect 24728 42656 24961 42684
rect 24728 42644 24734 42656
rect 24949 42653 24961 42656
rect 24995 42653 25007 42687
rect 25608 42684 25636 42712
rect 28718 42684 28724 42696
rect 25608 42656 28724 42684
rect 24949 42647 25007 42653
rect 28718 42644 28724 42656
rect 28776 42644 28782 42696
rect 30193 42687 30251 42693
rect 30193 42653 30205 42687
rect 30239 42684 30251 42687
rect 30742 42684 30748 42696
rect 30239 42656 30748 42684
rect 30239 42653 30251 42656
rect 30193 42647 30251 42653
rect 30742 42644 30748 42656
rect 30800 42644 30806 42696
rect 32674 42684 32680 42696
rect 32635 42656 32680 42684
rect 32674 42644 32680 42656
rect 32732 42644 32738 42696
rect 34517 42687 34575 42693
rect 34517 42653 34529 42687
rect 34563 42684 34575 42687
rect 34698 42684 34704 42696
rect 34563 42656 34704 42684
rect 34563 42653 34575 42656
rect 34517 42647 34575 42653
rect 34698 42644 34704 42656
rect 34756 42684 34762 42696
rect 36814 42684 36820 42696
rect 34756 42656 36820 42684
rect 34756 42644 34762 42656
rect 36814 42644 36820 42656
rect 36872 42644 36878 42696
rect 38470 42644 38476 42696
rect 38528 42684 38534 42696
rect 39206 42684 39212 42696
rect 38528 42656 39212 42684
rect 38528 42644 38534 42656
rect 39206 42644 39212 42656
rect 39264 42644 39270 42696
rect 42610 42684 42616 42696
rect 41017 42656 42616 42684
rect 17037 42619 17095 42625
rect 17037 42585 17049 42619
rect 17083 42616 17095 42619
rect 17126 42616 17132 42628
rect 17083 42588 17132 42616
rect 17083 42585 17095 42588
rect 17037 42579 17095 42585
rect 17126 42576 17132 42588
rect 17184 42616 17190 42628
rect 19705 42619 19763 42625
rect 19705 42616 19717 42619
rect 17184 42588 19717 42616
rect 17184 42576 17190 42588
rect 19705 42585 19717 42588
rect 19751 42616 19763 42619
rect 22554 42616 22560 42628
rect 19751 42588 22560 42616
rect 19751 42585 19763 42588
rect 19705 42579 19763 42585
rect 22554 42576 22560 42588
rect 22612 42576 22618 42628
rect 27062 42576 27068 42628
rect 27120 42616 27126 42628
rect 28074 42616 28080 42628
rect 27120 42588 28080 42616
rect 27120 42576 27126 42588
rect 28074 42576 28080 42588
rect 28132 42616 28138 42628
rect 32950 42616 32956 42628
rect 28132 42588 32956 42616
rect 28132 42576 28138 42588
rect 32950 42576 32956 42588
rect 33008 42576 33014 42628
rect 36170 42576 36176 42628
rect 36228 42616 36234 42628
rect 40310 42616 40316 42628
rect 36228 42588 40316 42616
rect 36228 42576 36234 42588
rect 40310 42576 40316 42588
rect 40368 42616 40374 42628
rect 41017 42616 41045 42656
rect 42610 42644 42616 42656
rect 42668 42644 42674 42696
rect 43438 42684 43444 42696
rect 43399 42656 43444 42684
rect 43438 42644 43444 42656
rect 43496 42644 43502 42696
rect 43717 42687 43775 42693
rect 43717 42653 43729 42687
rect 43763 42653 43775 42687
rect 43717 42647 43775 42653
rect 40368 42588 41045 42616
rect 40368 42576 40374 42588
rect 41782 42576 41788 42628
rect 41840 42616 41846 42628
rect 43732 42616 43760 42647
rect 41840 42588 43760 42616
rect 41840 42576 41846 42588
rect 15930 42548 15936 42560
rect 15891 42520 15936 42548
rect 15930 42508 15936 42520
rect 15988 42508 15994 42560
rect 21726 42548 21732 42560
rect 21687 42520 21732 42548
rect 21726 42508 21732 42520
rect 21784 42508 21790 42560
rect 28810 42508 28816 42560
rect 28868 42548 28874 42560
rect 29086 42548 29092 42560
rect 28868 42520 29092 42548
rect 28868 42508 28874 42520
rect 29086 42508 29092 42520
rect 29144 42548 29150 42560
rect 31113 42551 31171 42557
rect 31113 42548 31125 42551
rect 29144 42520 31125 42548
rect 29144 42508 29150 42520
rect 31113 42517 31125 42520
rect 31159 42517 31171 42551
rect 31113 42511 31171 42517
rect 36403 42551 36461 42557
rect 36403 42517 36415 42551
rect 36449 42548 36461 42551
rect 36538 42548 36544 42560
rect 36449 42520 36544 42548
rect 36449 42517 36461 42520
rect 36403 42511 36461 42517
rect 36538 42508 36544 42520
rect 36596 42508 36602 42560
rect 38470 42548 38476 42560
rect 38431 42520 38476 42548
rect 38470 42508 38476 42520
rect 38528 42508 38534 42560
rect 40126 42548 40132 42560
rect 40087 42520 40132 42548
rect 40126 42508 40132 42520
rect 40184 42508 40190 42560
rect 42334 42548 42340 42560
rect 42295 42520 42340 42548
rect 42334 42508 42340 42520
rect 42392 42508 42398 42560
rect 1104 42458 48852 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 48852 42458
rect 1104 42384 48852 42406
rect 14691 42347 14749 42353
rect 14691 42313 14703 42347
rect 14737 42344 14749 42347
rect 16206 42344 16212 42356
rect 14737 42316 16212 42344
rect 14737 42313 14749 42316
rect 14691 42307 14749 42313
rect 16206 42304 16212 42316
rect 16264 42304 16270 42356
rect 16298 42304 16304 42356
rect 16356 42344 16362 42356
rect 16485 42347 16543 42353
rect 16485 42344 16497 42347
rect 16356 42316 16497 42344
rect 16356 42304 16362 42316
rect 16485 42313 16497 42316
rect 16531 42344 16543 42347
rect 16666 42344 16672 42356
rect 16531 42316 16672 42344
rect 16531 42313 16543 42316
rect 16485 42307 16543 42313
rect 16666 42304 16672 42316
rect 16724 42344 16730 42356
rect 16761 42347 16819 42353
rect 16761 42344 16773 42347
rect 16724 42316 16773 42344
rect 16724 42304 16730 42316
rect 16761 42313 16773 42316
rect 16807 42313 16819 42347
rect 16761 42307 16819 42313
rect 19150 42304 19156 42356
rect 19208 42344 19214 42356
rect 20717 42347 20775 42353
rect 20717 42344 20729 42347
rect 19208 42316 20729 42344
rect 19208 42304 19214 42316
rect 20717 42313 20729 42316
rect 20763 42313 20775 42347
rect 21358 42344 21364 42356
rect 21319 42316 21364 42344
rect 20717 42307 20775 42313
rect 21358 42304 21364 42316
rect 21416 42304 21422 42356
rect 22922 42344 22928 42356
rect 22883 42316 22928 42344
rect 22922 42304 22928 42316
rect 22980 42304 22986 42356
rect 26513 42347 26571 42353
rect 26513 42313 26525 42347
rect 26559 42344 26571 42347
rect 27338 42344 27344 42356
rect 26559 42316 27344 42344
rect 26559 42313 26571 42316
rect 26513 42307 26571 42313
rect 27338 42304 27344 42316
rect 27396 42304 27402 42356
rect 28307 42347 28365 42353
rect 28307 42313 28319 42347
rect 28353 42344 28365 42347
rect 28626 42344 28632 42356
rect 28353 42316 28632 42344
rect 28353 42313 28365 42316
rect 28307 42307 28365 42313
rect 28626 42304 28632 42316
rect 28684 42304 28690 42356
rect 29086 42344 29092 42356
rect 29047 42316 29092 42344
rect 29086 42304 29092 42316
rect 29144 42304 29150 42356
rect 31941 42347 31999 42353
rect 31941 42313 31953 42347
rect 31987 42344 31999 42347
rect 32214 42344 32220 42356
rect 31987 42316 32220 42344
rect 31987 42313 31999 42316
rect 31941 42307 31999 42313
rect 32214 42304 32220 42316
rect 32272 42304 32278 42356
rect 36170 42304 36176 42356
rect 36228 42344 36234 42356
rect 36265 42347 36323 42353
rect 36265 42344 36277 42347
rect 36228 42316 36277 42344
rect 36228 42304 36234 42316
rect 36265 42313 36277 42316
rect 36311 42313 36323 42347
rect 36265 42307 36323 42313
rect 40126 42304 40132 42356
rect 40184 42344 40190 42356
rect 40221 42347 40279 42353
rect 40221 42344 40233 42347
rect 40184 42316 40233 42344
rect 40184 42304 40190 42316
rect 40221 42313 40233 42316
rect 40267 42313 40279 42347
rect 43441 42347 43499 42353
rect 43441 42344 43453 42347
rect 40221 42307 40279 42313
rect 42766 42316 43453 42344
rect 16224 42276 16252 42304
rect 17129 42279 17187 42285
rect 17129 42276 17141 42279
rect 16224 42248 17141 42276
rect 17129 42245 17141 42248
rect 17175 42245 17187 42279
rect 17129 42239 17187 42245
rect 21039 42279 21097 42285
rect 21039 42245 21051 42279
rect 21085 42276 21097 42279
rect 21726 42276 21732 42288
rect 21085 42248 21732 42276
rect 21085 42245 21097 42248
rect 21039 42239 21097 42245
rect 21726 42236 21732 42248
rect 21784 42236 21790 42288
rect 21818 42236 21824 42288
rect 21876 42276 21882 42288
rect 23293 42279 23351 42285
rect 23293 42276 23305 42279
rect 21876 42248 23305 42276
rect 21876 42236 21882 42248
rect 23293 42245 23305 42248
rect 23339 42245 23351 42279
rect 23293 42239 23351 42245
rect 24946 42236 24952 42288
rect 25004 42276 25010 42288
rect 26053 42279 26111 42285
rect 26053 42276 26065 42279
rect 25004 42248 26065 42276
rect 25004 42236 25010 42248
rect 26053 42245 26065 42248
rect 26099 42276 26111 42279
rect 26329 42279 26387 42285
rect 26329 42276 26341 42279
rect 26099 42248 26341 42276
rect 26099 42245 26111 42248
rect 26053 42239 26111 42245
rect 26329 42245 26341 42248
rect 26375 42245 26387 42279
rect 26329 42239 26387 42245
rect 27154 42236 27160 42288
rect 27212 42276 27218 42288
rect 27617 42279 27675 42285
rect 27617 42276 27629 42279
rect 27212 42248 27629 42276
rect 27212 42236 27218 42248
rect 27617 42245 27629 42248
rect 27663 42245 27675 42279
rect 33502 42276 33508 42288
rect 27617 42239 27675 42245
rect 32048 42248 33508 42276
rect 22002 42208 22008 42220
rect 21963 42180 22008 42208
rect 22002 42168 22008 42180
rect 22060 42168 22066 42220
rect 24167 42211 24225 42217
rect 24167 42177 24179 42211
rect 24213 42208 24225 42211
rect 26697 42211 26755 42217
rect 26697 42208 26709 42211
rect 24213 42180 26709 42208
rect 24213 42177 24225 42180
rect 24167 42171 24225 42177
rect 26697 42177 26709 42180
rect 26743 42208 26755 42211
rect 27985 42211 28043 42217
rect 27985 42208 27997 42211
rect 26743 42180 27997 42208
rect 26743 42177 26755 42180
rect 26697 42171 26755 42177
rect 27985 42177 27997 42180
rect 28031 42177 28043 42211
rect 27985 42171 28043 42177
rect 28350 42168 28356 42220
rect 28408 42208 28414 42220
rect 28408 42180 30880 42208
rect 28408 42168 28414 42180
rect 14620 42143 14678 42149
rect 14620 42109 14632 42143
rect 14666 42140 14678 42143
rect 15562 42140 15568 42152
rect 14666 42112 14964 42140
rect 15523 42112 15568 42140
rect 14666 42109 14678 42112
rect 14620 42103 14678 42109
rect 14936 42016 14964 42112
rect 15562 42100 15568 42112
rect 15620 42100 15626 42152
rect 20162 42100 20168 42152
rect 20220 42140 20226 42152
rect 20968 42143 21026 42149
rect 20968 42140 20980 42143
rect 20220 42112 20980 42140
rect 20220 42100 20226 42112
rect 20968 42109 20980 42112
rect 21014 42140 21026 42143
rect 21542 42140 21548 42152
rect 21014 42112 21548 42140
rect 21014 42109 21026 42112
rect 20968 42103 21026 42109
rect 21542 42100 21548 42112
rect 21600 42140 21606 42152
rect 21729 42143 21787 42149
rect 21729 42140 21741 42143
rect 21600 42112 21741 42140
rect 21600 42100 21606 42112
rect 21729 42109 21741 42112
rect 21775 42109 21787 42143
rect 21729 42103 21787 42109
rect 24080 42143 24138 42149
rect 24080 42109 24092 42143
rect 24126 42140 24138 42143
rect 24126 42112 24624 42140
rect 24126 42109 24138 42112
rect 24080 42103 24138 42109
rect 15473 42075 15531 42081
rect 15473 42041 15485 42075
rect 15519 42072 15531 42075
rect 15927 42075 15985 42081
rect 15927 42072 15939 42075
rect 15519 42044 15939 42072
rect 15519 42041 15531 42044
rect 15473 42035 15531 42041
rect 15927 42041 15939 42044
rect 15973 42072 15985 42075
rect 16206 42072 16212 42084
rect 15973 42044 16212 42072
rect 15973 42041 15985 42044
rect 15927 42035 15985 42041
rect 16206 42032 16212 42044
rect 16264 42032 16270 42084
rect 18325 42075 18383 42081
rect 18325 42041 18337 42075
rect 18371 42072 18383 42075
rect 19153 42075 19211 42081
rect 19153 42072 19165 42075
rect 18371 42044 19165 42072
rect 18371 42041 18383 42044
rect 18325 42035 18383 42041
rect 19153 42041 19165 42044
rect 19199 42072 19211 42075
rect 19429 42075 19487 42081
rect 19429 42072 19441 42075
rect 19199 42044 19441 42072
rect 19199 42041 19211 42044
rect 19153 42035 19211 42041
rect 19429 42041 19441 42044
rect 19475 42041 19487 42075
rect 19429 42035 19487 42041
rect 19521 42075 19579 42081
rect 19521 42041 19533 42075
rect 19567 42041 19579 42075
rect 19521 42035 19579 42041
rect 14918 41964 14924 42016
rect 14976 42004 14982 42016
rect 15013 42007 15071 42013
rect 15013 42004 15025 42007
rect 14976 41976 15025 42004
rect 14976 41964 14982 41976
rect 15013 41973 15025 41976
rect 15059 41973 15071 42007
rect 15013 41967 15071 41973
rect 18877 42007 18935 42013
rect 18877 41973 18889 42007
rect 18923 42004 18935 42007
rect 18966 42004 18972 42016
rect 18923 41976 18972 42004
rect 18923 41973 18935 41976
rect 18877 41967 18935 41973
rect 18966 41964 18972 41976
rect 19024 41964 19030 42016
rect 19334 41964 19340 42016
rect 19392 42004 19398 42016
rect 19536 42004 19564 42035
rect 19886 42032 19892 42084
rect 19944 42072 19950 42084
rect 20073 42075 20131 42081
rect 20073 42072 20085 42075
rect 19944 42044 20085 42072
rect 19944 42032 19950 42044
rect 20073 42041 20085 42044
rect 20119 42072 20131 42075
rect 20119 42044 21864 42072
rect 20119 42041 20131 42044
rect 20073 42035 20131 42041
rect 20349 42007 20407 42013
rect 20349 42004 20361 42007
rect 19392 41976 20361 42004
rect 19392 41964 19398 41976
rect 20349 41973 20361 41976
rect 20395 41973 20407 42007
rect 21836 42004 21864 42044
rect 22094 42032 22100 42084
rect 22152 42072 22158 42084
rect 22646 42072 22652 42084
rect 22152 42044 22197 42072
rect 22607 42044 22652 42072
rect 22152 42032 22158 42044
rect 22646 42032 22652 42044
rect 22704 42032 22710 42084
rect 22664 42004 22692 42032
rect 24596 42016 24624 42112
rect 25774 42100 25780 42152
rect 25832 42140 25838 42152
rect 26510 42140 26516 42152
rect 25832 42112 26516 42140
rect 25832 42100 25838 42112
rect 26510 42100 26516 42112
rect 26568 42100 26574 42152
rect 27614 42100 27620 42152
rect 27672 42100 27678 42152
rect 30852 42149 30880 42180
rect 28236 42143 28294 42149
rect 28236 42109 28248 42143
rect 28282 42140 28294 42143
rect 30561 42143 30619 42149
rect 28282 42112 28764 42140
rect 28282 42109 28294 42112
rect 28236 42103 28294 42109
rect 25130 42072 25136 42084
rect 25091 42044 25136 42072
rect 25130 42032 25136 42044
rect 25188 42032 25194 42084
rect 25225 42075 25283 42081
rect 25225 42041 25237 42075
rect 25271 42041 25283 42075
rect 25225 42035 25283 42041
rect 26329 42075 26387 42081
rect 26329 42041 26341 42075
rect 26375 42072 26387 42075
rect 26789 42075 26847 42081
rect 26789 42072 26801 42075
rect 26375 42044 26801 42072
rect 26375 42041 26387 42044
rect 26329 42035 26387 42041
rect 26789 42041 26801 42044
rect 26835 42072 26847 42075
rect 26970 42072 26976 42084
rect 26835 42044 26976 42072
rect 26835 42041 26847 42044
rect 26789 42035 26847 42041
rect 23842 42004 23848 42016
rect 21836 41976 22692 42004
rect 23803 41976 23848 42004
rect 20349 41967 20407 41973
rect 23842 41964 23848 41976
rect 23900 41964 23906 42016
rect 24578 42004 24584 42016
rect 24539 41976 24584 42004
rect 24578 41964 24584 41976
rect 24636 41964 24642 42016
rect 24949 42007 25007 42013
rect 24949 41973 24961 42007
rect 24995 42004 25007 42007
rect 25038 42004 25044 42016
rect 24995 41976 25044 42004
rect 24995 41973 25007 41976
rect 24949 41967 25007 41973
rect 25038 41964 25044 41976
rect 25096 42004 25102 42016
rect 25240 42004 25268 42035
rect 26970 42032 26976 42044
rect 27028 42032 27034 42084
rect 27341 42075 27399 42081
rect 27341 42041 27353 42075
rect 27387 42072 27399 42075
rect 27632 42072 27660 42100
rect 27890 42072 27896 42084
rect 27387 42044 27896 42072
rect 27387 42041 27399 42044
rect 27341 42035 27399 42041
rect 25958 42004 25964 42016
rect 25096 41976 25964 42004
rect 25096 41964 25102 41976
rect 25958 41964 25964 41976
rect 26016 41964 26022 42016
rect 26510 41964 26516 42016
rect 26568 42004 26574 42016
rect 27356 42004 27384 42035
rect 27890 42032 27896 42044
rect 27948 42032 27954 42084
rect 28736 42013 28764 42112
rect 30561 42109 30573 42143
rect 30607 42109 30619 42143
rect 30561 42103 30619 42109
rect 30837 42143 30895 42149
rect 30837 42109 30849 42143
rect 30883 42140 30895 42143
rect 31202 42140 31208 42152
rect 30883 42112 31208 42140
rect 30883 42109 30895 42112
rect 30837 42103 30895 42109
rect 29825 42075 29883 42081
rect 29825 42041 29837 42075
rect 29871 42072 29883 42075
rect 30576 42072 30604 42103
rect 31202 42100 31208 42112
rect 31260 42100 31266 42152
rect 32048 42149 32076 42248
rect 33502 42236 33508 42248
rect 33560 42276 33566 42288
rect 37918 42276 37924 42288
rect 33560 42248 37924 42276
rect 33560 42236 33566 42248
rect 37918 42236 37924 42248
rect 37976 42236 37982 42288
rect 41877 42279 41935 42285
rect 41877 42245 41889 42279
rect 41923 42276 41935 42279
rect 42766 42276 42794 42316
rect 43441 42313 43453 42316
rect 43487 42344 43499 42347
rect 43530 42344 43536 42356
rect 43487 42316 43536 42344
rect 43487 42313 43499 42316
rect 43441 42307 43499 42313
rect 43530 42304 43536 42316
rect 43588 42304 43594 42356
rect 41923 42248 42794 42276
rect 42889 42279 42947 42285
rect 41923 42245 41935 42248
rect 41877 42239 41935 42245
rect 42889 42245 42901 42279
rect 42935 42276 42947 42279
rect 43070 42276 43076 42288
rect 42935 42248 43076 42276
rect 42935 42245 42947 42248
rect 42889 42239 42947 42245
rect 43070 42236 43076 42248
rect 43128 42276 43134 42288
rect 43714 42276 43720 42288
rect 43128 42248 43720 42276
rect 43128 42236 43134 42248
rect 43714 42236 43720 42248
rect 43772 42236 43778 42288
rect 43806 42236 43812 42288
rect 43864 42276 43870 42288
rect 44174 42276 44180 42288
rect 43864 42248 44180 42276
rect 43864 42236 43870 42248
rect 44174 42236 44180 42248
rect 44232 42276 44238 42288
rect 44453 42279 44511 42285
rect 44453 42276 44465 42279
rect 44232 42248 44465 42276
rect 44232 42236 44238 42248
rect 44453 42245 44465 42248
rect 44499 42245 44511 42279
rect 44453 42239 44511 42245
rect 32674 42208 32680 42220
rect 32635 42180 32680 42208
rect 32674 42168 32680 42180
rect 32732 42208 32738 42220
rect 33413 42211 33471 42217
rect 33413 42208 33425 42211
rect 32732 42180 33425 42208
rect 32732 42168 32738 42180
rect 33413 42177 33425 42180
rect 33459 42177 33471 42211
rect 35618 42208 35624 42220
rect 35579 42180 35624 42208
rect 33413 42171 33471 42177
rect 35618 42168 35624 42180
rect 35676 42168 35682 42220
rect 35989 42211 36047 42217
rect 35989 42177 36001 42211
rect 36035 42208 36047 42211
rect 36538 42208 36544 42220
rect 36035 42180 36544 42208
rect 36035 42177 36047 42180
rect 35989 42171 36047 42177
rect 36538 42168 36544 42180
rect 36596 42168 36602 42220
rect 36814 42208 36820 42220
rect 36775 42180 36820 42208
rect 36814 42168 36820 42180
rect 36872 42168 36878 42220
rect 37829 42211 37887 42217
rect 37829 42177 37841 42211
rect 37875 42208 37887 42211
rect 38010 42208 38016 42220
rect 37875 42180 38016 42208
rect 37875 42177 37887 42180
rect 37829 42171 37887 42177
rect 38010 42168 38016 42180
rect 38068 42208 38074 42220
rect 39482 42208 39488 42220
rect 38068 42180 39488 42208
rect 38068 42168 38074 42180
rect 39482 42168 39488 42180
rect 39540 42168 39546 42220
rect 40770 42208 40776 42220
rect 40731 42180 40776 42208
rect 40770 42168 40776 42180
rect 40828 42168 40834 42220
rect 43438 42168 43444 42220
rect 43496 42208 43502 42220
rect 44821 42211 44879 42217
rect 44821 42208 44833 42211
rect 43496 42180 44833 42208
rect 43496 42168 43502 42180
rect 44821 42177 44833 42180
rect 44867 42177 44879 42211
rect 44821 42171 44879 42177
rect 32033 42143 32091 42149
rect 32033 42140 32045 42143
rect 31588 42112 32045 42140
rect 31588 42072 31616 42112
rect 32033 42109 32045 42112
rect 32079 42109 32091 42143
rect 32033 42103 32091 42109
rect 32214 42100 32220 42152
rect 32272 42140 32278 42152
rect 32493 42143 32551 42149
rect 32493 42140 32505 42143
rect 32272 42112 32505 42140
rect 32272 42100 32278 42112
rect 32493 42109 32505 42112
rect 32539 42109 32551 42143
rect 32493 42103 32551 42109
rect 33648 42143 33706 42149
rect 33648 42109 33660 42143
rect 33694 42140 33706 42143
rect 33694 42112 33870 42140
rect 33694 42109 33706 42112
rect 33648 42103 33706 42109
rect 29871 42044 31616 42072
rect 33842 42072 33870 42112
rect 34054 42100 34060 42152
rect 34112 42140 34118 42152
rect 34609 42143 34667 42149
rect 34609 42140 34621 42143
rect 34112 42112 34621 42140
rect 34112 42100 34118 42112
rect 34609 42109 34621 42112
rect 34655 42109 34667 42143
rect 38194 42140 38200 42152
rect 38107 42112 38200 42140
rect 34609 42103 34667 42109
rect 33842 42044 34192 42072
rect 29871 42041 29883 42044
rect 29825 42035 29883 42041
rect 26568 41976 27384 42004
rect 28721 42007 28779 42013
rect 26568 41964 26574 41976
rect 28721 41973 28733 42007
rect 28767 42004 28779 42007
rect 28810 42004 28816 42016
rect 28767 41976 28816 42004
rect 28767 41973 28779 41976
rect 28721 41967 28779 41973
rect 28810 41964 28816 41976
rect 28868 41964 28874 42016
rect 30190 42004 30196 42016
rect 30151 41976 30196 42004
rect 30190 41964 30196 41976
rect 30248 41964 30254 42016
rect 30561 42007 30619 42013
rect 30561 41973 30573 42007
rect 30607 42004 30619 42007
rect 30742 42004 30748 42016
rect 30607 41976 30748 42004
rect 30607 41973 30619 41976
rect 30561 41967 30619 41973
rect 30742 41964 30748 41976
rect 30800 41964 30806 42016
rect 31588 42013 31616 42044
rect 34164 42016 34192 42044
rect 31573 42007 31631 42013
rect 31573 42004 31585 42007
rect 31531 41976 31585 42004
rect 31573 41973 31585 41976
rect 31619 41973 31631 42007
rect 33042 42004 33048 42016
rect 33003 41976 33048 42004
rect 31573 41967 31631 41973
rect 33042 41964 33048 41976
rect 33100 41964 33106 42016
rect 33735 42007 33793 42013
rect 33735 41973 33747 42007
rect 33781 42004 33793 42007
rect 33962 42004 33968 42016
rect 33781 41976 33968 42004
rect 33781 41973 33793 41976
rect 33735 41967 33793 41973
rect 33962 41964 33968 41976
rect 34020 41964 34026 42016
rect 34146 42004 34152 42016
rect 34107 41976 34152 42004
rect 34146 41964 34152 41976
rect 34204 41964 34210 42016
rect 34624 42004 34652 42103
rect 38194 42100 38200 42112
rect 38252 42140 38258 42152
rect 38657 42143 38715 42149
rect 38657 42140 38669 42143
rect 38252 42112 38669 42140
rect 38252 42100 38258 42112
rect 38657 42109 38669 42112
rect 38703 42109 38715 42143
rect 38657 42103 38715 42109
rect 34974 42072 34980 42084
rect 34935 42044 34980 42072
rect 34974 42032 34980 42044
rect 35032 42032 35038 42084
rect 35069 42075 35127 42081
rect 35069 42041 35081 42075
rect 35115 42041 35127 42075
rect 36630 42072 36636 42084
rect 36591 42044 36636 42072
rect 35069 42035 35127 42041
rect 35084 42004 35112 42035
rect 36630 42032 36636 42044
rect 36688 42032 36694 42084
rect 38286 42032 38292 42084
rect 38344 42072 38350 42084
rect 38565 42075 38623 42081
rect 38565 42072 38577 42075
rect 38344 42044 38577 42072
rect 38344 42032 38350 42044
rect 38565 42041 38577 42044
rect 38611 42072 38623 42075
rect 38978 42075 39036 42081
rect 38978 42072 38990 42075
rect 38611 42044 38990 42072
rect 38611 42041 38623 42044
rect 38565 42035 38623 42041
rect 38978 42041 38990 42044
rect 39024 42072 39036 42075
rect 39024 42044 39988 42072
rect 39024 42041 39036 42044
rect 38978 42035 39036 42041
rect 39960 42016 39988 42044
rect 40126 42032 40132 42084
rect 40184 42072 40190 42084
rect 40865 42075 40923 42081
rect 40865 42072 40877 42075
rect 40184 42044 40877 42072
rect 40184 42032 40190 42044
rect 40865 42041 40877 42044
rect 40911 42041 40923 42075
rect 40865 42035 40923 42041
rect 41417 42075 41475 42081
rect 41417 42041 41429 42075
rect 41463 42072 41475 42075
rect 41966 42072 41972 42084
rect 41463 42044 41972 42072
rect 41463 42041 41475 42044
rect 41417 42035 41475 42041
rect 41966 42032 41972 42044
rect 42024 42032 42030 42084
rect 42334 42072 42340 42084
rect 42295 42044 42340 42072
rect 42334 42032 42340 42044
rect 42392 42032 42398 42084
rect 42429 42075 42487 42081
rect 42429 42041 42441 42075
rect 42475 42041 42487 42075
rect 43898 42072 43904 42084
rect 43859 42044 43904 42072
rect 42429 42035 42487 42041
rect 39574 42004 39580 42016
rect 34624 41976 35112 42004
rect 39535 41976 39580 42004
rect 39574 41964 39580 41976
rect 39632 41964 39638 42016
rect 39942 42004 39948 42016
rect 39903 41976 39948 42004
rect 39942 41964 39948 41976
rect 40000 41964 40006 42016
rect 41322 41964 41328 42016
rect 41380 42004 41386 42016
rect 41693 42007 41751 42013
rect 41693 42004 41705 42007
rect 41380 41976 41705 42004
rect 41380 41964 41386 41976
rect 41693 41973 41705 41976
rect 41739 42004 41751 42007
rect 41877 42007 41935 42013
rect 41877 42004 41889 42007
rect 41739 41976 41889 42004
rect 41739 41973 41751 41976
rect 41693 41967 41751 41973
rect 41877 41973 41889 41976
rect 41923 41973 41935 42007
rect 42058 42004 42064 42016
rect 42019 41976 42064 42004
rect 41877 41967 41935 41973
rect 42058 41964 42064 41976
rect 42116 42004 42122 42016
rect 42444 42004 42472 42035
rect 43898 42032 43904 42044
rect 43956 42032 43962 42084
rect 43990 42032 43996 42084
rect 44048 42072 44054 42084
rect 44048 42044 44093 42072
rect 44048 42032 44054 42044
rect 42116 41976 42472 42004
rect 42116 41964 42122 41976
rect 1104 41914 48852 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 48852 41914
rect 1104 41840 48852 41862
rect 19334 41760 19340 41812
rect 19392 41800 19398 41812
rect 19521 41803 19579 41809
rect 19521 41800 19533 41803
rect 19392 41772 19533 41800
rect 19392 41760 19398 41772
rect 19521 41769 19533 41772
rect 19567 41800 19579 41803
rect 19797 41803 19855 41809
rect 19797 41800 19809 41803
rect 19567 41772 19809 41800
rect 19567 41769 19579 41772
rect 19521 41763 19579 41769
rect 19797 41769 19809 41772
rect 19843 41769 19855 41803
rect 21266 41800 21272 41812
rect 21227 41772 21272 41800
rect 19797 41763 19855 41769
rect 21266 41760 21272 41772
rect 21324 41760 21330 41812
rect 21821 41803 21879 41809
rect 21821 41769 21833 41803
rect 21867 41800 21879 41803
rect 22094 41800 22100 41812
rect 21867 41772 22100 41800
rect 21867 41769 21879 41772
rect 21821 41763 21879 41769
rect 22094 41760 22100 41772
rect 22152 41760 22158 41812
rect 24670 41800 24676 41812
rect 24631 41772 24676 41800
rect 24670 41760 24676 41772
rect 24728 41760 24734 41812
rect 26970 41800 26976 41812
rect 26931 41772 26976 41800
rect 26970 41760 26976 41772
rect 27028 41760 27034 41812
rect 28718 41760 28724 41812
rect 28776 41800 28782 41812
rect 28813 41803 28871 41809
rect 28813 41800 28825 41803
rect 28776 41772 28825 41800
rect 28776 41760 28782 41772
rect 28813 41769 28825 41772
rect 28859 41769 28871 41803
rect 30742 41800 30748 41812
rect 30703 41772 30748 41800
rect 28813 41763 28871 41769
rect 30742 41760 30748 41772
rect 30800 41760 30806 41812
rect 31113 41803 31171 41809
rect 31113 41769 31125 41803
rect 31159 41800 31171 41803
rect 31202 41800 31208 41812
rect 31159 41772 31208 41800
rect 31159 41769 31171 41772
rect 31113 41763 31171 41769
rect 16666 41732 16672 41744
rect 16627 41704 16672 41732
rect 16666 41692 16672 41704
rect 16724 41692 16730 41744
rect 17218 41732 17224 41744
rect 17179 41704 17224 41732
rect 17218 41692 17224 41704
rect 17276 41692 17282 41744
rect 18690 41692 18696 41744
rect 18748 41732 18754 41744
rect 18963 41735 19021 41741
rect 18963 41732 18975 41735
rect 18748 41704 18975 41732
rect 18748 41692 18754 41704
rect 18963 41701 18975 41704
rect 19009 41732 19021 41735
rect 21284 41732 21312 41760
rect 19009 41704 21312 41732
rect 19009 41701 19021 41704
rect 18963 41695 19021 41701
rect 22002 41692 22008 41744
rect 22060 41732 22066 41744
rect 22465 41735 22523 41741
rect 22465 41732 22477 41735
rect 22060 41704 22477 41732
rect 22060 41692 22066 41704
rect 22465 41701 22477 41704
rect 22511 41701 22523 41735
rect 22830 41732 22836 41744
rect 22791 41704 22836 41732
rect 22465 41695 22523 41701
rect 22830 41692 22836 41704
rect 22888 41692 22894 41744
rect 23382 41732 23388 41744
rect 23343 41704 23388 41732
rect 23382 41692 23388 41704
rect 23440 41692 23446 41744
rect 24946 41692 24952 41744
rect 25004 41732 25010 41744
rect 25041 41735 25099 41741
rect 25041 41732 25053 41735
rect 25004 41704 25053 41732
rect 25004 41692 25010 41704
rect 25041 41701 25053 41704
rect 25087 41701 25099 41735
rect 25041 41695 25099 41701
rect 25593 41735 25651 41741
rect 25593 41701 25605 41735
rect 25639 41732 25651 41735
rect 25866 41732 25872 41744
rect 25639 41704 25872 41732
rect 25639 41701 25651 41704
rect 25593 41695 25651 41701
rect 25866 41692 25872 41704
rect 25924 41692 25930 41744
rect 27982 41732 27988 41744
rect 27943 41704 27988 41732
rect 27982 41692 27988 41704
rect 28040 41692 28046 41744
rect 29546 41732 29552 41744
rect 29507 41704 29552 41732
rect 29546 41692 29552 41704
rect 29604 41692 29610 41744
rect 30469 41735 30527 41741
rect 30469 41701 30481 41735
rect 30515 41732 30527 41735
rect 31128 41732 31156 41763
rect 31202 41760 31208 41772
rect 31260 41760 31266 41812
rect 34790 41760 34796 41812
rect 34848 41800 34854 41812
rect 34885 41803 34943 41809
rect 34885 41800 34897 41803
rect 34848 41772 34897 41800
rect 34848 41760 34854 41772
rect 34885 41769 34897 41772
rect 34931 41769 34943 41803
rect 34885 41763 34943 41769
rect 36541 41803 36599 41809
rect 36541 41769 36553 41803
rect 36587 41800 36599 41803
rect 36630 41800 36636 41812
rect 36587 41772 36636 41800
rect 36587 41769 36599 41772
rect 36541 41763 36599 41769
rect 36630 41760 36636 41772
rect 36688 41760 36694 41812
rect 38194 41800 38200 41812
rect 38155 41772 38200 41800
rect 38194 41760 38200 41772
rect 38252 41760 38258 41812
rect 39206 41800 39212 41812
rect 39167 41772 39212 41800
rect 39206 41760 39212 41772
rect 39264 41760 39270 41812
rect 40862 41760 40868 41812
rect 40920 41800 40926 41812
rect 41049 41803 41107 41809
rect 41049 41800 41061 41803
rect 40920 41772 41061 41800
rect 40920 41760 40926 41772
rect 41049 41769 41061 41772
rect 41095 41769 41107 41803
rect 41049 41763 41107 41769
rect 43487 41803 43545 41809
rect 43487 41769 43499 41803
rect 43533 41800 43545 41803
rect 43898 41800 43904 41812
rect 43533 41772 43904 41800
rect 43533 41769 43545 41772
rect 43487 41763 43545 41769
rect 43898 41760 43904 41772
rect 43956 41800 43962 41812
rect 44177 41803 44235 41809
rect 44177 41800 44189 41803
rect 43956 41772 44189 41800
rect 43956 41760 43962 41772
rect 44177 41769 44189 41772
rect 44223 41769 44235 41803
rect 44177 41763 44235 41769
rect 33962 41732 33968 41744
rect 30515 41704 31156 41732
rect 33923 41704 33968 41732
rect 30515 41701 30527 41704
rect 30469 41695 30527 41701
rect 33962 41692 33968 41704
rect 34020 41692 34026 41744
rect 34054 41692 34060 41744
rect 34112 41732 34118 41744
rect 34609 41735 34667 41741
rect 34112 41704 34157 41732
rect 34112 41692 34118 41704
rect 34609 41701 34621 41735
rect 34655 41732 34667 41735
rect 34698 41732 34704 41744
rect 34655 41704 34704 41732
rect 34655 41701 34667 41704
rect 34609 41695 34667 41701
rect 34698 41692 34704 41704
rect 34756 41692 34762 41744
rect 35618 41732 35624 41744
rect 35579 41704 35624 41732
rect 35618 41692 35624 41704
rect 35676 41692 35682 41744
rect 39942 41692 39948 41744
rect 40000 41732 40006 41744
rect 40174 41735 40232 41741
rect 40174 41732 40186 41735
rect 40000 41704 40186 41732
rect 40000 41692 40006 41704
rect 40174 41701 40186 41704
rect 40220 41701 40232 41735
rect 40174 41695 40232 41701
rect 40770 41692 40776 41744
rect 40828 41732 40834 41744
rect 41877 41735 41935 41741
rect 41877 41732 41889 41735
rect 40828 41704 41889 41732
rect 40828 41692 40834 41704
rect 41877 41701 41889 41704
rect 41923 41701 41935 41735
rect 41877 41695 41935 41701
rect 41966 41692 41972 41744
rect 42024 41732 42030 41744
rect 42429 41735 42487 41741
rect 42429 41732 42441 41735
rect 42024 41704 42441 41732
rect 42024 41692 42030 41704
rect 42429 41701 42441 41704
rect 42475 41732 42487 41735
rect 42610 41732 42616 41744
rect 42475 41704 42616 41732
rect 42475 41701 42487 41704
rect 42429 41695 42487 41701
rect 42610 41692 42616 41704
rect 42668 41692 42674 41744
rect 26421 41667 26479 41673
rect 26421 41633 26433 41667
rect 26467 41664 26479 41667
rect 26510 41664 26516 41676
rect 26467 41636 26516 41664
rect 26467 41633 26479 41636
rect 26421 41627 26479 41633
rect 26510 41624 26516 41636
rect 26568 41624 26574 41676
rect 30929 41667 30987 41673
rect 30929 41633 30941 41667
rect 30975 41664 30987 41667
rect 31386 41664 31392 41676
rect 30975 41636 31392 41664
rect 30975 41633 30987 41636
rect 30929 41627 30987 41633
rect 31386 41624 31392 41636
rect 31444 41624 31450 41676
rect 32306 41624 32312 41676
rect 32364 41664 32370 41676
rect 32896 41667 32954 41673
rect 32896 41664 32908 41667
rect 32364 41636 32908 41664
rect 32364 41624 32370 41636
rect 32896 41633 32908 41636
rect 32942 41633 32954 41667
rect 37918 41664 37924 41676
rect 37879 41636 37924 41664
rect 32896 41627 32954 41633
rect 37918 41624 37924 41636
rect 37976 41624 37982 41676
rect 38102 41624 38108 41676
rect 38160 41664 38166 41676
rect 38381 41667 38439 41673
rect 38381 41664 38393 41667
rect 38160 41636 38393 41664
rect 38160 41624 38166 41636
rect 38381 41633 38393 41636
rect 38427 41633 38439 41667
rect 38381 41627 38439 41633
rect 43257 41667 43315 41673
rect 43257 41633 43269 41667
rect 43303 41664 43315 41667
rect 43346 41664 43352 41676
rect 43303 41636 43352 41664
rect 43303 41633 43315 41636
rect 43257 41627 43315 41633
rect 43346 41624 43352 41636
rect 43404 41624 43410 41676
rect 15611 41599 15669 41605
rect 15611 41565 15623 41599
rect 15657 41596 15669 41599
rect 16577 41599 16635 41605
rect 16577 41596 16589 41599
rect 15657 41568 16589 41596
rect 15657 41565 15669 41568
rect 15611 41559 15669 41565
rect 16577 41565 16589 41568
rect 16623 41596 16635 41599
rect 17402 41596 17408 41608
rect 16623 41568 17408 41596
rect 16623 41565 16635 41568
rect 16577 41559 16635 41565
rect 17402 41556 17408 41568
rect 17460 41556 17466 41608
rect 18601 41599 18659 41605
rect 18601 41565 18613 41599
rect 18647 41596 18659 41599
rect 18874 41596 18880 41608
rect 18647 41568 18880 41596
rect 18647 41565 18659 41568
rect 18601 41559 18659 41565
rect 18874 41556 18880 41568
rect 18932 41556 18938 41608
rect 20901 41599 20959 41605
rect 20901 41565 20913 41599
rect 20947 41596 20959 41599
rect 21174 41596 21180 41608
rect 20947 41568 21180 41596
rect 20947 41565 20959 41568
rect 20901 41559 20959 41565
rect 21174 41556 21180 41568
rect 21232 41556 21238 41608
rect 22741 41599 22799 41605
rect 22741 41565 22753 41599
rect 22787 41596 22799 41599
rect 23382 41596 23388 41608
rect 22787 41568 23388 41596
rect 22787 41565 22799 41568
rect 22741 41559 22799 41565
rect 23382 41556 23388 41568
rect 23440 41556 23446 41608
rect 24394 41556 24400 41608
rect 24452 41596 24458 41608
rect 24949 41599 25007 41605
rect 24949 41596 24961 41599
rect 24452 41568 24961 41596
rect 24452 41556 24458 41568
rect 24949 41565 24961 41568
rect 24995 41596 25007 41599
rect 26651 41599 26709 41605
rect 26651 41596 26663 41599
rect 24995 41568 26663 41596
rect 24995 41565 25007 41568
rect 24949 41559 25007 41565
rect 26651 41565 26663 41568
rect 26697 41565 26709 41599
rect 27890 41596 27896 41608
rect 27851 41568 27896 41596
rect 26651 41559 26709 41565
rect 27890 41556 27896 41568
rect 27948 41556 27954 41608
rect 29454 41596 29460 41608
rect 29415 41568 29460 41596
rect 29454 41556 29460 41568
rect 29512 41556 29518 41608
rect 29638 41556 29644 41608
rect 29696 41596 29702 41608
rect 29733 41599 29791 41605
rect 29733 41596 29745 41599
rect 29696 41568 29745 41596
rect 29696 41556 29702 41568
rect 29733 41565 29745 41568
rect 29779 41565 29791 41599
rect 35529 41599 35587 41605
rect 35529 41596 35541 41599
rect 29733 41559 29791 41565
rect 34624 41568 35541 41596
rect 15378 41528 15384 41540
rect 15339 41500 15384 41528
rect 15378 41488 15384 41500
rect 15436 41488 15442 41540
rect 26786 41488 26792 41540
rect 26844 41528 26850 41540
rect 28445 41531 28503 41537
rect 28445 41528 28457 41531
rect 26844 41500 28457 41528
rect 26844 41488 26850 41500
rect 28445 41497 28457 41500
rect 28491 41528 28503 41531
rect 29656 41528 29684 41556
rect 28491 41500 29684 41528
rect 28491 41497 28503 41500
rect 28445 41491 28503 41497
rect 34624 41472 34652 41568
rect 35529 41565 35541 41568
rect 35575 41565 35587 41599
rect 35986 41596 35992 41608
rect 35947 41568 35992 41596
rect 35529 41559 35587 41565
rect 35986 41556 35992 41568
rect 36044 41556 36050 41608
rect 39850 41596 39856 41608
rect 39811 41568 39856 41596
rect 39850 41556 39856 41568
rect 39908 41556 39914 41608
rect 41598 41556 41604 41608
rect 41656 41596 41662 41608
rect 41782 41596 41788 41608
rect 41656 41568 41788 41596
rect 41656 41556 41662 41568
rect 41782 41556 41788 41568
rect 41840 41556 41846 41608
rect 43809 41599 43867 41605
rect 43809 41596 43821 41599
rect 42076 41568 43821 41596
rect 42076 41540 42104 41568
rect 43809 41565 43821 41568
rect 43855 41596 43867 41599
rect 43990 41596 43996 41608
rect 43855 41568 43996 41596
rect 43855 41565 43867 41568
rect 43809 41559 43867 41565
rect 43990 41556 43996 41568
rect 44048 41556 44054 41608
rect 34974 41488 34980 41540
rect 35032 41488 35038 41540
rect 40773 41531 40831 41537
rect 40773 41497 40785 41531
rect 40819 41528 40831 41531
rect 42058 41528 42064 41540
rect 40819 41500 42064 41528
rect 40819 41497 40831 41500
rect 40773 41491 40831 41497
rect 42058 41488 42064 41500
rect 42116 41488 42122 41540
rect 13906 41420 13912 41472
rect 13964 41460 13970 41472
rect 15562 41460 15568 41472
rect 13964 41432 15568 41460
rect 13964 41420 13970 41432
rect 15562 41420 15568 41432
rect 15620 41460 15626 41472
rect 15933 41463 15991 41469
rect 15933 41460 15945 41463
rect 15620 41432 15945 41460
rect 15620 41420 15626 41432
rect 15933 41429 15945 41432
rect 15979 41429 15991 41463
rect 15933 41423 15991 41429
rect 25130 41420 25136 41472
rect 25188 41460 25194 41472
rect 25869 41463 25927 41469
rect 25869 41460 25881 41463
rect 25188 41432 25881 41460
rect 25188 41420 25194 41432
rect 25869 41429 25881 41432
rect 25915 41429 25927 41463
rect 25869 41423 25927 41429
rect 27525 41463 27583 41469
rect 27525 41429 27537 41463
rect 27571 41460 27583 41463
rect 27614 41460 27620 41472
rect 27571 41432 27620 41460
rect 27571 41429 27583 41432
rect 27525 41423 27583 41429
rect 27614 41420 27620 41432
rect 27672 41420 27678 41472
rect 32674 41460 32680 41472
rect 32635 41432 32680 41460
rect 32674 41420 32680 41432
rect 32732 41420 32738 41472
rect 32999 41463 33057 41469
rect 32999 41429 33011 41463
rect 33045 41460 33057 41463
rect 34606 41460 34612 41472
rect 33045 41432 34612 41460
rect 33045 41429 33057 41432
rect 32999 41423 33057 41429
rect 34606 41420 34612 41432
rect 34664 41420 34670 41472
rect 34790 41420 34796 41472
rect 34848 41460 34854 41472
rect 34992 41460 35020 41488
rect 35253 41463 35311 41469
rect 35253 41460 35265 41463
rect 34848 41432 35265 41460
rect 34848 41420 34854 41432
rect 35253 41429 35265 41432
rect 35299 41429 35311 41463
rect 37366 41460 37372 41472
rect 37327 41432 37372 41460
rect 35253 41423 35311 41429
rect 37366 41420 37372 41432
rect 37424 41420 37430 41472
rect 1104 41370 48852 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 48852 41370
rect 1104 41296 48852 41318
rect 16301 41259 16359 41265
rect 16301 41225 16313 41259
rect 16347 41256 16359 41259
rect 16666 41256 16672 41268
rect 16347 41228 16672 41256
rect 16347 41225 16359 41228
rect 16301 41219 16359 41225
rect 16666 41216 16672 41228
rect 16724 41216 16730 41268
rect 17402 41256 17408 41268
rect 17363 41228 17408 41256
rect 17402 41216 17408 41228
rect 17460 41216 17466 41268
rect 18690 41256 18696 41268
rect 18651 41228 18696 41256
rect 18690 41216 18696 41228
rect 18748 41216 18754 41268
rect 21913 41259 21971 41265
rect 21913 41225 21925 41259
rect 21959 41256 21971 41259
rect 22186 41256 22192 41268
rect 21959 41228 22192 41256
rect 21959 41225 21971 41228
rect 21913 41219 21971 41225
rect 22186 41216 22192 41228
rect 22244 41256 22250 41268
rect 22830 41256 22836 41268
rect 22244 41228 22836 41256
rect 22244 41216 22250 41228
rect 22830 41216 22836 41228
rect 22888 41256 22894 41268
rect 23017 41259 23075 41265
rect 23017 41256 23029 41259
rect 22888 41228 23029 41256
rect 22888 41216 22894 41228
rect 23017 41225 23029 41228
rect 23063 41225 23075 41259
rect 23017 41219 23075 41225
rect 23983 41259 24041 41265
rect 23983 41225 23995 41259
rect 24029 41256 24041 41259
rect 25130 41256 25136 41268
rect 24029 41228 25136 41256
rect 24029 41225 24041 41228
rect 23983 41219 24041 41225
rect 25130 41216 25136 41228
rect 25188 41216 25194 41268
rect 25866 41216 25872 41268
rect 25924 41256 25930 41268
rect 25924 41228 27476 41256
rect 25924 41216 25930 41228
rect 20993 41191 21051 41197
rect 20993 41157 21005 41191
rect 21039 41188 21051 41191
rect 21266 41188 21272 41200
rect 21039 41160 21272 41188
rect 21039 41157 21051 41160
rect 20993 41151 21051 41157
rect 21266 41148 21272 41160
rect 21324 41188 21330 41200
rect 21324 41160 23060 41188
rect 21324 41148 21330 41160
rect 23032 41132 23060 41160
rect 24946 41148 24952 41200
rect 25004 41188 25010 41200
rect 25777 41191 25835 41197
rect 25777 41188 25789 41191
rect 25004 41160 25789 41188
rect 25004 41148 25010 41160
rect 25777 41157 25789 41160
rect 25823 41188 25835 41191
rect 26053 41191 26111 41197
rect 26053 41188 26065 41191
rect 25823 41160 26065 41188
rect 25823 41157 25835 41160
rect 25777 41151 25835 41157
rect 26053 41157 26065 41160
rect 26099 41157 26111 41191
rect 26053 41151 26111 41157
rect 16485 41123 16543 41129
rect 16485 41089 16497 41123
rect 16531 41120 16543 41123
rect 17126 41120 17132 41132
rect 16531 41092 17132 41120
rect 16531 41089 16543 41092
rect 16485 41083 16543 41089
rect 17126 41080 17132 41092
rect 17184 41080 17190 41132
rect 19886 41120 19892 41132
rect 19847 41092 19892 41120
rect 19886 41080 19892 41092
rect 19944 41080 19950 41132
rect 22554 41120 22560 41132
rect 22515 41092 22560 41120
rect 22554 41080 22560 41092
rect 22612 41080 22618 41132
rect 23014 41080 23020 41132
rect 23072 41120 23078 41132
rect 24673 41123 24731 41129
rect 24673 41120 24685 41123
rect 23072 41092 24685 41120
rect 23072 41080 23078 41092
rect 24673 41089 24685 41092
rect 24719 41089 24731 41123
rect 24673 41083 24731 41089
rect 23912 41055 23970 41061
rect 23912 41052 23924 41055
rect 23446 41024 23924 41052
rect 15933 40987 15991 40993
rect 15933 40953 15945 40987
rect 15979 40984 15991 40987
rect 16577 40987 16635 40993
rect 15979 40956 16436 40984
rect 15979 40953 15991 40956
rect 15933 40947 15991 40953
rect 16408 40928 16436 40956
rect 16577 40953 16589 40987
rect 16623 40953 16635 40987
rect 16577 40947 16635 40953
rect 17129 40987 17187 40993
rect 17129 40953 17141 40987
rect 17175 40984 17187 40987
rect 17954 40984 17960 40996
rect 17175 40956 17960 40984
rect 17175 40953 17187 40956
rect 17129 40947 17187 40953
rect 13998 40876 14004 40928
rect 14056 40916 14062 40928
rect 15378 40916 15384 40928
rect 14056 40888 15384 40916
rect 14056 40876 14062 40888
rect 15378 40876 15384 40888
rect 15436 40916 15442 40928
rect 15473 40919 15531 40925
rect 15473 40916 15485 40919
rect 15436 40888 15485 40916
rect 15436 40876 15442 40888
rect 15473 40885 15485 40888
rect 15519 40885 15531 40919
rect 16390 40916 16396 40928
rect 16303 40888 16396 40916
rect 15473 40879 15531 40885
rect 16390 40876 16396 40888
rect 16448 40916 16454 40928
rect 16592 40916 16620 40947
rect 17954 40944 17960 40956
rect 18012 40944 18018 40996
rect 19426 40944 19432 40996
rect 19484 40984 19490 40996
rect 19705 40987 19763 40993
rect 19705 40984 19717 40987
rect 19484 40956 19717 40984
rect 19484 40944 19490 40956
rect 19705 40953 19717 40956
rect 19751 40984 19763 40987
rect 19958 40987 20016 40993
rect 19958 40984 19970 40987
rect 19751 40956 19970 40984
rect 19751 40953 19763 40956
rect 19705 40947 19763 40953
rect 19958 40953 19970 40956
rect 20004 40953 20016 40987
rect 20530 40984 20536 40996
rect 20491 40956 20536 40984
rect 19958 40947 20016 40953
rect 20530 40944 20536 40956
rect 20588 40944 20594 40996
rect 21726 40944 21732 40996
rect 21784 40984 21790 40996
rect 22097 40987 22155 40993
rect 22097 40984 22109 40987
rect 21784 40956 22109 40984
rect 21784 40944 21790 40956
rect 22097 40953 22109 40956
rect 22143 40953 22155 40987
rect 22097 40947 22155 40953
rect 22186 40944 22192 40996
rect 22244 40984 22250 40996
rect 22244 40956 22289 40984
rect 22244 40944 22250 40956
rect 22462 40944 22468 40996
rect 22520 40984 22526 40996
rect 23446 40984 23474 41024
rect 23912 41021 23924 41024
rect 23958 41052 23970 41055
rect 24305 41055 24363 41061
rect 24305 41052 24317 41055
rect 23958 41024 24317 41052
rect 23958 41021 23970 41024
rect 23912 41015 23970 41021
rect 24305 41021 24317 41024
rect 24351 41021 24363 41055
rect 24305 41015 24363 41021
rect 22520 40956 23474 40984
rect 24688 40984 24716 41083
rect 24762 41080 24768 41132
rect 24820 41120 24826 41132
rect 24857 41123 24915 41129
rect 24857 41120 24869 41123
rect 24820 41092 24869 41120
rect 24820 41080 24826 41092
rect 24857 41089 24869 41092
rect 24903 41120 24915 41123
rect 26878 41120 26884 41132
rect 24903 41092 26884 41120
rect 24903 41089 24915 41092
rect 24857 41083 24915 41089
rect 26878 41080 26884 41092
rect 26936 41080 26942 41132
rect 27448 41120 27476 41228
rect 27982 41216 27988 41268
rect 28040 41256 28046 41268
rect 28353 41259 28411 41265
rect 28353 41256 28365 41259
rect 28040 41228 28365 41256
rect 28040 41216 28046 41228
rect 28353 41225 28365 41228
rect 28399 41256 28411 41259
rect 28629 41259 28687 41265
rect 28629 41256 28641 41259
rect 28399 41228 28641 41256
rect 28399 41225 28411 41228
rect 28353 41219 28411 41225
rect 28629 41225 28641 41228
rect 28675 41225 28687 41259
rect 29546 41256 29552 41268
rect 29507 41228 29552 41256
rect 28629 41219 28687 41225
rect 29546 41216 29552 41228
rect 29604 41216 29610 41268
rect 33597 41259 33655 41265
rect 33597 41225 33609 41259
rect 33643 41256 33655 41259
rect 33873 41259 33931 41265
rect 33873 41256 33885 41259
rect 33643 41228 33885 41256
rect 33643 41225 33655 41228
rect 33597 41219 33655 41225
rect 33873 41225 33885 41228
rect 33919 41225 33931 41259
rect 33873 41219 33931 41225
rect 28442 41148 28448 41200
rect 28500 41188 28506 41200
rect 31297 41191 31355 41197
rect 31297 41188 31309 41191
rect 28500 41160 31309 41188
rect 28500 41148 28506 41160
rect 31297 41157 31309 41160
rect 31343 41157 31355 41191
rect 33888 41188 33916 41219
rect 33962 41216 33968 41268
rect 34020 41256 34026 41268
rect 34241 41259 34299 41265
rect 34241 41256 34253 41259
rect 34020 41228 34253 41256
rect 34020 41216 34026 41228
rect 34241 41225 34253 41228
rect 34287 41225 34299 41259
rect 34606 41256 34612 41268
rect 34567 41228 34612 41256
rect 34241 41219 34299 41225
rect 34606 41216 34612 41228
rect 34664 41216 34670 41268
rect 37185 41259 37243 41265
rect 37185 41225 37197 41259
rect 37231 41256 37243 41259
rect 38102 41256 38108 41268
rect 37231 41228 38108 41256
rect 37231 41225 37243 41228
rect 37185 41219 37243 41225
rect 38102 41216 38108 41228
rect 38160 41216 38166 41268
rect 39574 41216 39580 41268
rect 39632 41256 39638 41268
rect 40770 41256 40776 41268
rect 39632 41228 40776 41256
rect 39632 41216 39638 41228
rect 40770 41216 40776 41228
rect 40828 41216 40834 41268
rect 41095 41259 41153 41265
rect 41095 41225 41107 41259
rect 41141 41256 41153 41259
rect 42334 41256 42340 41268
rect 41141 41228 42340 41256
rect 41141 41225 41153 41228
rect 41095 41219 41153 41225
rect 42334 41216 42340 41228
rect 42392 41216 42398 41268
rect 43070 41256 43076 41268
rect 42766 41228 43076 41256
rect 34054 41188 34060 41200
rect 33888 41160 34060 41188
rect 31297 41151 31355 41157
rect 34054 41148 34060 41160
rect 34112 41188 34118 41200
rect 35437 41191 35495 41197
rect 35437 41188 35449 41191
rect 34112 41160 35449 41188
rect 34112 41148 34118 41160
rect 35437 41157 35449 41160
rect 35483 41188 35495 41191
rect 35618 41188 35624 41200
rect 35483 41160 35624 41188
rect 35483 41157 35495 41160
rect 35437 41151 35495 41157
rect 35618 41148 35624 41160
rect 35676 41148 35682 41200
rect 36004 41160 37688 41188
rect 36004 41132 36032 41160
rect 28997 41123 29055 41129
rect 28997 41120 29009 41123
rect 27448 41092 29009 41120
rect 28997 41089 29009 41092
rect 29043 41120 29055 41123
rect 29454 41120 29460 41132
rect 29043 41092 29460 41120
rect 29043 41089 29055 41092
rect 28997 41083 29055 41089
rect 29454 41080 29460 41092
rect 29512 41080 29518 41132
rect 32217 41123 32275 41129
rect 32217 41089 32229 41123
rect 32263 41120 32275 41123
rect 32306 41120 32312 41132
rect 32263 41092 32312 41120
rect 32263 41089 32275 41092
rect 32217 41083 32275 41089
rect 32306 41080 32312 41092
rect 32364 41080 32370 41132
rect 32674 41120 32680 41132
rect 32635 41092 32680 41120
rect 32674 41080 32680 41092
rect 32732 41080 32738 41132
rect 35805 41123 35863 41129
rect 35805 41089 35817 41123
rect 35851 41120 35863 41123
rect 35986 41120 35992 41132
rect 35851 41092 35992 41120
rect 35851 41089 35863 41092
rect 35805 41083 35863 41089
rect 35986 41080 35992 41092
rect 36044 41080 36050 41132
rect 36078 41080 36084 41132
rect 36136 41120 36142 41132
rect 37366 41120 37372 41132
rect 36136 41092 36181 41120
rect 37327 41092 37372 41120
rect 36136 41080 36142 41092
rect 37366 41080 37372 41092
rect 37424 41080 37430 41132
rect 37660 41129 37688 41160
rect 37918 41148 37924 41200
rect 37976 41188 37982 41200
rect 38381 41191 38439 41197
rect 38381 41188 38393 41191
rect 37976 41160 38393 41188
rect 37976 41148 37982 41160
rect 38381 41157 38393 41160
rect 38427 41157 38439 41191
rect 42610 41188 42616 41200
rect 42571 41160 42616 41188
rect 38381 41151 38439 41157
rect 42610 41148 42616 41160
rect 42668 41148 42674 41200
rect 37645 41123 37703 41129
rect 37645 41089 37657 41123
rect 37691 41089 37703 41123
rect 37645 41083 37703 41089
rect 38102 41080 38108 41132
rect 38160 41120 38166 41132
rect 38930 41120 38936 41132
rect 38160 41092 38936 41120
rect 38160 41080 38166 41092
rect 38930 41080 38936 41092
rect 38988 41120 38994 41132
rect 39577 41123 39635 41129
rect 38988 41092 39344 41120
rect 38988 41080 38994 41092
rect 27433 41055 27491 41061
rect 27433 41021 27445 41055
rect 27479 41052 27491 41055
rect 27614 41052 27620 41064
rect 27479 41024 27620 41052
rect 27479 41021 27491 41024
rect 27433 41015 27491 41021
rect 27614 41012 27620 41024
rect 27672 41012 27678 41064
rect 29917 41055 29975 41061
rect 29917 41021 29929 41055
rect 29963 41052 29975 41055
rect 30377 41055 30435 41061
rect 30377 41052 30389 41055
rect 29963 41024 30389 41052
rect 29963 41021 29975 41024
rect 29917 41015 29975 41021
rect 30377 41021 30389 41024
rect 30423 41052 30435 41055
rect 30558 41052 30564 41064
rect 30423 41024 30564 41052
rect 30423 41021 30435 41024
rect 30377 41015 30435 41021
rect 30558 41012 30564 41024
rect 30616 41012 30622 41064
rect 39316 41061 39344 41092
rect 39577 41089 39589 41123
rect 39623 41120 39635 41123
rect 39850 41120 39856 41132
rect 39623 41092 39856 41120
rect 39623 41089 39635 41092
rect 39577 41083 39635 41089
rect 39850 41080 39856 41092
rect 39908 41120 39914 41132
rect 40221 41123 40279 41129
rect 40221 41120 40233 41123
rect 39908 41092 40233 41120
rect 39908 41080 39914 41092
rect 40221 41089 40233 41092
rect 40267 41089 40279 41123
rect 40221 41083 40279 41089
rect 42061 41123 42119 41129
rect 42061 41089 42073 41123
rect 42107 41120 42119 41123
rect 42766 41120 42794 41228
rect 43070 41216 43076 41228
rect 43128 41216 43134 41268
rect 43346 41120 43352 41132
rect 42107 41092 42794 41120
rect 43307 41092 43352 41120
rect 42107 41089 42119 41092
rect 42061 41083 42119 41089
rect 43346 41080 43352 41092
rect 43404 41080 43410 41132
rect 38841 41055 38899 41061
rect 38841 41052 38853 41055
rect 38672 41024 38853 41052
rect 25130 40984 25136 40996
rect 24688 40956 25136 40984
rect 22520 40944 22526 40956
rect 25130 40944 25136 40956
rect 25188 40993 25194 40996
rect 25188 40987 25236 40993
rect 25188 40953 25190 40987
rect 25224 40984 25236 40987
rect 27249 40987 27307 40993
rect 27249 40984 27261 40987
rect 25224 40956 27261 40984
rect 25224 40953 25236 40956
rect 25188 40947 25236 40953
rect 27249 40953 27261 40956
rect 27295 40984 27307 40987
rect 27754 40987 27812 40993
rect 27754 40984 27766 40987
rect 27295 40956 27766 40984
rect 27295 40953 27307 40956
rect 27249 40947 27307 40953
rect 27754 40953 27766 40956
rect 27800 40984 27812 40987
rect 28534 40984 28540 40996
rect 27800 40956 28540 40984
rect 27800 40953 27812 40956
rect 27754 40947 27812 40953
rect 25188 40944 25194 40947
rect 28534 40944 28540 40956
rect 28592 40944 28598 40996
rect 30190 40944 30196 40996
rect 30248 40984 30254 40996
rect 33042 40993 33048 40996
rect 30285 40987 30343 40993
rect 30285 40984 30297 40987
rect 30248 40956 30297 40984
rect 30248 40944 30254 40956
rect 30285 40953 30297 40956
rect 30331 40984 30343 40987
rect 30739 40987 30797 40993
rect 30739 40984 30751 40987
rect 30331 40956 30751 40984
rect 30331 40953 30343 40956
rect 30285 40947 30343 40953
rect 30739 40953 30751 40956
rect 30785 40984 30797 40987
rect 32585 40987 32643 40993
rect 32585 40984 32597 40987
rect 30785 40956 32597 40984
rect 30785 40953 30797 40956
rect 30739 40947 30797 40953
rect 32585 40953 32597 40956
rect 32631 40984 32643 40987
rect 33039 40984 33048 40993
rect 32631 40956 33048 40984
rect 32631 40953 32643 40956
rect 32585 40947 32643 40953
rect 33039 40947 33048 40956
rect 33100 40984 33106 40996
rect 33318 40984 33324 40996
rect 33100 40956 33324 40984
rect 33042 40944 33048 40947
rect 33100 40944 33106 40956
rect 33318 40944 33324 40956
rect 33376 40944 33382 40996
rect 35894 40944 35900 40996
rect 35952 40984 35958 40996
rect 35952 40956 35997 40984
rect 35952 40944 35958 40956
rect 36630 40944 36636 40996
rect 36688 40984 36694 40996
rect 37182 40984 37188 40996
rect 36688 40956 37188 40984
rect 36688 40944 36694 40956
rect 37182 40944 37188 40956
rect 37240 40984 37246 40996
rect 37461 40987 37519 40993
rect 37461 40984 37473 40987
rect 37240 40956 37473 40984
rect 37240 40944 37246 40956
rect 37461 40953 37473 40956
rect 37507 40953 37519 40987
rect 37461 40947 37519 40953
rect 16448 40888 16620 40916
rect 16448 40876 16454 40888
rect 18874 40876 18880 40928
rect 18932 40916 18938 40928
rect 18969 40919 19027 40925
rect 18969 40916 18981 40919
rect 18932 40888 18981 40916
rect 18932 40876 18938 40888
rect 18969 40885 18981 40888
rect 19015 40885 19027 40919
rect 18969 40879 19027 40885
rect 21174 40876 21180 40928
rect 21232 40916 21238 40928
rect 21269 40919 21327 40925
rect 21269 40916 21281 40919
rect 21232 40888 21281 40916
rect 21232 40876 21238 40888
rect 21269 40885 21281 40888
rect 21315 40885 21327 40919
rect 23382 40916 23388 40928
rect 23343 40888 23388 40916
rect 21269 40879 21327 40885
rect 23382 40876 23388 40888
rect 23440 40876 23446 40928
rect 26510 40916 26516 40928
rect 26471 40888 26516 40916
rect 26510 40876 26516 40888
rect 26568 40876 26574 40928
rect 31386 40876 31392 40928
rect 31444 40916 31450 40928
rect 31573 40919 31631 40925
rect 31573 40916 31585 40919
rect 31444 40888 31585 40916
rect 31444 40876 31450 40888
rect 31573 40885 31585 40888
rect 31619 40885 31631 40919
rect 35158 40916 35164 40928
rect 35119 40888 35164 40916
rect 31573 40879 31631 40885
rect 35158 40876 35164 40888
rect 35216 40876 35222 40928
rect 38378 40876 38384 40928
rect 38436 40916 38442 40928
rect 38672 40925 38700 41024
rect 38841 41021 38853 41024
rect 38887 41021 38899 41055
rect 38841 41015 38899 41021
rect 39301 41055 39359 41061
rect 39301 41021 39313 41055
rect 39347 41021 39359 41055
rect 39301 41015 39359 41021
rect 39666 41012 39672 41064
rect 39724 41052 39730 41064
rect 40992 41055 41050 41061
rect 40992 41052 41004 41055
rect 39724 41024 41004 41052
rect 39724 41012 39730 41024
rect 40992 41021 41004 41024
rect 41038 41052 41050 41055
rect 41414 41052 41420 41064
rect 41038 41024 41420 41052
rect 41038 41021 41050 41024
rect 40992 41015 41050 41021
rect 41414 41012 41420 41024
rect 41472 41012 41478 41064
rect 42153 40987 42211 40993
rect 42153 40953 42165 40987
rect 42199 40953 42211 40987
rect 42153 40947 42211 40953
rect 38657 40919 38715 40925
rect 38657 40916 38669 40919
rect 38436 40888 38669 40916
rect 38436 40876 38442 40888
rect 38657 40885 38669 40888
rect 38703 40885 38715 40919
rect 38657 40879 38715 40885
rect 39114 40876 39120 40928
rect 39172 40916 39178 40928
rect 39853 40919 39911 40925
rect 39853 40916 39865 40919
rect 39172 40888 39865 40916
rect 39172 40876 39178 40888
rect 39853 40885 39865 40888
rect 39899 40916 39911 40919
rect 39942 40916 39948 40928
rect 39899 40888 39948 40916
rect 39899 40885 39911 40888
rect 39853 40879 39911 40885
rect 39942 40876 39948 40888
rect 40000 40876 40006 40928
rect 41690 40876 41696 40928
rect 41748 40916 41754 40928
rect 41785 40919 41843 40925
rect 41785 40916 41797 40919
rect 41748 40888 41797 40916
rect 41748 40876 41754 40888
rect 41785 40885 41797 40888
rect 41831 40916 41843 40919
rect 42168 40916 42196 40947
rect 41831 40888 42196 40916
rect 41831 40885 41843 40888
rect 41785 40879 41843 40885
rect 1104 40826 48852 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 48852 40826
rect 1104 40752 48852 40774
rect 16390 40712 16396 40724
rect 16351 40684 16396 40712
rect 16390 40672 16396 40684
rect 16448 40672 16454 40724
rect 17126 40712 17132 40724
rect 17087 40684 17132 40712
rect 17126 40672 17132 40684
rect 17184 40672 17190 40724
rect 18138 40672 18144 40724
rect 18196 40712 18202 40724
rect 19058 40712 19064 40724
rect 18196 40684 19064 40712
rect 18196 40672 18202 40684
rect 19058 40672 19064 40684
rect 19116 40672 19122 40724
rect 21315 40715 21373 40721
rect 21315 40681 21327 40715
rect 21361 40712 21373 40715
rect 21726 40712 21732 40724
rect 21361 40684 21732 40712
rect 21361 40681 21373 40684
rect 21315 40675 21373 40681
rect 21726 40672 21732 40684
rect 21784 40672 21790 40724
rect 22097 40715 22155 40721
rect 22097 40681 22109 40715
rect 22143 40712 22155 40715
rect 22186 40712 22192 40724
rect 22143 40684 22192 40712
rect 22143 40681 22155 40684
rect 22097 40675 22155 40681
rect 22186 40672 22192 40684
rect 22244 40712 22250 40724
rect 24394 40712 24400 40724
rect 22244 40684 22416 40712
rect 24355 40684 24400 40712
rect 22244 40672 22250 40684
rect 15835 40647 15893 40653
rect 15835 40613 15847 40647
rect 15881 40644 15893 40647
rect 16206 40644 16212 40656
rect 15881 40616 16212 40644
rect 15881 40613 15893 40616
rect 15835 40607 15893 40613
rect 16206 40604 16212 40616
rect 16264 40604 16270 40656
rect 17402 40644 17408 40656
rect 17363 40616 17408 40644
rect 17402 40604 17408 40616
rect 17460 40604 17466 40656
rect 19886 40644 19892 40656
rect 19847 40616 19892 40644
rect 19886 40604 19892 40616
rect 19944 40604 19950 40656
rect 22388 40653 22416 40684
rect 24394 40672 24400 40684
rect 24452 40672 24458 40724
rect 24762 40712 24768 40724
rect 24723 40684 24768 40712
rect 24762 40672 24768 40684
rect 24820 40672 24826 40724
rect 27890 40712 27896 40724
rect 27851 40684 27896 40712
rect 27890 40672 27896 40684
rect 27948 40672 27954 40724
rect 28534 40672 28540 40724
rect 28592 40712 28598 40724
rect 28629 40715 28687 40721
rect 28629 40712 28641 40715
rect 28592 40684 28641 40712
rect 28592 40672 28598 40684
rect 28629 40681 28641 40684
rect 28675 40681 28687 40715
rect 28629 40675 28687 40681
rect 29181 40715 29239 40721
rect 29181 40681 29193 40715
rect 29227 40712 29239 40715
rect 29546 40712 29552 40724
rect 29227 40684 29552 40712
rect 29227 40681 29239 40684
rect 29181 40675 29239 40681
rect 29546 40672 29552 40684
rect 29604 40672 29610 40724
rect 30558 40712 30564 40724
rect 30519 40684 30564 40712
rect 30558 40672 30564 40684
rect 30616 40672 30622 40724
rect 33827 40715 33885 40721
rect 33827 40681 33839 40715
rect 33873 40712 33885 40715
rect 34790 40712 34796 40724
rect 33873 40684 34796 40712
rect 33873 40681 33885 40684
rect 33827 40675 33885 40681
rect 34790 40672 34796 40684
rect 34848 40672 34854 40724
rect 35158 40672 35164 40724
rect 35216 40712 35222 40724
rect 35621 40715 35679 40721
rect 35621 40712 35633 40715
rect 35216 40684 35633 40712
rect 35216 40672 35222 40684
rect 35621 40681 35633 40684
rect 35667 40712 35679 40715
rect 35894 40712 35900 40724
rect 35667 40684 35900 40712
rect 35667 40681 35679 40684
rect 35621 40675 35679 40681
rect 35894 40672 35900 40684
rect 35952 40672 35958 40724
rect 35986 40672 35992 40724
rect 36044 40712 36050 40724
rect 36587 40715 36645 40721
rect 36044 40684 36089 40712
rect 36044 40672 36050 40684
rect 36587 40681 36599 40715
rect 36633 40712 36645 40715
rect 37366 40712 37372 40724
rect 36633 40684 37372 40712
rect 36633 40681 36645 40684
rect 36587 40675 36645 40681
rect 37366 40672 37372 40684
rect 37424 40672 37430 40724
rect 38930 40712 38936 40724
rect 38891 40684 38936 40712
rect 38930 40672 38936 40684
rect 38988 40672 38994 40724
rect 41598 40712 41604 40724
rect 41559 40684 41604 40712
rect 41598 40672 41604 40684
rect 41656 40672 41662 40724
rect 22373 40647 22431 40653
rect 22373 40613 22385 40647
rect 22419 40613 22431 40647
rect 22373 40607 22431 40613
rect 22646 40604 22652 40656
rect 22704 40644 22710 40656
rect 22925 40647 22983 40653
rect 22925 40644 22937 40647
rect 22704 40616 22937 40644
rect 22704 40604 22710 40616
rect 22925 40613 22937 40616
rect 22971 40613 22983 40647
rect 25038 40644 25044 40656
rect 24999 40616 25044 40644
rect 22925 40607 22983 40613
rect 25038 40604 25044 40616
rect 25096 40604 25102 40656
rect 25593 40647 25651 40653
rect 25593 40613 25605 40647
rect 25639 40644 25651 40647
rect 25866 40644 25872 40656
rect 25639 40616 25872 40644
rect 25639 40613 25651 40616
rect 25593 40607 25651 40613
rect 25866 40604 25872 40616
rect 25924 40604 25930 40656
rect 33318 40604 33324 40656
rect 33376 40644 33382 40656
rect 35022 40647 35080 40653
rect 35022 40644 35034 40647
rect 33376 40616 35034 40644
rect 33376 40604 33382 40616
rect 35022 40613 35034 40616
rect 35068 40644 35080 40647
rect 35250 40644 35256 40656
rect 35068 40616 35256 40644
rect 35068 40613 35080 40616
rect 35022 40607 35080 40613
rect 35250 40604 35256 40616
rect 35308 40604 35314 40656
rect 37182 40604 37188 40656
rect 37240 40644 37246 40656
rect 37277 40647 37335 40653
rect 37277 40644 37289 40647
rect 37240 40616 37289 40644
rect 37240 40604 37246 40616
rect 37277 40613 37289 40616
rect 37323 40613 37335 40647
rect 38948 40644 38976 40672
rect 41874 40644 41880 40656
rect 38948 40616 39620 40644
rect 41835 40616 41880 40644
rect 37277 40607 37335 40613
rect 39592 40588 39620 40616
rect 41874 40604 41880 40616
rect 41932 40604 41938 40656
rect 42426 40644 42432 40656
rect 42339 40616 42432 40644
rect 42426 40604 42432 40616
rect 42484 40644 42490 40656
rect 42610 40644 42616 40656
rect 42484 40616 42616 40644
rect 42484 40604 42490 40616
rect 42610 40604 42616 40616
rect 42668 40604 42674 40656
rect 18598 40536 18604 40588
rect 18656 40576 18662 40588
rect 18969 40579 19027 40585
rect 18969 40576 18981 40579
rect 18656 40548 18981 40576
rect 18656 40536 18662 40548
rect 18969 40545 18981 40548
rect 19015 40545 19027 40579
rect 18969 40539 19027 40545
rect 21244 40579 21302 40585
rect 21244 40545 21256 40579
rect 21290 40576 21302 40579
rect 21542 40576 21548 40588
rect 21290 40548 21548 40576
rect 21290 40545 21302 40548
rect 21244 40539 21302 40545
rect 21542 40536 21548 40548
rect 21600 40536 21606 40588
rect 23804 40579 23862 40585
rect 23804 40545 23816 40579
rect 23850 40576 23862 40579
rect 24302 40576 24308 40588
rect 23850 40548 24308 40576
rect 23850 40545 23862 40548
rect 23804 40539 23862 40545
rect 24302 40536 24308 40548
rect 24360 40536 24366 40588
rect 26970 40576 26976 40588
rect 26931 40548 26976 40576
rect 26970 40536 26976 40548
rect 27028 40536 27034 40588
rect 27249 40579 27307 40585
rect 27249 40545 27261 40579
rect 27295 40576 27307 40579
rect 27338 40576 27344 40588
rect 27295 40548 27344 40576
rect 27295 40545 27307 40548
rect 27249 40539 27307 40545
rect 27338 40536 27344 40548
rect 27396 40536 27402 40588
rect 30558 40576 30564 40588
rect 30519 40548 30564 40576
rect 30558 40536 30564 40548
rect 30616 40536 30622 40588
rect 31021 40579 31079 40585
rect 31021 40545 31033 40579
rect 31067 40576 31079 40579
rect 31386 40576 31392 40588
rect 31067 40548 31392 40576
rect 31067 40545 31079 40548
rect 31021 40539 31079 40545
rect 31386 40536 31392 40548
rect 31444 40536 31450 40588
rect 32125 40579 32183 40585
rect 32125 40545 32137 40579
rect 32171 40545 32183 40579
rect 32125 40539 32183 40545
rect 15286 40468 15292 40520
rect 15344 40508 15350 40520
rect 15473 40511 15531 40517
rect 15473 40508 15485 40511
rect 15344 40480 15485 40508
rect 15344 40468 15350 40480
rect 15473 40477 15485 40480
rect 15519 40477 15531 40511
rect 17310 40508 17316 40520
rect 17271 40480 17316 40508
rect 15473 40471 15531 40477
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 17954 40508 17960 40520
rect 17867 40480 17960 40508
rect 17954 40468 17960 40480
rect 18012 40508 18018 40520
rect 18690 40508 18696 40520
rect 18012 40480 18696 40508
rect 18012 40468 18018 40480
rect 18690 40468 18696 40480
rect 18748 40468 18754 40520
rect 22281 40511 22339 40517
rect 22281 40477 22293 40511
rect 22327 40508 22339 40511
rect 22738 40508 22744 40520
rect 22327 40480 22744 40508
rect 22327 40477 22339 40480
rect 22281 40471 22339 40477
rect 22738 40468 22744 40480
rect 22796 40508 22802 40520
rect 23891 40511 23949 40517
rect 23891 40508 23903 40511
rect 22796 40480 23903 40508
rect 22796 40468 22802 40480
rect 23891 40477 23903 40480
rect 23937 40477 23949 40511
rect 24946 40508 24952 40520
rect 24907 40480 24952 40508
rect 23891 40471 23949 40477
rect 24946 40468 24952 40480
rect 25004 40468 25010 40520
rect 27433 40511 27491 40517
rect 27433 40477 27445 40511
rect 27479 40508 27491 40511
rect 28261 40511 28319 40517
rect 28261 40508 28273 40511
rect 27479 40480 28273 40508
rect 27479 40477 27491 40480
rect 27433 40471 27491 40477
rect 28261 40477 28273 40480
rect 28307 40508 28319 40511
rect 28902 40508 28908 40520
rect 28307 40480 28908 40508
rect 28307 40477 28319 40480
rect 28261 40471 28319 40477
rect 28902 40468 28908 40480
rect 28960 40468 28966 40520
rect 32140 40508 32168 40539
rect 32214 40536 32220 40588
rect 32272 40576 32278 40588
rect 32585 40579 32643 40585
rect 32585 40576 32597 40579
rect 32272 40548 32597 40576
rect 32272 40536 32278 40548
rect 32585 40545 32597 40548
rect 32631 40545 32643 40579
rect 32585 40539 32643 40545
rect 33756 40579 33814 40585
rect 33756 40545 33768 40579
rect 33802 40576 33814 40579
rect 34238 40576 34244 40588
rect 33802 40548 34244 40576
rect 33802 40545 33814 40548
rect 33756 40539 33814 40545
rect 34238 40536 34244 40548
rect 34296 40576 34302 40588
rect 36449 40579 36507 40585
rect 34296 40548 36400 40576
rect 34296 40536 34302 40548
rect 32490 40508 32496 40520
rect 31449 40480 32496 40508
rect 27154 40400 27160 40452
rect 27212 40440 27218 40452
rect 31449 40440 31477 40480
rect 32490 40468 32496 40480
rect 32548 40468 32554 40520
rect 32674 40508 32680 40520
rect 32635 40480 32680 40508
rect 32674 40468 32680 40480
rect 32732 40468 32738 40520
rect 34698 40508 34704 40520
rect 34659 40480 34704 40508
rect 34698 40468 34704 40480
rect 34756 40468 34762 40520
rect 36372 40508 36400 40548
rect 36449 40545 36461 40579
rect 36495 40576 36507 40579
rect 36538 40576 36544 40588
rect 36495 40548 36544 40576
rect 36495 40545 36507 40548
rect 36449 40539 36507 40545
rect 36538 40536 36544 40548
rect 36596 40536 36602 40588
rect 38930 40536 38936 40588
rect 38988 40576 38994 40588
rect 39117 40579 39175 40585
rect 39117 40576 39129 40579
rect 38988 40548 39129 40576
rect 38988 40536 38994 40548
rect 39117 40545 39129 40548
rect 39163 40545 39175 40579
rect 39574 40576 39580 40588
rect 39487 40548 39580 40576
rect 39117 40539 39175 40545
rect 39574 40536 39580 40548
rect 39632 40536 39638 40588
rect 43416 40579 43474 40585
rect 43416 40545 43428 40579
rect 43462 40576 43474 40579
rect 43806 40576 43812 40588
rect 43462 40548 43812 40576
rect 43462 40545 43474 40548
rect 43416 40539 43474 40545
rect 43806 40536 43812 40548
rect 43864 40536 43870 40588
rect 39666 40508 39672 40520
rect 36372 40480 39672 40508
rect 39666 40468 39672 40480
rect 39724 40468 39730 40520
rect 39850 40508 39856 40520
rect 39811 40480 39856 40508
rect 39850 40468 39856 40480
rect 39908 40468 39914 40520
rect 41782 40508 41788 40520
rect 41743 40480 41788 40508
rect 41782 40468 41788 40480
rect 41840 40468 41846 40520
rect 27212 40412 31477 40440
rect 32508 40440 32536 40468
rect 38378 40440 38384 40452
rect 32508 40412 38384 40440
rect 27212 40400 27218 40412
rect 38378 40400 38384 40412
rect 38436 40400 38442 40452
rect 16114 40332 16120 40384
rect 16172 40372 16178 40384
rect 16669 40375 16727 40381
rect 16669 40372 16681 40375
rect 16172 40344 16681 40372
rect 16172 40332 16178 40344
rect 16669 40341 16681 40344
rect 16715 40341 16727 40375
rect 19150 40372 19156 40384
rect 19111 40344 19156 40372
rect 16669 40335 16727 40341
rect 19150 40332 19156 40344
rect 19208 40332 19214 40384
rect 38010 40372 38016 40384
rect 37971 40344 38016 40372
rect 38010 40332 38016 40344
rect 38068 40332 38074 40384
rect 40494 40372 40500 40384
rect 40455 40344 40500 40372
rect 40494 40332 40500 40344
rect 40552 40332 40558 40384
rect 42794 40332 42800 40384
rect 42852 40372 42858 40384
rect 43487 40375 43545 40381
rect 43487 40372 43499 40375
rect 42852 40344 43499 40372
rect 42852 40332 42858 40344
rect 43487 40341 43499 40344
rect 43533 40341 43545 40375
rect 43487 40335 43545 40341
rect 1104 40282 48852 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 48852 40282
rect 1104 40208 48852 40230
rect 17037 40171 17095 40177
rect 17037 40137 17049 40171
rect 17083 40168 17095 40171
rect 17402 40168 17408 40180
rect 17083 40140 17408 40168
rect 17083 40137 17095 40140
rect 17037 40131 17095 40137
rect 17402 40128 17408 40140
rect 17460 40128 17466 40180
rect 18598 40168 18604 40180
rect 18559 40140 18604 40168
rect 18598 40128 18604 40140
rect 18656 40128 18662 40180
rect 19426 40128 19432 40180
rect 19484 40168 19490 40180
rect 19981 40171 20039 40177
rect 19981 40168 19993 40171
rect 19484 40140 19993 40168
rect 19484 40128 19490 40140
rect 19981 40137 19993 40140
rect 20027 40137 20039 40171
rect 19981 40131 20039 40137
rect 21545 40171 21603 40177
rect 21545 40137 21557 40171
rect 21591 40168 21603 40171
rect 22462 40168 22468 40180
rect 21591 40140 22468 40168
rect 21591 40137 21603 40140
rect 21545 40131 21603 40137
rect 17310 40060 17316 40112
rect 17368 40100 17374 40112
rect 17681 40103 17739 40109
rect 17681 40100 17693 40103
rect 17368 40072 17693 40100
rect 17368 40060 17374 40072
rect 17681 40069 17693 40072
rect 17727 40069 17739 40103
rect 21560 40100 21588 40131
rect 22462 40128 22468 40140
rect 22520 40128 22526 40180
rect 22830 40128 22836 40180
rect 22888 40168 22894 40180
rect 23017 40171 23075 40177
rect 23017 40168 23029 40171
rect 22888 40140 23029 40168
rect 22888 40128 22894 40140
rect 23017 40137 23029 40140
rect 23063 40137 23075 40171
rect 23017 40131 23075 40137
rect 25038 40128 25044 40180
rect 25096 40168 25102 40180
rect 25593 40171 25651 40177
rect 25593 40168 25605 40171
rect 25096 40140 25605 40168
rect 25096 40128 25102 40140
rect 25593 40137 25605 40140
rect 25639 40137 25651 40171
rect 25593 40131 25651 40137
rect 26421 40171 26479 40177
rect 26421 40137 26433 40171
rect 26467 40168 26479 40171
rect 27338 40168 27344 40180
rect 26467 40140 27344 40168
rect 26467 40137 26479 40140
rect 26421 40131 26479 40137
rect 27338 40128 27344 40140
rect 27396 40128 27402 40180
rect 28534 40168 28540 40180
rect 28495 40140 28540 40168
rect 28534 40128 28540 40140
rect 28592 40128 28598 40180
rect 28902 40168 28908 40180
rect 28863 40140 28908 40168
rect 28902 40128 28908 40140
rect 28960 40128 28966 40180
rect 32214 40168 32220 40180
rect 32175 40140 32220 40168
rect 32214 40128 32220 40140
rect 32272 40168 32278 40180
rect 32858 40168 32864 40180
rect 32272 40140 32864 40168
rect 32272 40128 32278 40140
rect 32858 40128 32864 40140
rect 32916 40168 32922 40180
rect 33045 40171 33103 40177
rect 33045 40168 33057 40171
rect 32916 40140 33057 40168
rect 32916 40128 32922 40140
rect 33045 40137 33057 40140
rect 33091 40168 33103 40171
rect 34238 40168 34244 40180
rect 33091 40140 33732 40168
rect 34199 40140 34244 40168
rect 33091 40137 33103 40140
rect 33045 40131 33103 40137
rect 17681 40063 17739 40069
rect 21054 40072 21588 40100
rect 16114 39964 16120 39976
rect 16075 39936 16120 39964
rect 16114 39924 16120 39936
rect 16172 39924 16178 39976
rect 19058 39964 19064 39976
rect 19019 39936 19064 39964
rect 19058 39924 19064 39936
rect 19116 39924 19122 39976
rect 20254 39924 20260 39976
rect 20312 39964 20318 39976
rect 21054 39973 21082 40072
rect 22370 40060 22376 40112
rect 22428 40100 22434 40112
rect 22649 40103 22707 40109
rect 22649 40100 22661 40103
rect 22428 40072 22661 40100
rect 22428 40060 22434 40072
rect 22649 40069 22661 40072
rect 22695 40069 22707 40103
rect 22649 40063 22707 40069
rect 23106 40060 23112 40112
rect 23164 40100 23170 40112
rect 23845 40103 23903 40109
rect 23845 40100 23857 40103
rect 23164 40072 23857 40100
rect 23164 40060 23170 40072
rect 23845 40069 23857 40072
rect 23891 40069 23903 40103
rect 26970 40100 26976 40112
rect 26931 40072 26976 40100
rect 23845 40063 23903 40069
rect 26970 40060 26976 40072
rect 27028 40060 27034 40112
rect 21131 40035 21189 40041
rect 21131 40001 21143 40035
rect 21177 40032 21189 40035
rect 22097 40035 22155 40041
rect 22097 40032 22109 40035
rect 21177 40004 22109 40032
rect 21177 40001 21189 40004
rect 21131 39995 21189 40001
rect 22097 40001 22109 40004
rect 22143 40032 22155 40035
rect 23385 40035 23443 40041
rect 23385 40032 23397 40035
rect 22143 40004 23397 40032
rect 22143 40001 22155 40004
rect 22097 39995 22155 40001
rect 23385 40001 23397 40004
rect 23431 40001 23443 40035
rect 27356 40032 27384 40128
rect 32490 40100 32496 40112
rect 32451 40072 32496 40100
rect 32490 40060 32496 40072
rect 32548 40060 32554 40112
rect 27706 40032 27712 40044
rect 27356 40004 27712 40032
rect 23385 39995 23443 40001
rect 27706 39992 27712 40004
rect 27764 40032 27770 40044
rect 27764 40004 28028 40032
rect 27764 39992 27770 40004
rect 21039 39967 21097 39973
rect 21039 39964 21051 39967
rect 20312 39936 21051 39964
rect 20312 39924 20318 39936
rect 21039 39933 21051 39936
rect 21085 39933 21097 39967
rect 21039 39927 21097 39933
rect 23661 39967 23719 39973
rect 23661 39933 23673 39967
rect 23707 39964 23719 39967
rect 23750 39964 23756 39976
rect 23707 39936 23756 39964
rect 23707 39933 23719 39936
rect 23661 39927 23719 39933
rect 23750 39924 23756 39936
rect 23808 39964 23814 39976
rect 24489 39967 24547 39973
rect 24489 39964 24501 39967
rect 23808 39936 24501 39964
rect 23808 39924 23814 39936
rect 24489 39933 24501 39936
rect 24535 39933 24547 39967
rect 24489 39927 24547 39933
rect 24832 39967 24890 39973
rect 24832 39933 24844 39967
rect 24878 39964 24890 39967
rect 25961 39967 26019 39973
rect 24878 39936 25360 39964
rect 24878 39933 24890 39936
rect 24832 39927 24890 39933
rect 15565 39899 15623 39905
rect 15565 39865 15577 39899
rect 15611 39896 15623 39899
rect 16025 39899 16083 39905
rect 16025 39896 16037 39899
rect 15611 39868 16037 39896
rect 15611 39865 15623 39868
rect 15565 39859 15623 39865
rect 16025 39865 16037 39868
rect 16071 39896 16083 39899
rect 16206 39896 16212 39908
rect 16071 39868 16212 39896
rect 16071 39865 16083 39868
rect 16025 39859 16083 39865
rect 16206 39856 16212 39868
rect 16264 39896 16270 39908
rect 16479 39899 16537 39905
rect 16479 39896 16491 39899
rect 16264 39868 16491 39896
rect 16264 39856 16270 39868
rect 16479 39865 16491 39868
rect 16525 39896 16537 39899
rect 18969 39899 19027 39905
rect 18969 39896 18981 39899
rect 16525 39868 18981 39896
rect 16525 39865 16537 39868
rect 16479 39859 16537 39865
rect 18969 39865 18981 39868
rect 19015 39896 19027 39899
rect 19423 39899 19481 39905
rect 19423 39896 19435 39899
rect 19015 39868 19435 39896
rect 19015 39865 19027 39868
rect 18969 39859 19027 39865
rect 19423 39865 19435 39868
rect 19469 39896 19481 39899
rect 20622 39896 20628 39908
rect 19469 39868 20628 39896
rect 19469 39865 19481 39868
rect 19423 39859 19481 39865
rect 20622 39856 20628 39868
rect 20680 39856 20686 39908
rect 22186 39896 22192 39908
rect 22147 39868 22192 39896
rect 22186 39856 22192 39868
rect 22244 39856 22250 39908
rect 24946 39856 24952 39908
rect 25004 39896 25010 39908
rect 25041 39899 25099 39905
rect 25041 39896 25053 39899
rect 25004 39868 25053 39896
rect 25004 39856 25010 39868
rect 25041 39865 25053 39868
rect 25087 39865 25099 39899
rect 25041 39859 25099 39865
rect 15197 39831 15255 39837
rect 15197 39797 15209 39831
rect 15243 39828 15255 39831
rect 15286 39828 15292 39840
rect 15243 39800 15292 39828
rect 15243 39797 15255 39800
rect 15197 39791 15255 39797
rect 15286 39788 15292 39800
rect 15344 39788 15350 39840
rect 21542 39788 21548 39840
rect 21600 39828 21606 39840
rect 21913 39831 21971 39837
rect 21913 39828 21925 39831
rect 21600 39800 21925 39828
rect 21600 39788 21606 39800
rect 21913 39797 21925 39800
rect 21959 39828 21971 39831
rect 22646 39828 22652 39840
rect 21959 39800 22652 39828
rect 21959 39797 21971 39800
rect 21913 39791 21971 39797
rect 22646 39788 22652 39800
rect 22704 39828 22710 39840
rect 23842 39828 23848 39840
rect 22704 39800 23848 39828
rect 22704 39788 22710 39800
rect 23842 39788 23848 39800
rect 23900 39788 23906 39840
rect 24213 39831 24271 39837
rect 24213 39797 24225 39831
rect 24259 39828 24271 39831
rect 24302 39828 24308 39840
rect 24259 39800 24308 39828
rect 24259 39797 24271 39800
rect 24213 39791 24271 39797
rect 24302 39788 24308 39800
rect 24360 39788 24366 39840
rect 25332 39837 25360 39936
rect 25961 39933 25973 39967
rect 26007 39964 26019 39967
rect 26564 39967 26622 39973
rect 26564 39964 26576 39967
rect 26007 39936 26576 39964
rect 26007 39933 26019 39936
rect 25961 39927 26019 39933
rect 26564 39933 26576 39936
rect 26610 39964 26622 39967
rect 26786 39964 26792 39976
rect 26610 39936 26792 39964
rect 26610 39933 26622 39936
rect 26564 39927 26622 39933
rect 26786 39924 26792 39936
rect 26844 39924 26850 39976
rect 28000 39973 28028 40004
rect 27525 39967 27583 39973
rect 27525 39964 27537 39967
rect 27448 39936 27537 39964
rect 26050 39856 26056 39908
rect 26108 39896 26114 39908
rect 26651 39899 26709 39905
rect 26651 39896 26663 39899
rect 26108 39868 26663 39896
rect 26108 39856 26114 39868
rect 26651 39865 26663 39868
rect 26697 39865 26709 39899
rect 26651 39859 26709 39865
rect 27448 39840 27476 39936
rect 27525 39933 27537 39936
rect 27571 39933 27583 39967
rect 27525 39927 27583 39933
rect 27985 39967 28043 39973
rect 27985 39933 27997 39967
rect 28031 39933 28043 39967
rect 30926 39964 30932 39976
rect 30887 39936 30932 39964
rect 27985 39927 28043 39933
rect 30926 39924 30932 39936
rect 30984 39924 30990 39976
rect 31386 39964 31392 39976
rect 31347 39936 31392 39964
rect 31386 39924 31392 39936
rect 31444 39924 31450 39976
rect 33226 39964 33232 39976
rect 33187 39936 33232 39964
rect 33226 39924 33232 39936
rect 33284 39924 33290 39976
rect 33704 39973 33732 40140
rect 34238 40128 34244 40140
rect 34296 40128 34302 40180
rect 35161 40171 35219 40177
rect 35161 40137 35173 40171
rect 35207 40168 35219 40171
rect 35250 40168 35256 40180
rect 35207 40140 35256 40168
rect 35207 40137 35219 40140
rect 35161 40131 35219 40137
rect 35250 40128 35256 40140
rect 35308 40128 35314 40180
rect 35342 40128 35348 40180
rect 35400 40168 35406 40180
rect 37737 40171 37795 40177
rect 37737 40168 37749 40171
rect 35400 40140 37749 40168
rect 35400 40128 35406 40140
rect 37737 40137 37749 40140
rect 37783 40168 37795 40171
rect 37918 40168 37924 40180
rect 37783 40140 37924 40168
rect 37783 40137 37795 40140
rect 37737 40131 37795 40137
rect 37918 40128 37924 40140
rect 37976 40128 37982 40180
rect 39574 40168 39580 40180
rect 39535 40140 39580 40168
rect 39574 40128 39580 40140
rect 39632 40128 39638 40180
rect 41417 40171 41475 40177
rect 41417 40137 41429 40171
rect 41463 40168 41475 40171
rect 41690 40168 41696 40180
rect 41463 40140 41696 40168
rect 41463 40137 41475 40140
rect 41417 40131 41475 40137
rect 41690 40128 41696 40140
rect 41748 40128 41754 40180
rect 41782 40128 41788 40180
rect 41840 40168 41846 40180
rect 42153 40171 42211 40177
rect 42153 40168 42165 40171
rect 41840 40140 42165 40168
rect 41840 40128 41846 40140
rect 42153 40137 42165 40140
rect 42199 40168 42211 40171
rect 44174 40168 44180 40180
rect 42199 40140 44180 40168
rect 42199 40137 42211 40140
rect 42153 40131 42211 40137
rect 44174 40128 44180 40140
rect 44232 40128 44238 40180
rect 36265 40103 36323 40109
rect 36265 40069 36277 40103
rect 36311 40100 36323 40103
rect 36538 40100 36544 40112
rect 36311 40072 36544 40100
rect 36311 40069 36323 40072
rect 36265 40063 36323 40069
rect 36538 40060 36544 40072
rect 36596 40100 36602 40112
rect 42242 40100 42248 40112
rect 36596 40072 42248 40100
rect 36596 40060 36602 40072
rect 42242 40060 42248 40072
rect 42300 40060 42306 40112
rect 33965 40035 34023 40041
rect 33965 40001 33977 40035
rect 34011 40032 34023 40035
rect 34609 40035 34667 40041
rect 34609 40032 34621 40035
rect 34011 40004 34621 40032
rect 34011 40001 34023 40004
rect 33965 39995 34023 40001
rect 34609 40001 34621 40004
rect 34655 40032 34667 40035
rect 34698 40032 34704 40044
rect 34655 40004 34704 40032
rect 34655 40001 34667 40004
rect 34609 39995 34667 40001
rect 34698 39992 34704 40004
rect 34756 39992 34762 40044
rect 35526 39992 35532 40044
rect 35584 40032 35590 40044
rect 36725 40035 36783 40041
rect 36725 40032 36737 40035
rect 35584 40004 36737 40032
rect 35584 39992 35590 40004
rect 36725 40001 36737 40004
rect 36771 40032 36783 40035
rect 36906 40032 36912 40044
rect 36771 40004 36912 40032
rect 36771 40001 36783 40004
rect 36725 39995 36783 40001
rect 36906 39992 36912 40004
rect 36964 39992 36970 40044
rect 38562 40032 38568 40044
rect 38523 40004 38568 40032
rect 38562 39992 38568 40004
rect 38620 39992 38626 40044
rect 39114 39992 39120 40044
rect 39172 40032 39178 40044
rect 40221 40035 40279 40041
rect 40221 40032 40233 40035
rect 39172 40004 40233 40032
rect 39172 39992 39178 40004
rect 40221 40001 40233 40004
rect 40267 40032 40279 40035
rect 41785 40035 41843 40041
rect 40267 40004 40791 40032
rect 40267 40001 40279 40004
rect 40221 39995 40279 40001
rect 33689 39967 33747 39973
rect 33689 39933 33701 39967
rect 33735 39933 33747 39967
rect 33689 39927 33747 39933
rect 35396 39967 35454 39973
rect 35396 39933 35408 39967
rect 35442 39964 35454 39967
rect 35802 39964 35808 39976
rect 35442 39936 35808 39964
rect 35442 39933 35454 39936
rect 35396 39927 35454 39933
rect 35802 39924 35808 39936
rect 35860 39924 35866 39976
rect 37918 39964 37924 39976
rect 37879 39936 37924 39964
rect 37918 39924 37924 39936
rect 37976 39924 37982 39976
rect 38010 39924 38016 39976
rect 38068 39964 38074 39976
rect 38381 39967 38439 39973
rect 38381 39964 38393 39967
rect 38068 39936 38393 39964
rect 38068 39924 38074 39936
rect 38381 39933 38393 39936
rect 38427 39933 38439 39967
rect 38381 39927 38439 39933
rect 39574 39924 39580 39976
rect 39632 39964 39638 39976
rect 40494 39964 40500 39976
rect 39632 39936 40500 39964
rect 39632 39924 39638 39936
rect 40494 39924 40500 39936
rect 40552 39924 40558 39976
rect 40763 39908 40791 40004
rect 41785 40001 41797 40035
rect 41831 40032 41843 40035
rect 41874 40032 41880 40044
rect 41831 40004 41880 40032
rect 41831 40001 41843 40004
rect 41785 39995 41843 40001
rect 41874 39992 41880 40004
rect 41932 39992 41938 40044
rect 42794 39992 42800 40044
rect 42852 40032 42858 40044
rect 43070 40032 43076 40044
rect 42852 40004 42897 40032
rect 43031 40004 43076 40032
rect 42852 39992 42858 40004
rect 43070 39992 43076 40004
rect 43128 39992 43134 40044
rect 35483 39899 35541 39905
rect 35483 39865 35495 39899
rect 35529 39896 35541 39899
rect 36449 39899 36507 39905
rect 36449 39896 36461 39899
rect 35529 39868 36461 39896
rect 35529 39865 35541 39868
rect 35483 39859 35541 39865
rect 36449 39865 36461 39868
rect 36495 39865 36507 39899
rect 36449 39859 36507 39865
rect 36541 39899 36599 39905
rect 36541 39865 36553 39899
rect 36587 39896 36599 39899
rect 36630 39896 36636 39908
rect 36587 39868 36636 39896
rect 36587 39865 36599 39868
rect 36541 39859 36599 39865
rect 25317 39831 25375 39837
rect 25317 39797 25329 39831
rect 25363 39828 25375 39831
rect 25498 39828 25504 39840
rect 25363 39800 25504 39828
rect 25363 39797 25375 39800
rect 25317 39791 25375 39797
rect 25498 39788 25504 39800
rect 25556 39788 25562 39840
rect 27430 39828 27436 39840
rect 27391 39800 27436 39828
rect 27430 39788 27436 39800
rect 27488 39788 27494 39840
rect 27614 39828 27620 39840
rect 27575 39800 27620 39828
rect 27614 39788 27620 39800
rect 27672 39788 27678 39840
rect 30190 39828 30196 39840
rect 30151 39800 30196 39828
rect 30190 39788 30196 39800
rect 30248 39788 30254 39840
rect 30558 39828 30564 39840
rect 30519 39800 30564 39828
rect 30558 39788 30564 39800
rect 30616 39788 30622 39840
rect 30834 39788 30840 39840
rect 30892 39828 30898 39840
rect 30929 39831 30987 39837
rect 30929 39828 30941 39831
rect 30892 39800 30941 39828
rect 30892 39788 30898 39800
rect 30929 39797 30941 39800
rect 30975 39797 30987 39831
rect 36464 39828 36492 39859
rect 36630 39856 36636 39868
rect 36688 39856 36694 39908
rect 40763 39905 40776 39908
rect 40748 39899 40776 39905
rect 40748 39896 40760 39899
rect 40683 39868 40760 39896
rect 40748 39865 40760 39868
rect 40748 39859 40776 39865
rect 40770 39856 40776 39859
rect 40828 39856 40834 39908
rect 42889 39899 42947 39905
rect 42889 39865 42901 39899
rect 42935 39865 42947 39899
rect 42889 39859 42947 39865
rect 36814 39828 36820 39840
rect 36464 39800 36820 39828
rect 30929 39791 30987 39797
rect 36814 39788 36820 39800
rect 36872 39788 36878 39840
rect 38930 39788 38936 39840
rect 38988 39828 38994 39840
rect 39117 39831 39175 39837
rect 39117 39828 39129 39831
rect 38988 39800 39129 39828
rect 38988 39788 38994 39800
rect 39117 39797 39129 39800
rect 39163 39797 39175 39831
rect 39117 39791 39175 39797
rect 41322 39788 41328 39840
rect 41380 39828 41386 39840
rect 42521 39831 42579 39837
rect 42521 39828 42533 39831
rect 41380 39800 42533 39828
rect 41380 39788 41386 39800
rect 42521 39797 42533 39800
rect 42567 39828 42579 39831
rect 42904 39828 42932 39859
rect 43346 39828 43352 39840
rect 42567 39800 43352 39828
rect 42567 39797 42579 39800
rect 42521 39791 42579 39797
rect 43346 39788 43352 39800
rect 43404 39788 43410 39840
rect 43806 39828 43812 39840
rect 43767 39800 43812 39828
rect 43806 39788 43812 39800
rect 43864 39788 43870 39840
rect 1104 39738 48852 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 48852 39738
rect 1104 39664 48852 39686
rect 17129 39627 17187 39633
rect 17129 39593 17141 39627
rect 17175 39624 17187 39627
rect 17954 39624 17960 39636
rect 17175 39596 17960 39624
rect 17175 39593 17187 39596
rect 17129 39587 17187 39593
rect 17954 39584 17960 39596
rect 18012 39624 18018 39636
rect 18012 39596 18184 39624
rect 18012 39584 18018 39596
rect 16206 39516 16212 39568
rect 16264 39556 16270 39568
rect 16530 39559 16588 39565
rect 16530 39556 16542 39559
rect 16264 39528 16542 39556
rect 16264 39516 16270 39528
rect 16530 39525 16542 39528
rect 16576 39525 16588 39559
rect 18046 39556 18052 39568
rect 18007 39528 18052 39556
rect 16530 39519 16588 39525
rect 18046 39516 18052 39528
rect 18104 39516 18110 39568
rect 18156 39565 18184 39596
rect 22186 39584 22192 39636
rect 22244 39624 22250 39636
rect 22373 39627 22431 39633
rect 22373 39624 22385 39627
rect 22244 39596 22385 39624
rect 22244 39584 22250 39596
rect 22373 39593 22385 39596
rect 22419 39593 22431 39627
rect 22738 39624 22744 39636
rect 22699 39596 22744 39624
rect 22373 39587 22431 39593
rect 22738 39584 22744 39596
rect 22796 39584 22802 39636
rect 24946 39624 24952 39636
rect 24907 39596 24952 39624
rect 24946 39584 24952 39596
rect 25004 39584 25010 39636
rect 25958 39584 25964 39636
rect 26016 39624 26022 39636
rect 26697 39627 26755 39633
rect 26697 39624 26709 39627
rect 26016 39596 26709 39624
rect 26016 39584 26022 39596
rect 26697 39593 26709 39596
rect 26743 39593 26755 39627
rect 27706 39624 27712 39636
rect 27667 39596 27712 39624
rect 26697 39587 26755 39593
rect 27706 39584 27712 39596
rect 27764 39584 27770 39636
rect 28534 39584 28540 39636
rect 28592 39624 28598 39636
rect 28629 39627 28687 39633
rect 28629 39624 28641 39627
rect 28592 39596 28641 39624
rect 28592 39584 28598 39596
rect 28629 39593 28641 39596
rect 28675 39593 28687 39627
rect 30926 39624 30932 39636
rect 30887 39596 30932 39624
rect 28629 39587 28687 39593
rect 30926 39584 30932 39596
rect 30984 39584 30990 39636
rect 32214 39624 32220 39636
rect 32175 39596 32220 39624
rect 32214 39584 32220 39596
rect 32272 39584 32278 39636
rect 33226 39624 33232 39636
rect 33187 39596 33232 39624
rect 33226 39584 33232 39596
rect 33284 39624 33290 39636
rect 33410 39624 33416 39636
rect 33284 39596 33416 39624
rect 33284 39584 33290 39596
rect 33410 39584 33416 39596
rect 33468 39624 33474 39636
rect 36541 39627 36599 39633
rect 33468 39596 36492 39624
rect 33468 39584 33474 39596
rect 18141 39559 18199 39565
rect 18141 39525 18153 39559
rect 18187 39525 18199 39559
rect 18690 39556 18696 39568
rect 18603 39528 18696 39556
rect 18141 39519 18199 39525
rect 18690 39516 18696 39528
rect 18748 39556 18754 39568
rect 18748 39528 20576 39556
rect 18748 39516 18754 39528
rect 20548 39500 20576 39528
rect 20622 39516 20628 39568
rect 20680 39556 20686 39568
rect 21815 39559 21873 39565
rect 21815 39556 21827 39559
rect 20680 39528 21827 39556
rect 20680 39516 20686 39528
rect 21815 39525 21827 39528
rect 21861 39556 21873 39559
rect 22002 39556 22008 39568
rect 21861 39528 22008 39556
rect 21861 39525 21873 39528
rect 21815 39519 21873 39525
rect 22002 39516 22008 39528
rect 22060 39516 22066 39568
rect 27154 39556 27160 39568
rect 26896 39528 27160 39556
rect 19521 39491 19579 39497
rect 19521 39457 19533 39491
rect 19567 39488 19579 39491
rect 19610 39488 19616 39500
rect 19567 39460 19616 39488
rect 19567 39457 19579 39460
rect 19521 39451 19579 39457
rect 19610 39448 19616 39460
rect 19668 39448 19674 39500
rect 20530 39448 20536 39500
rect 20588 39488 20594 39500
rect 23201 39491 23259 39497
rect 23201 39488 23213 39491
rect 20588 39460 23213 39488
rect 20588 39448 20594 39460
rect 23201 39457 23213 39460
rect 23247 39488 23259 39491
rect 23290 39488 23296 39500
rect 23247 39460 23296 39488
rect 23247 39457 23259 39460
rect 23201 39451 23259 39457
rect 23290 39448 23296 39460
rect 23348 39448 23354 39500
rect 24118 39448 24124 39500
rect 24176 39488 24182 39500
rect 24213 39491 24271 39497
rect 24213 39488 24225 39491
rect 24176 39460 24225 39488
rect 24176 39448 24182 39460
rect 24213 39457 24225 39460
rect 24259 39457 24271 39491
rect 24213 39451 24271 39457
rect 24578 39448 24584 39500
rect 24636 39488 24642 39500
rect 26896 39497 26924 39528
rect 27154 39516 27160 39528
rect 27212 39516 27218 39568
rect 30190 39516 30196 39568
rect 30248 39556 30254 39568
rect 30561 39559 30619 39565
rect 30561 39556 30573 39559
rect 30248 39528 30573 39556
rect 30248 39516 30254 39528
rect 30561 39525 30573 39528
rect 30607 39556 30619 39559
rect 31386 39556 31392 39568
rect 30607 39528 31392 39556
rect 30607 39525 30619 39528
rect 30561 39519 30619 39525
rect 31386 39516 31392 39528
rect 31444 39516 31450 39568
rect 33318 39516 33324 39568
rect 33376 39556 33382 39568
rect 34010 39559 34068 39565
rect 34010 39556 34022 39559
rect 33376 39528 34022 39556
rect 33376 39516 33382 39528
rect 34010 39525 34022 39528
rect 34056 39525 34068 39559
rect 35621 39559 35679 39565
rect 35621 39556 35633 39559
rect 34010 39519 34068 39525
rect 34624 39528 35633 39556
rect 34624 39500 34652 39528
rect 35621 39525 35633 39528
rect 35667 39525 35679 39559
rect 36464 39556 36492 39596
rect 36541 39593 36553 39627
rect 36587 39624 36599 39627
rect 36630 39624 36636 39636
rect 36587 39596 36636 39624
rect 36587 39593 36599 39596
rect 36541 39587 36599 39593
rect 36630 39584 36636 39596
rect 36688 39584 36694 39636
rect 36814 39624 36820 39636
rect 36775 39596 36820 39624
rect 36814 39584 36820 39596
rect 36872 39584 36878 39636
rect 37921 39627 37979 39633
rect 37921 39593 37933 39627
rect 37967 39624 37979 39627
rect 38102 39624 38108 39636
rect 37967 39596 38108 39624
rect 37967 39593 37979 39596
rect 37921 39587 37979 39593
rect 38102 39584 38108 39596
rect 38160 39584 38166 39636
rect 39114 39624 39120 39636
rect 39075 39596 39120 39624
rect 39114 39584 39120 39596
rect 39172 39584 39178 39636
rect 39669 39627 39727 39633
rect 39669 39593 39681 39627
rect 39715 39624 39727 39627
rect 41322 39624 41328 39636
rect 39715 39596 41328 39624
rect 39715 39593 39727 39596
rect 39669 39587 39727 39593
rect 41322 39584 41328 39596
rect 41380 39584 41386 39636
rect 41417 39627 41475 39633
rect 41417 39593 41429 39627
rect 41463 39624 41475 39627
rect 41874 39624 41880 39636
rect 41463 39596 41880 39624
rect 41463 39593 41475 39596
rect 41417 39587 41475 39593
rect 41874 39584 41880 39596
rect 41932 39584 41938 39636
rect 42794 39584 42800 39636
rect 42852 39624 42858 39636
rect 42852 39596 42897 39624
rect 42852 39584 42858 39596
rect 38654 39556 38660 39568
rect 36464 39528 38660 39556
rect 35621 39519 35679 39525
rect 38654 39516 38660 39528
rect 38712 39556 38718 39568
rect 38930 39556 38936 39568
rect 38712 39528 38936 39556
rect 38712 39516 38718 39528
rect 38930 39516 38936 39528
rect 38988 39516 38994 39568
rect 40770 39556 40776 39568
rect 40731 39528 40776 39556
rect 40770 39516 40776 39528
rect 40828 39516 40834 39568
rect 41782 39556 41788 39568
rect 41695 39528 41788 39556
rect 41782 39516 41788 39528
rect 41840 39556 41846 39568
rect 42426 39556 42432 39568
rect 41840 39528 42432 39556
rect 41840 39516 41846 39528
rect 42426 39516 42432 39528
rect 42484 39516 42490 39568
rect 43438 39516 43444 39568
rect 43496 39556 43502 39568
rect 43533 39559 43591 39565
rect 43533 39556 43545 39559
rect 43496 39528 43545 39556
rect 43496 39516 43502 39528
rect 43533 39525 43545 39528
rect 43579 39525 43591 39559
rect 43533 39519 43591 39525
rect 44085 39559 44143 39565
rect 44085 39525 44097 39559
rect 44131 39556 44143 39559
rect 44174 39556 44180 39568
rect 44131 39528 44180 39556
rect 44131 39525 44143 39528
rect 44085 39519 44143 39525
rect 44174 39516 44180 39528
rect 44232 39516 44238 39568
rect 25292 39491 25350 39497
rect 25292 39488 25304 39491
rect 24636 39460 25304 39488
rect 24636 39448 24642 39460
rect 25292 39457 25304 39460
rect 25338 39488 25350 39491
rect 26881 39491 26939 39497
rect 25338 39460 25820 39488
rect 25338 39457 25350 39460
rect 25292 39451 25350 39457
rect 16209 39423 16267 39429
rect 16209 39389 16221 39423
rect 16255 39420 16267 39423
rect 16758 39420 16764 39432
rect 16255 39392 16764 39420
rect 16255 39389 16267 39392
rect 16209 39383 16267 39389
rect 16758 39380 16764 39392
rect 16816 39380 16822 39432
rect 21450 39420 21456 39432
rect 21411 39392 21456 39420
rect 21450 39380 21456 39392
rect 21508 39380 21514 39432
rect 21358 39312 21364 39364
rect 21416 39352 21422 39364
rect 25792 39361 25820 39460
rect 26881 39457 26893 39491
rect 26927 39457 26939 39491
rect 26881 39451 26939 39457
rect 27065 39491 27123 39497
rect 27065 39457 27077 39491
rect 27111 39488 27123 39491
rect 27246 39488 27252 39500
rect 27111 39460 27252 39488
rect 27111 39457 27123 39460
rect 27065 39451 27123 39457
rect 27246 39448 27252 39460
rect 27304 39448 27310 39500
rect 31018 39488 31024 39500
rect 30979 39460 31024 39488
rect 31018 39448 31024 39460
rect 31076 39448 31082 39500
rect 32030 39448 32036 39500
rect 32088 39488 32094 39500
rect 32125 39491 32183 39497
rect 32125 39488 32137 39491
rect 32088 39460 32137 39488
rect 32088 39448 32094 39460
rect 32125 39457 32137 39460
rect 32171 39457 32183 39491
rect 32125 39451 32183 39457
rect 32585 39491 32643 39497
rect 32585 39457 32597 39491
rect 32631 39457 32643 39491
rect 34606 39488 34612 39500
rect 34519 39460 34612 39488
rect 32585 39451 32643 39457
rect 28258 39420 28264 39432
rect 28219 39392 28264 39420
rect 28258 39380 28264 39392
rect 28316 39380 28322 39432
rect 32306 39420 32312 39432
rect 28552 39392 32312 39420
rect 24397 39355 24455 39361
rect 24397 39352 24409 39355
rect 21416 39324 24409 39352
rect 21416 39312 21422 39324
rect 24397 39321 24409 39324
rect 24443 39321 24455 39355
rect 24397 39315 24455 39321
rect 25777 39355 25835 39361
rect 25777 39321 25789 39355
rect 25823 39352 25835 39355
rect 28552 39352 28580 39392
rect 32306 39380 32312 39392
rect 32364 39380 32370 39432
rect 25823 39324 28580 39352
rect 31205 39355 31263 39361
rect 25823 39321 25835 39324
rect 25777 39315 25835 39321
rect 31205 39321 31217 39355
rect 31251 39352 31263 39355
rect 31846 39352 31852 39364
rect 31251 39324 31852 39352
rect 31251 39321 31263 39324
rect 31205 39315 31263 39321
rect 31846 39312 31852 39324
rect 31904 39352 31910 39364
rect 32600 39352 32628 39451
rect 34606 39448 34612 39460
rect 34664 39448 34670 39500
rect 37737 39491 37795 39497
rect 37737 39457 37749 39491
rect 37783 39488 37795 39491
rect 38010 39488 38016 39500
rect 37783 39460 38016 39488
rect 37783 39457 37795 39460
rect 37737 39451 37795 39457
rect 38010 39448 38016 39460
rect 38068 39448 38074 39500
rect 39850 39448 39856 39500
rect 39908 39488 39914 39500
rect 40218 39488 40224 39500
rect 39908 39460 40224 39488
rect 39908 39448 39914 39460
rect 40218 39448 40224 39460
rect 40276 39488 40282 39500
rect 40497 39491 40555 39497
rect 40497 39488 40509 39491
rect 40276 39460 40509 39488
rect 40276 39448 40282 39460
rect 40497 39457 40509 39460
rect 40543 39457 40555 39491
rect 42242 39488 42248 39500
rect 42203 39460 42248 39488
rect 40497 39451 40555 39457
rect 42242 39448 42248 39460
rect 42300 39448 42306 39500
rect 33686 39420 33692 39432
rect 33647 39392 33692 39420
rect 33686 39380 33692 39392
rect 33744 39380 33750 39432
rect 35526 39420 35532 39432
rect 35487 39392 35532 39420
rect 35526 39380 35532 39392
rect 35584 39380 35590 39432
rect 38746 39420 38752 39432
rect 38707 39392 38752 39420
rect 38746 39380 38752 39392
rect 38804 39380 38810 39432
rect 42383 39423 42441 39429
rect 42383 39389 42395 39423
rect 42429 39420 42441 39423
rect 42702 39420 42708 39432
rect 42429 39392 42708 39420
rect 42429 39389 42441 39392
rect 42383 39383 42441 39389
rect 42702 39380 42708 39392
rect 42760 39420 42766 39432
rect 43441 39423 43499 39429
rect 43441 39420 43453 39423
rect 42760 39392 43453 39420
rect 42760 39380 42766 39392
rect 43441 39389 43453 39392
rect 43487 39389 43499 39423
rect 43441 39383 43499 39389
rect 36078 39352 36084 39364
rect 31904 39324 32628 39352
rect 36039 39324 36084 39352
rect 31904 39312 31910 39324
rect 36078 39312 36084 39324
rect 36136 39312 36142 39364
rect 19058 39284 19064 39296
rect 19019 39256 19064 39284
rect 19058 39244 19064 39256
rect 19116 39244 19122 39296
rect 19426 39244 19432 39296
rect 19484 39284 19490 39296
rect 19659 39287 19717 39293
rect 19659 39284 19671 39287
rect 19484 39256 19671 39284
rect 19484 39244 19490 39256
rect 19659 39253 19671 39256
rect 19705 39253 19717 39287
rect 19659 39247 19717 39253
rect 21082 39244 21088 39296
rect 21140 39284 21146 39296
rect 23339 39287 23397 39293
rect 23339 39284 23351 39287
rect 21140 39256 23351 39284
rect 21140 39244 21146 39256
rect 23339 39253 23351 39256
rect 23385 39253 23397 39287
rect 23339 39247 23397 39253
rect 24946 39244 24952 39296
rect 25004 39284 25010 39296
rect 25363 39287 25421 39293
rect 25363 39284 25375 39287
rect 25004 39256 25375 39284
rect 25004 39244 25010 39256
rect 25363 39253 25375 39256
rect 25409 39253 25421 39287
rect 25363 39247 25421 39253
rect 25498 39244 25504 39296
rect 25556 39284 25562 39296
rect 28626 39284 28632 39296
rect 25556 39256 28632 39284
rect 25556 39244 25562 39256
rect 28626 39244 28632 39256
rect 28684 39244 28690 39296
rect 29178 39284 29184 39296
rect 29139 39256 29184 39284
rect 29178 39244 29184 39256
rect 29236 39244 29242 39296
rect 29454 39284 29460 39296
rect 29415 39256 29460 39284
rect 29454 39244 29460 39256
rect 29512 39244 29518 39296
rect 30926 39244 30932 39296
rect 30984 39284 30990 39296
rect 35342 39284 35348 39296
rect 30984 39256 35348 39284
rect 30984 39244 30990 39256
rect 35342 39244 35348 39256
rect 35400 39244 35406 39296
rect 1104 39194 48852 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 48852 39194
rect 1104 39120 48852 39142
rect 16206 39080 16212 39092
rect 16167 39052 16212 39080
rect 16206 39040 16212 39052
rect 16264 39040 16270 39092
rect 17497 39083 17555 39089
rect 17497 39049 17509 39083
rect 17543 39080 17555 39083
rect 18046 39080 18052 39092
rect 17543 39052 18052 39080
rect 17543 39049 17555 39052
rect 17497 39043 17555 39049
rect 18046 39040 18052 39052
rect 18104 39040 18110 39092
rect 18598 39040 18604 39092
rect 18656 39080 18662 39092
rect 20349 39083 20407 39089
rect 20349 39080 20361 39083
rect 18656 39052 20361 39080
rect 18656 39040 18662 39052
rect 20349 39049 20361 39052
rect 20395 39049 20407 39083
rect 20349 39043 20407 39049
rect 22603 39083 22661 39089
rect 22603 39049 22615 39083
rect 22649 39080 22661 39083
rect 23382 39080 23388 39092
rect 22649 39052 23388 39080
rect 22649 39049 22661 39052
rect 22603 39043 22661 39049
rect 13906 38944 13912 38956
rect 13867 38916 13912 38944
rect 13906 38904 13912 38916
rect 13964 38904 13970 38956
rect 15286 38944 15292 38956
rect 15247 38916 15292 38944
rect 15286 38904 15292 38916
rect 15344 38904 15350 38956
rect 19058 38944 19064 38956
rect 15672 38916 16528 38944
rect 19019 38916 19064 38944
rect 13081 38879 13139 38885
rect 13081 38845 13093 38879
rect 13127 38876 13139 38879
rect 13449 38879 13507 38885
rect 13449 38876 13461 38879
rect 13127 38848 13461 38876
rect 13127 38845 13139 38848
rect 13081 38839 13139 38845
rect 13449 38845 13461 38848
rect 13495 38876 13507 38879
rect 13630 38876 13636 38888
rect 13495 38848 13636 38876
rect 13495 38845 13507 38848
rect 13449 38839 13507 38845
rect 13630 38836 13636 38848
rect 13688 38836 13694 38888
rect 13725 38879 13783 38885
rect 13725 38845 13737 38879
rect 13771 38876 13783 38879
rect 13814 38876 13820 38888
rect 13771 38848 13820 38876
rect 13771 38845 13783 38848
rect 13725 38839 13783 38845
rect 13814 38836 13820 38848
rect 13872 38836 13878 38888
rect 14645 38879 14703 38885
rect 14645 38845 14657 38879
rect 14691 38876 14703 38879
rect 14737 38879 14795 38885
rect 14737 38876 14749 38879
rect 14691 38848 14749 38876
rect 14691 38845 14703 38848
rect 14645 38839 14703 38845
rect 14737 38845 14749 38848
rect 14783 38845 14795 38879
rect 14737 38839 14795 38845
rect 15197 38879 15255 38885
rect 15197 38845 15209 38879
rect 15243 38876 15255 38879
rect 15672 38876 15700 38916
rect 16500 38888 16528 38916
rect 19058 38904 19064 38916
rect 19116 38904 19122 38956
rect 20364 38944 20392 39043
rect 23382 39040 23388 39052
rect 23440 39040 23446 39092
rect 26697 39083 26755 39089
rect 26697 39049 26709 39083
rect 26743 39080 26755 39083
rect 27154 39080 27160 39092
rect 26743 39052 27160 39080
rect 26743 39049 26755 39052
rect 26697 39043 26755 39049
rect 27154 39040 27160 39052
rect 27212 39040 27218 39092
rect 28534 39040 28540 39092
rect 28592 39080 28598 39092
rect 28629 39083 28687 39089
rect 28629 39080 28641 39083
rect 28592 39052 28641 39080
rect 28592 39040 28598 39052
rect 28629 39049 28641 39052
rect 28675 39080 28687 39083
rect 28718 39080 28724 39092
rect 28675 39052 28724 39080
rect 28675 39049 28687 39052
rect 28629 39043 28687 39049
rect 28718 39040 28724 39052
rect 28776 39040 28782 39092
rect 29089 39083 29147 39089
rect 29089 39049 29101 39083
rect 29135 39080 29147 39083
rect 29178 39080 29184 39092
rect 29135 39052 29184 39080
rect 29135 39049 29147 39052
rect 29089 39043 29147 39049
rect 29178 39040 29184 39052
rect 29236 39040 29242 39092
rect 30377 39083 30435 39089
rect 30377 39049 30389 39083
rect 30423 39080 30435 39083
rect 31018 39080 31024 39092
rect 30423 39052 31024 39080
rect 30423 39049 30435 39052
rect 30377 39043 30435 39049
rect 31018 39040 31024 39052
rect 31076 39040 31082 39092
rect 32030 39040 32036 39092
rect 32088 39080 32094 39092
rect 32125 39083 32183 39089
rect 32125 39080 32137 39083
rect 32088 39052 32137 39080
rect 32088 39040 32094 39052
rect 32125 39049 32137 39052
rect 32171 39049 32183 39083
rect 32858 39080 32864 39092
rect 32819 39052 32864 39080
rect 32125 39043 32183 39049
rect 32858 39040 32864 39052
rect 32916 39080 32922 39092
rect 34606 39080 34612 39092
rect 32916 39052 33548 39080
rect 34567 39052 34612 39080
rect 32916 39040 32922 39052
rect 22002 39012 22008 39024
rect 21915 38984 22008 39012
rect 22002 38972 22008 38984
rect 22060 39012 22066 39024
rect 23290 39012 23296 39024
rect 22060 38984 23060 39012
rect 23251 38984 23296 39012
rect 22060 38972 22066 38984
rect 23032 38956 23060 38984
rect 23290 38972 23296 38984
rect 23348 38972 23354 39024
rect 25130 39012 25136 39024
rect 25091 38984 25136 39012
rect 25130 38972 25136 38984
rect 25188 38972 25194 39024
rect 27062 38972 27068 39024
rect 27120 39012 27126 39024
rect 32493 39015 32551 39021
rect 32493 39012 32505 39015
rect 27120 38984 32505 39012
rect 27120 38972 27126 38984
rect 32493 38981 32505 38984
rect 32539 39012 32551 39015
rect 32539 38984 33088 39012
rect 32539 38981 32551 38984
rect 32493 38975 32551 38981
rect 20364 38916 21404 38944
rect 21376 38888 21404 38916
rect 21450 38904 21456 38956
rect 21508 38944 21514 38956
rect 21637 38947 21695 38953
rect 21637 38944 21649 38947
rect 21508 38916 21649 38944
rect 21508 38904 21514 38916
rect 21637 38913 21649 38916
rect 21683 38944 21695 38947
rect 22281 38947 22339 38953
rect 22281 38944 22293 38947
rect 21683 38916 22293 38944
rect 21683 38913 21695 38916
rect 21637 38907 21695 38913
rect 22281 38913 22293 38916
rect 22327 38913 22339 38947
rect 22281 38907 22339 38913
rect 23014 38904 23020 38956
rect 23072 38904 23078 38956
rect 25498 38944 25504 38956
rect 23354 38916 25504 38944
rect 16301 38879 16359 38885
rect 16301 38876 16313 38879
rect 15243 38848 15700 38876
rect 15764 38848 16313 38876
rect 15243 38845 15255 38848
rect 15197 38839 15255 38845
rect 13538 38700 13544 38752
rect 13596 38740 13602 38752
rect 14660 38740 14688 38839
rect 15764 38752 15792 38848
rect 16301 38845 16313 38848
rect 16347 38845 16359 38879
rect 16301 38839 16359 38845
rect 16482 38836 16488 38888
rect 16540 38876 16546 38888
rect 16853 38879 16911 38885
rect 16853 38876 16865 38879
rect 16540 38848 16865 38876
rect 16540 38836 16546 38848
rect 16853 38845 16865 38848
rect 16899 38876 16911 38879
rect 18325 38879 18383 38885
rect 16899 38848 17908 38876
rect 16899 38845 16911 38848
rect 16853 38839 16911 38845
rect 17880 38817 17908 38848
rect 18325 38845 18337 38879
rect 18371 38876 18383 38879
rect 18417 38879 18475 38885
rect 18417 38876 18429 38879
rect 18371 38848 18429 38876
rect 18371 38845 18383 38848
rect 18325 38839 18383 38845
rect 18417 38845 18429 38848
rect 18463 38876 18475 38879
rect 18782 38876 18788 38888
rect 18463 38848 18788 38876
rect 18463 38845 18475 38848
rect 18417 38839 18475 38845
rect 18782 38836 18788 38848
rect 18840 38836 18846 38888
rect 18969 38879 19027 38885
rect 18969 38845 18981 38879
rect 19015 38876 19027 38879
rect 19150 38876 19156 38888
rect 19015 38848 19156 38876
rect 19015 38845 19027 38848
rect 18969 38839 19027 38845
rect 17865 38811 17923 38817
rect 17865 38777 17877 38811
rect 17911 38808 17923 38811
rect 18046 38808 18052 38820
rect 17911 38780 18052 38808
rect 17911 38777 17923 38780
rect 17865 38771 17923 38777
rect 18046 38768 18052 38780
rect 18104 38808 18110 38820
rect 18984 38808 19012 38839
rect 19150 38836 19156 38848
rect 19208 38836 19214 38888
rect 19610 38876 19616 38888
rect 19523 38848 19616 38876
rect 19610 38836 19616 38848
rect 19668 38876 19674 38888
rect 21177 38879 21235 38885
rect 19668 38848 20392 38876
rect 19668 38836 19674 38848
rect 18104 38780 19012 38808
rect 18104 38768 18110 38780
rect 20364 38752 20392 38848
rect 21177 38845 21189 38879
rect 21223 38845 21235 38879
rect 21177 38839 21235 38845
rect 20809 38811 20867 38817
rect 20809 38777 20821 38811
rect 20855 38808 20867 38811
rect 21192 38808 21220 38839
rect 21358 38836 21364 38888
rect 21416 38876 21422 38888
rect 22532 38879 22590 38885
rect 22532 38876 22544 38879
rect 21416 38848 21509 38876
rect 22112 38848 22544 38876
rect 21416 38836 21422 38848
rect 22002 38808 22008 38820
rect 20855 38780 22008 38808
rect 20855 38777 20867 38780
rect 20809 38771 20867 38777
rect 22002 38768 22008 38780
rect 22060 38768 22066 38820
rect 15746 38740 15752 38752
rect 13596 38712 14688 38740
rect 15707 38712 15752 38740
rect 13596 38700 13602 38712
rect 15746 38700 15752 38712
rect 15804 38700 15810 38752
rect 16577 38743 16635 38749
rect 16577 38709 16589 38743
rect 16623 38740 16635 38743
rect 16758 38740 16764 38752
rect 16623 38712 16764 38740
rect 16623 38709 16635 38712
rect 16577 38703 16635 38709
rect 16758 38700 16764 38712
rect 16816 38700 16822 38752
rect 20346 38700 20352 38752
rect 20404 38740 20410 38752
rect 22112 38740 22140 38848
rect 22532 38845 22544 38848
rect 22578 38876 22590 38879
rect 22925 38879 22983 38885
rect 22925 38876 22937 38879
rect 22578 38848 22937 38876
rect 22578 38845 22590 38848
rect 22532 38839 22590 38845
rect 22925 38845 22937 38848
rect 22971 38876 22983 38879
rect 23354 38876 23382 38916
rect 25498 38904 25504 38916
rect 25556 38904 25562 38956
rect 28350 38904 28356 38956
rect 28408 38944 28414 38956
rect 29365 38947 29423 38953
rect 29365 38944 29377 38947
rect 28408 38916 29377 38944
rect 28408 38904 28414 38916
rect 29365 38913 29377 38916
rect 29411 38944 29423 38947
rect 29454 38944 29460 38956
rect 29411 38916 29460 38944
rect 29411 38913 29423 38916
rect 29365 38907 29423 38913
rect 29454 38904 29460 38916
rect 29512 38904 29518 38956
rect 29638 38944 29644 38956
rect 29599 38916 29644 38944
rect 29638 38904 29644 38916
rect 29696 38904 29702 38956
rect 22971 38848 23382 38876
rect 24280 38879 24338 38885
rect 22971 38845 22983 38848
rect 22925 38839 22983 38845
rect 24280 38845 24292 38879
rect 24326 38876 24338 38879
rect 24486 38876 24492 38888
rect 24326 38848 24492 38876
rect 24326 38845 24338 38848
rect 24280 38839 24338 38845
rect 24486 38836 24492 38848
rect 24544 38876 24550 38888
rect 24673 38879 24731 38885
rect 24673 38876 24685 38879
rect 24544 38848 24685 38876
rect 24544 38836 24550 38848
rect 24673 38845 24685 38848
rect 24719 38845 24731 38879
rect 24673 38839 24731 38845
rect 25225 38879 25283 38885
rect 25225 38845 25237 38879
rect 25271 38876 25283 38879
rect 25958 38876 25964 38888
rect 25271 38848 25964 38876
rect 25271 38845 25283 38848
rect 25225 38839 25283 38845
rect 25958 38836 25964 38848
rect 26016 38836 26022 38888
rect 27430 38836 27436 38888
rect 27488 38876 27494 38888
rect 27525 38879 27583 38885
rect 27525 38876 27537 38879
rect 27488 38848 27537 38876
rect 27488 38836 27494 38848
rect 27525 38845 27537 38848
rect 27571 38876 27583 38879
rect 27890 38876 27896 38888
rect 27571 38848 27896 38876
rect 27571 38845 27583 38848
rect 27525 38839 27583 38845
rect 27890 38836 27896 38848
rect 27948 38836 27954 38888
rect 28166 38876 28172 38888
rect 28127 38848 28172 38876
rect 28166 38836 28172 38848
rect 28224 38836 28230 38888
rect 30837 38879 30895 38885
rect 30837 38845 30849 38879
rect 30883 38876 30895 38879
rect 31478 38876 31484 38888
rect 30883 38848 31484 38876
rect 30883 38845 30895 38848
rect 30837 38839 30895 38845
rect 31478 38836 31484 38848
rect 31536 38836 31542 38888
rect 33060 38885 33088 38984
rect 33045 38879 33103 38885
rect 33045 38845 33057 38879
rect 33091 38876 33103 38879
rect 33226 38876 33232 38888
rect 33091 38848 33232 38876
rect 33091 38845 33103 38848
rect 33045 38839 33103 38845
rect 33226 38836 33232 38848
rect 33284 38836 33290 38888
rect 33520 38885 33548 39052
rect 34606 39040 34612 39052
rect 34664 39040 34670 39092
rect 36630 39080 36636 39092
rect 36591 39052 36636 39080
rect 36630 39040 36636 39052
rect 36688 39040 36694 39092
rect 36906 39080 36912 39092
rect 36867 39052 36912 39080
rect 36906 39040 36912 39052
rect 36964 39040 36970 39092
rect 38102 39040 38108 39092
rect 38160 39080 38166 39092
rect 38289 39083 38347 39089
rect 38289 39080 38301 39083
rect 38160 39052 38301 39080
rect 38160 39040 38166 39052
rect 38289 39049 38301 39052
rect 38335 39080 38347 39083
rect 40218 39080 40224 39092
rect 38335 39052 38654 39080
rect 40179 39052 40224 39080
rect 38335 39049 38347 39052
rect 38289 39043 38347 39049
rect 36078 38972 36084 39024
rect 36136 39012 36142 39024
rect 37277 39015 37335 39021
rect 37277 39012 37289 39015
rect 36136 38984 37289 39012
rect 36136 38972 36142 38984
rect 37277 38981 37289 38984
rect 37323 38981 37335 39015
rect 37277 38975 37335 38981
rect 33686 38944 33692 38956
rect 33647 38916 33692 38944
rect 33686 38904 33692 38916
rect 33744 38904 33750 38956
rect 33505 38879 33563 38885
rect 33505 38845 33517 38879
rect 33551 38845 33563 38879
rect 33505 38839 33563 38845
rect 24118 38808 24124 38820
rect 24031 38780 24124 38808
rect 24118 38768 24124 38780
rect 24176 38808 24182 38820
rect 24854 38808 24860 38820
rect 24176 38780 24860 38808
rect 24176 38768 24182 38780
rect 24854 38768 24860 38780
rect 24912 38768 24918 38820
rect 25130 38768 25136 38820
rect 25188 38808 25194 38820
rect 25546 38811 25604 38817
rect 25546 38808 25558 38811
rect 25188 38780 25558 38808
rect 25188 38768 25194 38780
rect 25546 38777 25558 38780
rect 25592 38777 25604 38811
rect 25546 38771 25604 38777
rect 27065 38811 27123 38817
rect 27065 38777 27077 38811
rect 27111 38808 27123 38811
rect 27246 38808 27252 38820
rect 27111 38780 27252 38808
rect 27111 38777 27123 38780
rect 27065 38771 27123 38777
rect 27246 38768 27252 38780
rect 27304 38808 27310 38820
rect 28184 38808 28212 38836
rect 27304 38780 28212 38808
rect 28353 38811 28411 38817
rect 27304 38768 27310 38780
rect 28353 38777 28365 38811
rect 28399 38808 28411 38811
rect 28534 38808 28540 38820
rect 28399 38780 28540 38808
rect 28399 38777 28411 38780
rect 28353 38771 28411 38777
rect 28534 38768 28540 38780
rect 28592 38768 28598 38820
rect 29457 38811 29515 38817
rect 29457 38777 29469 38811
rect 29503 38777 29515 38811
rect 29457 38771 29515 38777
rect 20404 38712 22140 38740
rect 24351 38743 24409 38749
rect 20404 38700 20410 38712
rect 24351 38709 24363 38743
rect 24397 38740 24409 38743
rect 24578 38740 24584 38752
rect 24397 38712 24584 38740
rect 24397 38709 24409 38712
rect 24351 38703 24409 38709
rect 24578 38700 24584 38712
rect 24636 38700 24642 38752
rect 26142 38740 26148 38752
rect 26103 38712 26148 38740
rect 26142 38700 26148 38712
rect 26200 38700 26206 38752
rect 29178 38700 29184 38752
rect 29236 38740 29242 38752
rect 29472 38740 29500 38771
rect 30282 38768 30288 38820
rect 30340 38808 30346 38820
rect 30745 38811 30803 38817
rect 30745 38808 30757 38811
rect 30340 38780 30757 38808
rect 30340 38768 30346 38780
rect 30745 38777 30757 38780
rect 30791 38808 30803 38811
rect 31199 38811 31257 38817
rect 31199 38808 31211 38811
rect 30791 38780 31211 38808
rect 30791 38777 30803 38780
rect 30745 38771 30803 38777
rect 31199 38777 31211 38780
rect 31245 38808 31257 38811
rect 31245 38780 32168 38808
rect 31245 38777 31257 38780
rect 31199 38771 31257 38777
rect 32140 38752 32168 38780
rect 33134 38768 33140 38820
rect 33192 38808 33198 38820
rect 33704 38808 33732 38904
rect 35250 38876 35256 38888
rect 35163 38848 35256 38876
rect 35250 38836 35256 38848
rect 35308 38876 35314 38888
rect 35713 38879 35771 38885
rect 35713 38876 35725 38879
rect 35308 38848 35725 38876
rect 35308 38836 35314 38848
rect 35713 38845 35725 38848
rect 35759 38845 35771 38879
rect 37292 38876 37320 38975
rect 38626 38944 38654 39052
rect 40218 39040 40224 39052
rect 40276 39040 40282 39092
rect 40770 39040 40776 39092
rect 40828 39080 40834 39092
rect 41049 39083 41107 39089
rect 41049 39080 41061 39083
rect 40828 39052 41061 39080
rect 40828 39040 40834 39052
rect 41049 39049 41061 39052
rect 41095 39049 41107 39083
rect 41414 39080 41420 39092
rect 41375 39052 41420 39080
rect 41049 39043 41107 39049
rect 41414 39040 41420 39052
rect 41472 39040 41478 39092
rect 42702 39040 42708 39092
rect 42760 39080 42766 39092
rect 42981 39083 43039 39089
rect 42981 39080 42993 39083
rect 42760 39052 42993 39080
rect 42760 39040 42766 39052
rect 42981 39049 42993 39052
rect 43027 39049 43039 39083
rect 43438 39080 43444 39092
rect 43399 39052 43444 39080
rect 42981 39043 43039 39049
rect 43438 39040 43444 39052
rect 43496 39040 43502 39092
rect 39574 38944 39580 38956
rect 38626 38916 39344 38944
rect 39535 38916 39580 38944
rect 37496 38879 37554 38885
rect 37496 38876 37508 38879
rect 37292 38848 37508 38876
rect 35713 38839 35771 38845
rect 37496 38845 37508 38848
rect 37542 38845 37554 38879
rect 38838 38876 38844 38888
rect 38799 38848 38844 38876
rect 37496 38839 37554 38845
rect 38838 38836 38844 38848
rect 38896 38836 38902 38888
rect 39316 38885 39344 38916
rect 39574 38904 39580 38916
rect 39632 38904 39638 38956
rect 39301 38879 39359 38885
rect 39301 38845 39313 38879
rect 39347 38845 39359 38879
rect 39301 38839 39359 38845
rect 40656 38879 40714 38885
rect 40656 38845 40668 38879
rect 40702 38876 40714 38879
rect 41230 38876 41236 38888
rect 40702 38848 41236 38876
rect 40702 38845 40714 38848
rect 40656 38839 40714 38845
rect 41230 38836 41236 38848
rect 41288 38876 41294 38888
rect 41414 38876 41420 38888
rect 41288 38848 41420 38876
rect 41288 38836 41294 38848
rect 41414 38836 41420 38848
rect 41472 38836 41478 38888
rect 41668 38879 41726 38885
rect 41668 38845 41680 38879
rect 41714 38876 41726 38879
rect 41782 38876 41788 38888
rect 41714 38848 41788 38876
rect 41714 38845 41726 38848
rect 41668 38839 41726 38845
rect 41782 38836 41788 38848
rect 41840 38836 41846 38888
rect 43876 38879 43934 38885
rect 43876 38845 43888 38879
rect 43922 38876 43934 38879
rect 44266 38876 44272 38888
rect 43922 38848 44272 38876
rect 43922 38845 43934 38848
rect 43876 38839 43934 38845
rect 44266 38836 44272 38848
rect 44324 38876 44330 38888
rect 44324 38848 44404 38876
rect 44324 38836 44330 38848
rect 36034 38811 36092 38817
rect 36034 38808 36046 38811
rect 33192 38780 33732 38808
rect 35544 38780 36046 38808
rect 33192 38768 33198 38780
rect 35544 38752 35572 38780
rect 36034 38777 36046 38780
rect 36080 38808 36092 38811
rect 38657 38811 38715 38817
rect 38657 38808 38669 38811
rect 36080 38780 38669 38808
rect 36080 38777 36092 38780
rect 36034 38771 36092 38777
rect 38657 38777 38669 38780
rect 38703 38808 38715 38811
rect 39114 38808 39120 38820
rect 38703 38780 39120 38808
rect 38703 38777 38715 38780
rect 38657 38771 38715 38777
rect 39114 38768 39120 38780
rect 39172 38768 39178 38820
rect 31754 38740 31760 38752
rect 29236 38712 29500 38740
rect 31715 38712 31760 38740
rect 29236 38700 29242 38712
rect 31754 38700 31760 38712
rect 31812 38700 31818 38752
rect 32122 38700 32128 38752
rect 32180 38740 32186 38752
rect 33318 38740 33324 38752
rect 32180 38712 33324 38740
rect 32180 38700 32186 38712
rect 33318 38700 33324 38712
rect 33376 38740 33382 38752
rect 33594 38740 33600 38752
rect 33376 38712 33600 38740
rect 33376 38700 33382 38712
rect 33594 38700 33600 38712
rect 33652 38740 33658 38752
rect 34057 38743 34115 38749
rect 34057 38740 34069 38743
rect 33652 38712 34069 38740
rect 33652 38700 33658 38712
rect 34057 38709 34069 38712
rect 34103 38740 34115 38743
rect 35526 38740 35532 38752
rect 34103 38712 35532 38740
rect 34103 38709 34115 38712
rect 34057 38703 34115 38709
rect 35526 38700 35532 38712
rect 35584 38700 35590 38752
rect 37366 38700 37372 38752
rect 37424 38740 37430 38752
rect 37599 38743 37657 38749
rect 37599 38740 37611 38743
rect 37424 38712 37611 38740
rect 37424 38700 37430 38712
rect 37599 38709 37611 38712
rect 37645 38709 37657 38743
rect 38010 38740 38016 38752
rect 37971 38712 38016 38740
rect 37599 38703 37657 38709
rect 38010 38700 38016 38712
rect 38068 38700 38074 38752
rect 40727 38743 40785 38749
rect 40727 38709 40739 38743
rect 40773 38740 40785 38743
rect 40954 38740 40960 38752
rect 40773 38712 40960 38740
rect 40773 38709 40785 38712
rect 40727 38703 40785 38709
rect 40954 38700 40960 38712
rect 41012 38700 41018 38752
rect 41739 38743 41797 38749
rect 41739 38709 41751 38743
rect 41785 38740 41797 38743
rect 41966 38740 41972 38752
rect 41785 38712 41972 38740
rect 41785 38709 41797 38712
rect 41739 38703 41797 38709
rect 41966 38700 41972 38712
rect 42024 38700 42030 38752
rect 42334 38740 42340 38752
rect 42295 38712 42340 38740
rect 42334 38700 42340 38712
rect 42392 38700 42398 38752
rect 43947 38743 44005 38749
rect 43947 38709 43959 38743
rect 43993 38740 44005 38743
rect 44174 38740 44180 38752
rect 43993 38712 44180 38740
rect 43993 38709 44005 38712
rect 43947 38703 44005 38709
rect 44174 38700 44180 38712
rect 44232 38700 44238 38752
rect 44376 38749 44404 38848
rect 44361 38743 44419 38749
rect 44361 38709 44373 38743
rect 44407 38740 44419 38743
rect 44450 38740 44456 38752
rect 44407 38712 44456 38740
rect 44407 38709 44419 38712
rect 44361 38703 44419 38709
rect 44450 38700 44456 38712
rect 44508 38700 44514 38752
rect 1104 38650 48852 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 48852 38650
rect 1104 38576 48852 38598
rect 16482 38536 16488 38548
rect 16443 38508 16488 38536
rect 16482 38496 16488 38508
rect 16540 38496 16546 38548
rect 16758 38536 16764 38548
rect 16719 38508 16764 38536
rect 16758 38496 16764 38508
rect 16816 38496 16822 38548
rect 17954 38536 17960 38548
rect 17915 38508 17960 38536
rect 17954 38496 17960 38508
rect 18012 38496 18018 38548
rect 19426 38496 19432 38548
rect 19484 38536 19490 38548
rect 19521 38539 19579 38545
rect 19521 38536 19533 38539
rect 19484 38508 19533 38536
rect 19484 38496 19490 38508
rect 19521 38505 19533 38508
rect 19567 38505 19579 38539
rect 21174 38536 21180 38548
rect 21135 38508 21180 38536
rect 19521 38499 19579 38505
rect 21174 38496 21180 38508
rect 21232 38496 21238 38548
rect 22278 38496 22284 38548
rect 22336 38536 22342 38548
rect 24486 38536 24492 38548
rect 22336 38508 24492 38536
rect 22336 38496 22342 38508
rect 24486 38496 24492 38508
rect 24544 38496 24550 38548
rect 25958 38536 25964 38548
rect 25919 38508 25964 38536
rect 25958 38496 25964 38508
rect 26016 38496 26022 38548
rect 28258 38536 28264 38548
rect 28219 38508 28264 38536
rect 28258 38496 28264 38508
rect 28316 38496 28322 38548
rect 31846 38536 31852 38548
rect 31807 38508 31852 38536
rect 31846 38496 31852 38508
rect 31904 38496 31910 38548
rect 32493 38539 32551 38545
rect 32493 38505 32505 38539
rect 32539 38505 32551 38539
rect 35250 38536 35256 38548
rect 35211 38508 35256 38536
rect 32493 38499 32551 38505
rect 13814 38468 13820 38480
rect 13786 38428 13820 38468
rect 13872 38468 13878 38480
rect 14829 38471 14887 38477
rect 14829 38468 14841 38471
rect 13872 38440 14841 38468
rect 13872 38428 13878 38440
rect 14829 38437 14841 38440
rect 14875 38468 14887 38471
rect 15562 38468 15568 38480
rect 14875 38440 15568 38468
rect 14875 38437 14887 38440
rect 14829 38431 14887 38437
rect 15562 38428 15568 38440
rect 15620 38468 15626 38480
rect 16114 38468 16120 38480
rect 15620 38440 15976 38468
rect 16075 38440 16120 38468
rect 15620 38428 15626 38440
rect 13265 38335 13323 38341
rect 13265 38301 13277 38335
rect 13311 38332 13323 38335
rect 13786 38332 13814 38428
rect 15654 38400 15660 38412
rect 15615 38372 15660 38400
rect 15654 38360 15660 38372
rect 15712 38360 15718 38412
rect 15948 38409 15976 38440
rect 16114 38428 16120 38440
rect 16172 38428 16178 38480
rect 15933 38403 15991 38409
rect 15933 38369 15945 38403
rect 15979 38400 15991 38403
rect 16500 38400 16528 38496
rect 18874 38468 18880 38480
rect 18835 38440 18880 38468
rect 18874 38428 18880 38440
rect 18932 38428 18938 38480
rect 23014 38428 23020 38480
rect 23072 38468 23078 38480
rect 23338 38471 23396 38477
rect 23338 38468 23350 38471
rect 23072 38440 23350 38468
rect 23072 38428 23078 38440
rect 23338 38437 23350 38440
rect 23384 38437 23396 38471
rect 24946 38468 24952 38480
rect 24907 38440 24952 38468
rect 23338 38431 23396 38437
rect 24946 38428 24952 38440
rect 25004 38428 25010 38480
rect 25041 38471 25099 38477
rect 25041 38437 25053 38471
rect 25087 38468 25099 38471
rect 26142 38468 26148 38480
rect 25087 38440 26148 38468
rect 25087 38437 25099 38440
rect 25041 38431 25099 38437
rect 26142 38428 26148 38440
rect 26200 38468 26206 38480
rect 26602 38468 26608 38480
rect 26200 38440 26608 38468
rect 26200 38428 26206 38440
rect 26602 38428 26608 38440
rect 26660 38468 26666 38480
rect 26697 38471 26755 38477
rect 26697 38468 26709 38471
rect 26660 38440 26709 38468
rect 26660 38428 26666 38440
rect 26697 38437 26709 38440
rect 26743 38437 26755 38471
rect 26697 38431 26755 38437
rect 28718 38428 28724 38480
rect 28776 38468 28782 38480
rect 28858 38471 28916 38477
rect 28858 38468 28870 38471
rect 28776 38440 28870 38468
rect 28776 38428 28782 38440
rect 28858 38437 28870 38440
rect 28904 38468 28916 38471
rect 30282 38468 30288 38480
rect 28904 38440 30288 38468
rect 28904 38437 28916 38440
rect 28858 38431 28916 38437
rect 30282 38428 30288 38440
rect 30340 38428 30346 38480
rect 30374 38428 30380 38480
rect 30432 38468 30438 38480
rect 30653 38471 30711 38477
rect 30653 38468 30665 38471
rect 30432 38440 30665 38468
rect 30432 38428 30438 38440
rect 30653 38437 30665 38440
rect 30699 38468 30711 38471
rect 31754 38468 31760 38480
rect 30699 38440 31760 38468
rect 30699 38437 30711 38440
rect 30653 38431 30711 38437
rect 31754 38428 31760 38440
rect 31812 38428 31818 38480
rect 15979 38372 16528 38400
rect 15979 38369 15991 38372
rect 15933 38363 15991 38369
rect 17862 38360 17868 38412
rect 17920 38400 17926 38412
rect 18141 38403 18199 38409
rect 18141 38400 18153 38403
rect 17920 38372 18153 38400
rect 17920 38360 17926 38372
rect 18141 38369 18153 38372
rect 18187 38369 18199 38403
rect 18141 38363 18199 38369
rect 18693 38403 18751 38409
rect 18693 38369 18705 38403
rect 18739 38400 18751 38403
rect 19150 38400 19156 38412
rect 18739 38372 19156 38400
rect 18739 38369 18751 38372
rect 18693 38363 18751 38369
rect 19150 38360 19156 38372
rect 19208 38360 19214 38412
rect 19864 38403 19922 38409
rect 19864 38369 19876 38403
rect 19910 38400 19922 38403
rect 20530 38400 20536 38412
rect 19910 38372 20536 38400
rect 19910 38369 19922 38372
rect 19864 38363 19922 38369
rect 20530 38360 20536 38372
rect 20588 38360 20594 38412
rect 20898 38400 20904 38412
rect 20859 38372 20904 38400
rect 20898 38360 20904 38372
rect 20956 38360 20962 38412
rect 21358 38400 21364 38412
rect 21319 38372 21364 38400
rect 21358 38360 21364 38372
rect 21416 38360 21422 38412
rect 32125 38403 32183 38409
rect 32125 38369 32137 38403
rect 32171 38400 32183 38403
rect 32214 38400 32220 38412
rect 32171 38372 32220 38400
rect 32171 38369 32183 38372
rect 32125 38363 32183 38369
rect 32214 38360 32220 38372
rect 32272 38360 32278 38412
rect 32508 38400 32536 38499
rect 35250 38496 35256 38508
rect 35308 38496 35314 38548
rect 36817 38539 36875 38545
rect 36817 38505 36829 38539
rect 36863 38536 36875 38539
rect 38010 38536 38016 38548
rect 36863 38508 38016 38536
rect 36863 38505 36875 38508
rect 36817 38499 36875 38505
rect 38010 38496 38016 38508
rect 38068 38496 38074 38548
rect 38838 38536 38844 38548
rect 38120 38508 38844 38536
rect 33318 38428 33324 38480
rect 33376 38468 33382 38480
rect 38120 38468 38148 38508
rect 38838 38496 38844 38508
rect 38896 38496 38902 38548
rect 33376 38440 38148 38468
rect 38473 38471 38531 38477
rect 33376 38428 33382 38440
rect 38473 38437 38485 38471
rect 38519 38468 38531 38471
rect 38746 38468 38752 38480
rect 38519 38440 38752 38468
rect 38519 38437 38531 38440
rect 38473 38431 38531 38437
rect 38746 38428 38752 38440
rect 38804 38468 38810 38480
rect 39209 38471 39267 38477
rect 39209 38468 39221 38471
rect 38804 38440 39221 38468
rect 38804 38428 38810 38440
rect 39209 38437 39221 38440
rect 39255 38437 39267 38471
rect 39209 38431 39267 38437
rect 40954 38428 40960 38480
rect 41012 38468 41018 38480
rect 41782 38468 41788 38480
rect 41012 38440 41788 38468
rect 41012 38428 41018 38440
rect 41782 38428 41788 38440
rect 41840 38428 41846 38480
rect 41874 38428 41880 38480
rect 41932 38468 41938 38480
rect 44085 38471 44143 38477
rect 41932 38440 41977 38468
rect 41932 38428 41938 38440
rect 44085 38437 44097 38471
rect 44131 38468 44143 38471
rect 44266 38468 44272 38480
rect 44131 38440 44272 38468
rect 44131 38437 44143 38440
rect 44085 38431 44143 38437
rect 44266 38428 44272 38440
rect 44324 38428 44330 38480
rect 33594 38400 33600 38412
rect 32508 38372 33600 38400
rect 33594 38360 33600 38372
rect 33652 38360 33658 38412
rect 33962 38400 33968 38412
rect 33923 38372 33968 38400
rect 33962 38360 33968 38372
rect 34020 38360 34026 38412
rect 35250 38400 35256 38412
rect 35211 38372 35256 38400
rect 35250 38360 35256 38372
rect 35308 38360 35314 38412
rect 35434 38400 35440 38412
rect 35395 38372 35440 38400
rect 35434 38360 35440 38372
rect 35492 38360 35498 38412
rect 36633 38403 36691 38409
rect 36633 38369 36645 38403
rect 36679 38400 36691 38403
rect 36906 38400 36912 38412
rect 36679 38372 36912 38400
rect 36679 38369 36691 38372
rect 36633 38363 36691 38369
rect 36906 38360 36912 38372
rect 36964 38360 36970 38412
rect 37734 38400 37740 38412
rect 37695 38372 37740 38400
rect 37734 38360 37740 38372
rect 37792 38360 37798 38412
rect 38010 38360 38016 38412
rect 38068 38400 38074 38412
rect 38289 38403 38347 38409
rect 38289 38400 38301 38403
rect 38068 38372 38301 38400
rect 38068 38360 38074 38372
rect 38289 38369 38301 38372
rect 38335 38400 38347 38403
rect 39022 38400 39028 38412
rect 38335 38372 39028 38400
rect 38335 38369 38347 38372
rect 38289 38363 38347 38369
rect 39022 38360 39028 38372
rect 39080 38360 39086 38412
rect 40310 38360 40316 38412
rect 40368 38400 40374 38412
rect 40624 38403 40682 38409
rect 40624 38400 40636 38403
rect 40368 38372 40636 38400
rect 40368 38360 40374 38372
rect 40624 38369 40636 38372
rect 40670 38369 40682 38403
rect 40624 38363 40682 38369
rect 13311 38304 13814 38332
rect 23017 38335 23075 38341
rect 13311 38301 13323 38304
rect 13265 38295 13323 38301
rect 23017 38301 23029 38335
rect 23063 38301 23075 38335
rect 23017 38295 23075 38301
rect 17034 38196 17040 38208
rect 16995 38168 17040 38196
rect 17034 38156 17040 38168
rect 17092 38156 17098 38208
rect 17267 38199 17325 38205
rect 17267 38165 17279 38199
rect 17313 38196 17325 38199
rect 17770 38196 17776 38208
rect 17313 38168 17776 38196
rect 17313 38165 17325 38168
rect 17267 38159 17325 38165
rect 17770 38156 17776 38168
rect 17828 38156 17834 38208
rect 19935 38199 19993 38205
rect 19935 38165 19947 38199
rect 19981 38196 19993 38199
rect 20714 38196 20720 38208
rect 19981 38168 20720 38196
rect 19981 38165 19993 38168
rect 19935 38159 19993 38165
rect 20714 38156 20720 38168
rect 20772 38156 20778 38208
rect 22738 38156 22744 38208
rect 22796 38196 22802 38208
rect 22833 38199 22891 38205
rect 22833 38196 22845 38199
rect 22796 38168 22845 38196
rect 22796 38156 22802 38168
rect 22833 38165 22845 38168
rect 22879 38196 22891 38199
rect 23032 38196 23060 38295
rect 24578 38292 24584 38344
rect 24636 38332 24642 38344
rect 26605 38335 26663 38341
rect 26605 38332 26617 38335
rect 24636 38304 26617 38332
rect 24636 38292 24642 38304
rect 26605 38301 26617 38304
rect 26651 38332 26663 38335
rect 26970 38332 26976 38344
rect 26651 38304 26976 38332
rect 26651 38301 26663 38304
rect 26605 38295 26663 38301
rect 26970 38292 26976 38304
rect 27028 38292 27034 38344
rect 27249 38335 27307 38341
rect 27249 38301 27261 38335
rect 27295 38332 27307 38335
rect 28350 38332 28356 38344
rect 27295 38304 28356 38332
rect 27295 38301 27307 38304
rect 27249 38295 27307 38301
rect 28350 38292 28356 38304
rect 28408 38292 28414 38344
rect 28534 38332 28540 38344
rect 28495 38304 28540 38332
rect 28534 38292 28540 38304
rect 28592 38292 28598 38344
rect 30561 38335 30619 38341
rect 30561 38301 30573 38335
rect 30607 38301 30619 38335
rect 30561 38295 30619 38301
rect 25501 38267 25559 38273
rect 25501 38233 25513 38267
rect 25547 38264 25559 38267
rect 26234 38264 26240 38276
rect 25547 38236 26240 38264
rect 25547 38233 25559 38236
rect 25501 38227 25559 38233
rect 26234 38224 26240 38236
rect 26292 38224 26298 38276
rect 30466 38224 30472 38276
rect 30524 38264 30530 38276
rect 30576 38264 30604 38295
rect 31202 38292 31208 38344
rect 31260 38332 31266 38344
rect 33502 38332 33508 38344
rect 31260 38304 33508 38332
rect 31260 38292 31266 38304
rect 33502 38292 33508 38304
rect 33560 38292 33566 38344
rect 39485 38335 39543 38341
rect 39485 38301 39497 38335
rect 39531 38332 39543 38335
rect 39666 38332 39672 38344
rect 39531 38304 39672 38332
rect 39531 38301 39543 38304
rect 39485 38295 39543 38301
rect 39666 38292 39672 38304
rect 39724 38292 39730 38344
rect 43990 38332 43996 38344
rect 43951 38304 43996 38332
rect 43990 38292 43996 38304
rect 44048 38292 44054 38344
rect 44637 38335 44695 38341
rect 44637 38301 44649 38335
rect 44683 38332 44695 38335
rect 46198 38332 46204 38344
rect 44683 38304 46204 38332
rect 44683 38301 44695 38304
rect 44637 38295 44695 38301
rect 30524 38236 30604 38264
rect 31113 38267 31171 38273
rect 30524 38224 30530 38236
rect 31113 38233 31125 38267
rect 31159 38264 31171 38267
rect 31570 38264 31576 38276
rect 31159 38236 31576 38264
rect 31159 38233 31171 38236
rect 31113 38227 31171 38233
rect 31570 38224 31576 38236
rect 31628 38224 31634 38276
rect 32858 38224 32864 38276
rect 32916 38264 32922 38276
rect 34149 38267 34207 38273
rect 34149 38264 34161 38267
rect 32916 38236 34161 38264
rect 32916 38224 32922 38236
rect 34149 38233 34161 38236
rect 34195 38233 34207 38267
rect 41417 38267 41475 38273
rect 41417 38264 41429 38267
rect 34149 38227 34207 38233
rect 40604 38236 41429 38264
rect 40604 38208 40632 38236
rect 41417 38233 41429 38236
rect 41463 38233 41475 38267
rect 41417 38227 41475 38233
rect 42337 38267 42395 38273
rect 42337 38233 42349 38267
rect 42383 38264 42395 38267
rect 43622 38264 43628 38276
rect 42383 38236 43628 38264
rect 42383 38233 42395 38236
rect 42337 38227 42395 38233
rect 43622 38224 43628 38236
rect 43680 38264 43686 38276
rect 44652 38264 44680 38295
rect 46198 38292 46204 38304
rect 46256 38292 46262 38344
rect 43680 38236 44680 38264
rect 43680 38224 43686 38236
rect 23934 38196 23940 38208
rect 22879 38168 23060 38196
rect 23895 38168 23940 38196
rect 22879 38165 22891 38168
rect 22833 38159 22891 38165
rect 23934 38156 23940 38168
rect 23992 38156 23998 38208
rect 27709 38199 27767 38205
rect 27709 38165 27721 38199
rect 27755 38196 27767 38199
rect 28166 38196 28172 38208
rect 27755 38168 28172 38196
rect 27755 38165 27767 38168
rect 27709 38159 27767 38165
rect 28166 38156 28172 38168
rect 28224 38156 28230 38208
rect 29454 38196 29460 38208
rect 29415 38168 29460 38196
rect 29454 38156 29460 38168
rect 29512 38156 29518 38208
rect 31478 38196 31484 38208
rect 31439 38168 31484 38196
rect 31478 38156 31484 38168
rect 31536 38156 31542 38208
rect 33042 38196 33048 38208
rect 33003 38168 33048 38196
rect 33042 38156 33048 38168
rect 33100 38156 33106 38208
rect 33134 38156 33140 38208
rect 33192 38196 33198 38208
rect 33689 38199 33747 38205
rect 33689 38196 33701 38199
rect 33192 38168 33701 38196
rect 33192 38156 33198 38168
rect 33689 38165 33701 38168
rect 33735 38165 33747 38199
rect 35986 38196 35992 38208
rect 35947 38168 35992 38196
rect 33689 38159 33747 38165
rect 35986 38156 35992 38168
rect 36044 38156 36050 38208
rect 39715 38199 39773 38205
rect 39715 38165 39727 38199
rect 39761 38196 39773 38199
rect 40586 38196 40592 38208
rect 39761 38168 40592 38196
rect 39761 38165 39773 38168
rect 39715 38159 39773 38165
rect 40586 38156 40592 38168
rect 40644 38156 40650 38208
rect 40727 38199 40785 38205
rect 40727 38165 40739 38199
rect 40773 38196 40785 38199
rect 40862 38196 40868 38208
rect 40773 38168 40868 38196
rect 40773 38165 40785 38168
rect 40727 38159 40785 38165
rect 40862 38156 40868 38168
rect 40920 38156 40926 38208
rect 41046 38196 41052 38208
rect 41007 38168 41052 38196
rect 41046 38156 41052 38168
rect 41104 38156 41110 38208
rect 1104 38106 48852 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 48852 38106
rect 1104 38032 48852 38054
rect 15654 37952 15660 38004
rect 15712 37992 15718 38004
rect 15749 37995 15807 38001
rect 15749 37992 15761 37995
rect 15712 37964 15761 37992
rect 15712 37952 15718 37964
rect 15749 37961 15761 37964
rect 15795 37961 15807 37995
rect 15749 37955 15807 37961
rect 17865 37995 17923 38001
rect 17865 37961 17877 37995
rect 17911 37992 17923 37995
rect 18046 37992 18052 38004
rect 17911 37964 18052 37992
rect 17911 37961 17923 37964
rect 17865 37955 17923 37961
rect 18046 37952 18052 37964
rect 18104 37952 18110 38004
rect 18601 37995 18659 38001
rect 18601 37961 18613 37995
rect 18647 37992 18659 37995
rect 20162 37992 20168 38004
rect 18647 37964 20168 37992
rect 18647 37961 18659 37964
rect 18601 37955 18659 37961
rect 15473 37927 15531 37933
rect 15473 37893 15485 37927
rect 15519 37924 15531 37927
rect 15930 37924 15936 37936
rect 15519 37896 15936 37924
rect 15519 37893 15531 37896
rect 15473 37887 15531 37893
rect 14988 37791 15046 37797
rect 14988 37757 15000 37791
rect 15034 37788 15046 37791
rect 15194 37788 15200 37800
rect 15034 37760 15200 37788
rect 15034 37757 15046 37760
rect 14988 37751 15046 37757
rect 15194 37748 15200 37760
rect 15252 37788 15258 37800
rect 15488 37788 15516 37887
rect 15930 37884 15936 37896
rect 15988 37884 15994 37936
rect 16574 37924 16580 37936
rect 16535 37896 16580 37924
rect 16574 37884 16580 37896
rect 16632 37884 16638 37936
rect 15252 37760 15516 37788
rect 18116 37791 18174 37797
rect 15252 37748 15258 37760
rect 18116 37757 18128 37791
rect 18162 37788 18174 37791
rect 18616 37788 18644 37955
rect 20162 37952 20168 37964
rect 20220 37952 20226 38004
rect 21358 37992 21364 38004
rect 21319 37964 21364 37992
rect 21358 37952 21364 37964
rect 21416 37952 21422 38004
rect 26602 37992 26608 38004
rect 26563 37964 26608 37992
rect 26602 37952 26608 37964
rect 26660 37952 26666 38004
rect 26970 37992 26976 38004
rect 26931 37964 26976 37992
rect 26970 37952 26976 37964
rect 27028 37952 27034 38004
rect 27062 37952 27068 38004
rect 27120 37992 27126 38004
rect 27433 37995 27491 38001
rect 27433 37992 27445 37995
rect 27120 37964 27445 37992
rect 27120 37952 27126 37964
rect 27433 37961 27445 37964
rect 27479 37992 27491 37995
rect 27614 37992 27620 38004
rect 27479 37964 27620 37992
rect 27479 37961 27491 37964
rect 27433 37955 27491 37961
rect 27614 37952 27620 37964
rect 27672 37952 27678 38004
rect 28718 37992 28724 38004
rect 28679 37964 28724 37992
rect 28718 37952 28724 37964
rect 28776 37952 28782 38004
rect 29638 37992 29644 38004
rect 28966 37964 29644 37992
rect 18690 37884 18696 37936
rect 18748 37924 18754 37936
rect 20898 37924 20904 37936
rect 18748 37896 20904 37924
rect 18748 37884 18754 37896
rect 20898 37884 20904 37896
rect 20956 37884 20962 37936
rect 26786 37884 26792 37936
rect 26844 37924 26850 37936
rect 28966 37924 28994 37964
rect 29638 37952 29644 37964
rect 29696 37992 29702 38004
rect 30374 37992 30380 38004
rect 29696 37964 29960 37992
rect 30335 37964 30380 37992
rect 29696 37952 29702 37964
rect 29932 37933 29960 37964
rect 30374 37952 30380 37964
rect 30432 37952 30438 38004
rect 32122 37992 32128 38004
rect 32083 37964 32128 37992
rect 32122 37952 32128 37964
rect 32180 37952 32186 38004
rect 32214 37952 32220 38004
rect 32272 37992 32278 38004
rect 33597 37995 33655 38001
rect 33597 37992 33609 37995
rect 32272 37964 33609 37992
rect 32272 37952 32278 37964
rect 33597 37961 33609 37964
rect 33643 37961 33655 37995
rect 33962 37992 33968 38004
rect 33923 37964 33968 37992
rect 33597 37955 33655 37961
rect 33962 37952 33968 37964
rect 34020 37992 34026 38004
rect 35069 37995 35127 38001
rect 35069 37992 35081 37995
rect 34020 37964 35081 37992
rect 34020 37952 34026 37964
rect 35069 37961 35081 37964
rect 35115 37992 35127 37995
rect 35434 37992 35440 38004
rect 35115 37964 35440 37992
rect 35115 37961 35127 37964
rect 35069 37955 35127 37961
rect 35434 37952 35440 37964
rect 35492 37952 35498 38004
rect 35526 37952 35532 38004
rect 35584 37992 35590 38004
rect 35584 37964 35629 37992
rect 35584 37952 35590 37964
rect 36446 37952 36452 38004
rect 36504 37992 36510 38004
rect 36541 37995 36599 38001
rect 36541 37992 36553 37995
rect 36504 37964 36553 37992
rect 36504 37952 36510 37964
rect 36541 37961 36553 37964
rect 36587 37961 36599 37995
rect 39022 37992 39028 38004
rect 38983 37964 39028 37992
rect 36541 37955 36599 37961
rect 39022 37952 39028 37964
rect 39080 37952 39086 38004
rect 40310 37992 40316 38004
rect 40271 37964 40316 37992
rect 40310 37952 40316 37964
rect 40368 37992 40374 38004
rect 43898 37992 43904 38004
rect 40368 37964 43904 37992
rect 40368 37952 40374 37964
rect 43898 37952 43904 37964
rect 43956 37952 43962 38004
rect 44082 37952 44088 38004
rect 44140 37992 44146 38004
rect 44634 37992 44640 38004
rect 44140 37964 44640 37992
rect 44140 37952 44146 37964
rect 44634 37952 44640 37964
rect 44692 37992 44698 38004
rect 46569 37995 46627 38001
rect 46569 37992 46581 37995
rect 44692 37964 46581 37992
rect 44692 37952 44698 37964
rect 26844 37896 28994 37924
rect 29917 37927 29975 37933
rect 26844 37884 26850 37896
rect 29917 37893 29929 37927
rect 29963 37924 29975 37927
rect 42981 37927 43039 37933
rect 29963 37896 31616 37924
rect 29963 37893 29975 37896
rect 29917 37887 29975 37893
rect 31588 37868 31616 37896
rect 42981 37893 42993 37927
rect 43027 37924 43039 37927
rect 44726 37924 44732 37936
rect 43027 37896 44732 37924
rect 43027 37893 43039 37896
rect 42981 37887 43039 37893
rect 44726 37884 44732 37896
rect 44784 37884 44790 37936
rect 19426 37816 19432 37868
rect 19484 37856 19490 37868
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19484 37828 19625 37856
rect 19484 37816 19490 37828
rect 19613 37825 19625 37828
rect 19659 37825 19671 37859
rect 19886 37856 19892 37868
rect 19847 37828 19892 37856
rect 19613 37819 19671 37825
rect 19886 37816 19892 37828
rect 19944 37816 19950 37868
rect 22738 37856 22744 37868
rect 22699 37828 22744 37856
rect 22738 37816 22744 37828
rect 22796 37816 22802 37868
rect 28258 37856 28264 37868
rect 28219 37828 28264 37856
rect 28258 37816 28264 37828
rect 28316 37816 28322 37868
rect 31478 37856 31484 37868
rect 31439 37828 31484 37856
rect 31478 37816 31484 37828
rect 31536 37816 31542 37868
rect 31570 37816 31576 37868
rect 31628 37856 31634 37868
rect 32953 37859 33011 37865
rect 32953 37856 32965 37859
rect 31628 37828 32965 37856
rect 31628 37816 31634 37828
rect 32953 37825 32965 37828
rect 32999 37825 33011 37859
rect 32953 37819 33011 37825
rect 35621 37859 35679 37865
rect 35621 37825 35633 37859
rect 35667 37856 35679 37859
rect 35986 37856 35992 37868
rect 35667 37828 35992 37856
rect 35667 37825 35679 37828
rect 35621 37819 35679 37825
rect 35986 37816 35992 37828
rect 36044 37816 36050 37868
rect 40586 37816 40592 37868
rect 40644 37856 40650 37868
rect 40865 37859 40923 37865
rect 40865 37856 40877 37859
rect 40644 37828 40877 37856
rect 40644 37816 40650 37828
rect 40865 37825 40877 37828
rect 40911 37825 40923 37859
rect 44174 37856 44180 37868
rect 44135 37828 44180 37856
rect 40865 37819 40923 37825
rect 44174 37816 44180 37828
rect 44232 37856 44238 37868
rect 45097 37859 45155 37865
rect 45097 37856 45109 37859
rect 44232 37828 45109 37856
rect 44232 37816 44238 37828
rect 45097 37825 45109 37828
rect 45143 37825 45155 37859
rect 45097 37819 45155 37825
rect 22002 37788 22008 37800
rect 18162 37760 18644 37788
rect 21963 37760 22008 37788
rect 18162 37757 18174 37760
rect 18116 37751 18174 37757
rect 22002 37748 22008 37760
rect 22060 37748 22066 37800
rect 22465 37791 22523 37797
rect 22465 37757 22477 37791
rect 22511 37757 22523 37791
rect 23658 37788 23664 37800
rect 23619 37760 23664 37788
rect 22465 37751 22523 37757
rect 14829 37723 14887 37729
rect 14829 37689 14841 37723
rect 14875 37720 14887 37723
rect 15470 37720 15476 37732
rect 14875 37692 15476 37720
rect 14875 37689 14887 37692
rect 14829 37683 14887 37689
rect 15470 37680 15476 37692
rect 15528 37720 15534 37732
rect 16025 37723 16083 37729
rect 16025 37720 16037 37723
rect 15528 37692 16037 37720
rect 15528 37680 15534 37692
rect 16025 37689 16037 37692
rect 16071 37689 16083 37723
rect 16025 37683 16083 37689
rect 16114 37680 16120 37732
rect 16172 37720 16178 37732
rect 16172 37692 16217 37720
rect 16172 37680 16178 37692
rect 17862 37680 17868 37732
rect 17920 37720 17926 37732
rect 18877 37723 18935 37729
rect 18877 37720 18889 37723
rect 17920 37692 18889 37720
rect 17920 37680 17926 37692
rect 18877 37689 18889 37692
rect 18923 37689 18935 37723
rect 18877 37683 18935 37689
rect 19705 37723 19763 37729
rect 19705 37689 19717 37723
rect 19751 37689 19763 37723
rect 22480 37720 22508 37751
rect 23658 37748 23664 37760
rect 23716 37748 23722 37800
rect 27614 37788 27620 37800
rect 27575 37760 27620 37788
rect 27614 37748 27620 37760
rect 27672 37748 27678 37800
rect 28166 37788 28172 37800
rect 28079 37760 28172 37788
rect 28166 37748 28172 37760
rect 28224 37788 28230 37800
rect 29178 37788 29184 37800
rect 28224 37760 29184 37788
rect 28224 37748 28230 37760
rect 29178 37748 29184 37760
rect 29236 37748 29242 37800
rect 30745 37791 30803 37797
rect 30745 37757 30757 37791
rect 30791 37788 30803 37791
rect 31113 37791 31171 37797
rect 31113 37788 31125 37791
rect 30791 37760 31125 37788
rect 30791 37757 30803 37760
rect 30745 37751 30803 37757
rect 31113 37757 31125 37760
rect 31159 37788 31171 37791
rect 31202 37788 31208 37800
rect 31159 37760 31208 37788
rect 31159 37757 31171 37760
rect 31113 37751 31171 37757
rect 31202 37748 31208 37760
rect 31260 37748 31266 37800
rect 31294 37748 31300 37800
rect 31352 37788 31358 37800
rect 31389 37791 31447 37797
rect 31389 37788 31401 37791
rect 31352 37760 31401 37788
rect 31352 37748 31358 37760
rect 31389 37757 31401 37760
rect 31435 37788 31447 37791
rect 31846 37788 31852 37800
rect 31435 37760 31852 37788
rect 31435 37757 31447 37760
rect 31389 37751 31447 37757
rect 31846 37748 31852 37760
rect 31904 37748 31910 37800
rect 37921 37791 37979 37797
rect 37921 37757 37933 37791
rect 37967 37788 37979 37791
rect 38286 37788 38292 37800
rect 37967 37760 38292 37788
rect 37967 37757 37979 37760
rect 37921 37751 37979 37757
rect 38286 37748 38292 37760
rect 38344 37748 38350 37800
rect 38470 37788 38476 37800
rect 38431 37760 38476 37788
rect 38470 37748 38476 37760
rect 38528 37748 38534 37800
rect 46159 37797 46187 37964
rect 46569 37961 46581 37964
rect 46615 37961 46627 37995
rect 46569 37955 46627 37961
rect 46144 37791 46202 37797
rect 46144 37757 46156 37791
rect 46190 37757 46202 37791
rect 46144 37751 46202 37757
rect 23982 37723 24040 37729
rect 23982 37720 23994 37723
rect 19705 37683 19763 37689
rect 21836 37692 22508 37720
rect 23400 37692 23994 37720
rect 15059 37655 15117 37661
rect 15059 37621 15071 37655
rect 15105 37652 15117 37655
rect 15286 37652 15292 37664
rect 15105 37624 15292 37652
rect 15105 37621 15117 37624
rect 15059 37615 15117 37621
rect 15286 37612 15292 37624
rect 15344 37612 15350 37664
rect 17034 37612 17040 37664
rect 17092 37652 17098 37664
rect 17221 37655 17279 37661
rect 17221 37652 17233 37655
rect 17092 37624 17233 37652
rect 17092 37612 17098 37624
rect 17221 37621 17233 37624
rect 17267 37652 17279 37655
rect 18046 37652 18052 37664
rect 17267 37624 18052 37652
rect 17267 37621 17279 37624
rect 17221 37615 17279 37621
rect 18046 37612 18052 37624
rect 18104 37612 18110 37664
rect 18187 37655 18245 37661
rect 18187 37621 18199 37655
rect 18233 37652 18245 37655
rect 18414 37652 18420 37664
rect 18233 37624 18420 37652
rect 18233 37621 18245 37624
rect 18187 37615 18245 37621
rect 18414 37612 18420 37624
rect 18472 37612 18478 37664
rect 19426 37652 19432 37664
rect 19387 37624 19432 37652
rect 19426 37612 19432 37624
rect 19484 37652 19490 37664
rect 19720 37652 19748 37683
rect 21836 37664 21864 37692
rect 20530 37652 20536 37664
rect 19484 37624 19748 37652
rect 20491 37624 20536 37652
rect 19484 37612 19490 37624
rect 20530 37612 20536 37624
rect 20588 37612 20594 37664
rect 21818 37652 21824 37664
rect 21779 37624 21824 37652
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 23014 37652 23020 37664
rect 22927 37624 23020 37652
rect 23014 37612 23020 37624
rect 23072 37652 23078 37664
rect 23400 37661 23428 37692
rect 23982 37689 23994 37692
rect 24028 37689 24040 37723
rect 25682 37720 25688 37732
rect 25643 37692 25688 37720
rect 23982 37683 24040 37689
rect 25682 37680 25688 37692
rect 25740 37680 25746 37732
rect 25777 37723 25835 37729
rect 25777 37689 25789 37723
rect 25823 37720 25835 37723
rect 26142 37720 26148 37732
rect 25823 37692 26148 37720
rect 25823 37689 25835 37692
rect 25777 37683 25835 37689
rect 23385 37655 23443 37661
rect 23385 37652 23397 37655
rect 23072 37624 23397 37652
rect 23072 37612 23078 37624
rect 23385 37621 23397 37624
rect 23431 37621 23443 37655
rect 23385 37615 23443 37621
rect 23842 37612 23848 37664
rect 23900 37652 23906 37664
rect 24581 37655 24639 37661
rect 24581 37652 24593 37655
rect 23900 37624 24593 37652
rect 23900 37612 23906 37624
rect 24581 37621 24593 37624
rect 24627 37621 24639 37655
rect 24581 37615 24639 37621
rect 24949 37655 25007 37661
rect 24949 37621 24961 37655
rect 24995 37652 25007 37655
rect 25501 37655 25559 37661
rect 25501 37652 25513 37655
rect 24995 37624 25513 37652
rect 24995 37621 25007 37624
rect 24949 37615 25007 37621
rect 25501 37621 25513 37624
rect 25547 37652 25559 37655
rect 25792 37652 25820 37683
rect 26142 37680 26148 37692
rect 26200 37680 26206 37732
rect 26329 37723 26387 37729
rect 26329 37689 26341 37723
rect 26375 37720 26387 37723
rect 26878 37720 26884 37732
rect 26375 37692 26884 37720
rect 26375 37689 26387 37692
rect 26329 37683 26387 37689
rect 26878 37680 26884 37692
rect 26936 37680 26942 37732
rect 29362 37720 29368 37732
rect 29323 37692 29368 37720
rect 29362 37680 29368 37692
rect 29420 37680 29426 37732
rect 29454 37680 29460 37732
rect 29512 37720 29518 37732
rect 32674 37720 32680 37732
rect 29512 37692 29557 37720
rect 32635 37692 32680 37720
rect 29512 37680 29518 37692
rect 32674 37680 32680 37692
rect 32732 37680 32738 37732
rect 32769 37723 32827 37729
rect 32769 37689 32781 37723
rect 32815 37720 32827 37723
rect 33042 37720 33048 37732
rect 32815 37692 33048 37720
rect 32815 37689 32827 37692
rect 32769 37683 32827 37689
rect 33042 37680 33048 37692
rect 33100 37680 33106 37732
rect 35526 37680 35532 37732
rect 35584 37720 35590 37732
rect 35942 37723 36000 37729
rect 35942 37720 35954 37723
rect 35584 37692 35954 37720
rect 35584 37680 35590 37692
rect 35942 37689 35954 37692
rect 35988 37720 36000 37723
rect 36630 37720 36636 37732
rect 35988 37692 36636 37720
rect 35988 37689 36000 37692
rect 35942 37683 36000 37689
rect 36630 37680 36636 37692
rect 36688 37680 36694 37732
rect 37461 37723 37519 37729
rect 37461 37720 37473 37723
rect 36740 37692 37473 37720
rect 25547 37624 25820 37652
rect 29089 37655 29147 37661
rect 25547 37621 25559 37624
rect 25501 37615 25559 37621
rect 29089 37621 29101 37655
rect 29135 37652 29147 37655
rect 29472 37652 29500 37680
rect 29135 37624 29500 37652
rect 29135 37621 29147 37624
rect 29089 37615 29147 37621
rect 30558 37612 30564 37664
rect 30616 37652 30622 37664
rect 34701 37655 34759 37661
rect 34701 37652 34713 37655
rect 30616 37624 34713 37652
rect 30616 37612 30622 37624
rect 34701 37621 34713 37624
rect 34747 37652 34759 37655
rect 35250 37652 35256 37664
rect 34747 37624 35256 37652
rect 34747 37621 34759 37624
rect 34701 37615 34759 37621
rect 35250 37612 35256 37624
rect 35308 37652 35314 37664
rect 36538 37652 36544 37664
rect 35308 37624 36544 37652
rect 35308 37612 35314 37624
rect 36538 37612 36544 37624
rect 36596 37652 36602 37664
rect 36740 37652 36768 37692
rect 37461 37689 37473 37692
rect 37507 37720 37519 37723
rect 37734 37720 37740 37732
rect 37507 37692 37740 37720
rect 37507 37689 37519 37692
rect 37461 37683 37519 37689
rect 37734 37680 37740 37692
rect 37792 37680 37798 37732
rect 38749 37723 38807 37729
rect 38749 37689 38761 37723
rect 38795 37720 38807 37723
rect 38930 37720 38936 37732
rect 38795 37692 38936 37720
rect 38795 37689 38807 37692
rect 38749 37683 38807 37689
rect 38930 37680 38936 37692
rect 38988 37680 38994 37732
rect 39758 37680 39764 37732
rect 39816 37720 39822 37732
rect 40957 37723 41015 37729
rect 40957 37720 40969 37723
rect 39816 37692 40969 37720
rect 39816 37680 39822 37692
rect 40957 37689 40969 37692
rect 41003 37720 41015 37723
rect 41046 37720 41052 37732
rect 41003 37692 41052 37720
rect 41003 37689 41015 37692
rect 40957 37683 41015 37689
rect 41046 37680 41052 37692
rect 41104 37680 41110 37732
rect 41506 37720 41512 37732
rect 41467 37692 41512 37720
rect 41506 37680 41512 37692
rect 41564 37680 41570 37732
rect 42426 37720 42432 37732
rect 42387 37692 42432 37720
rect 42426 37680 42432 37692
rect 42484 37680 42490 37732
rect 42521 37723 42579 37729
rect 42521 37689 42533 37723
rect 42567 37689 42579 37723
rect 42521 37683 42579 37689
rect 43625 37723 43683 37729
rect 43625 37689 43637 37723
rect 43671 37720 43683 37723
rect 43901 37723 43959 37729
rect 43901 37720 43913 37723
rect 43671 37692 43913 37720
rect 43671 37689 43683 37692
rect 43625 37683 43683 37689
rect 43901 37689 43913 37692
rect 43947 37720 43959 37723
rect 44266 37720 44272 37732
rect 43947 37692 44272 37720
rect 43947 37689 43959 37692
rect 43901 37683 43959 37689
rect 36906 37652 36912 37664
rect 36596 37624 36768 37652
rect 36867 37624 36912 37652
rect 36596 37612 36602 37624
rect 36906 37612 36912 37624
rect 36964 37612 36970 37664
rect 39666 37652 39672 37664
rect 39627 37624 39672 37652
rect 39666 37612 39672 37624
rect 39724 37612 39730 37664
rect 41064 37652 41092 37680
rect 41785 37655 41843 37661
rect 41785 37652 41797 37655
rect 41064 37624 41797 37652
rect 41785 37621 41797 37624
rect 41831 37652 41843 37655
rect 41874 37652 41880 37664
rect 41831 37624 41880 37652
rect 41831 37621 41843 37624
rect 41785 37615 41843 37621
rect 41874 37612 41880 37624
rect 41932 37652 41938 37664
rect 42153 37655 42211 37661
rect 42153 37652 42165 37655
rect 41932 37624 42165 37652
rect 41932 37612 41938 37624
rect 42153 37621 42165 37624
rect 42199 37652 42211 37655
rect 42536 37652 42564 37683
rect 44266 37680 44272 37692
rect 44324 37680 44330 37732
rect 42199 37624 42564 37652
rect 42199 37621 42211 37624
rect 42153 37615 42211 37621
rect 43990 37612 43996 37664
rect 44048 37652 44054 37664
rect 46247 37655 46305 37661
rect 46247 37652 46259 37655
rect 44048 37624 46259 37652
rect 44048 37612 44054 37624
rect 46247 37621 46259 37624
rect 46293 37621 46305 37655
rect 46247 37615 46305 37621
rect 1104 37562 48852 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 48852 37562
rect 1104 37488 48852 37510
rect 15562 37448 15568 37460
rect 15523 37420 15568 37448
rect 15562 37408 15568 37420
rect 15620 37408 15626 37460
rect 18414 37408 18420 37460
rect 18472 37448 18478 37460
rect 18693 37451 18751 37457
rect 18693 37448 18705 37451
rect 18472 37420 18705 37448
rect 18472 37408 18478 37420
rect 18693 37417 18705 37420
rect 18739 37417 18751 37451
rect 18693 37411 18751 37417
rect 20898 37408 20904 37460
rect 20956 37448 20962 37460
rect 23658 37448 23664 37460
rect 20956 37420 22784 37448
rect 20956 37408 20962 37420
rect 15286 37340 15292 37392
rect 15344 37380 15350 37392
rect 16025 37383 16083 37389
rect 16025 37380 16037 37383
rect 15344 37352 16037 37380
rect 15344 37340 15350 37352
rect 16025 37349 16037 37352
rect 16071 37349 16083 37383
rect 16025 37343 16083 37349
rect 16114 37340 16120 37392
rect 16172 37380 16178 37392
rect 16945 37383 17003 37389
rect 16945 37380 16957 37383
rect 16172 37352 16957 37380
rect 16172 37340 16178 37352
rect 16945 37349 16957 37352
rect 16991 37349 17003 37383
rect 17770 37380 17776 37392
rect 17731 37352 17776 37380
rect 16945 37343 17003 37349
rect 17770 37340 17776 37352
rect 17828 37340 17834 37392
rect 17865 37383 17923 37389
rect 17865 37349 17877 37383
rect 17911 37380 17923 37383
rect 17954 37380 17960 37392
rect 17911 37352 17960 37380
rect 17911 37349 17923 37352
rect 17865 37343 17923 37349
rect 17954 37340 17960 37352
rect 18012 37340 18018 37392
rect 19426 37380 19432 37392
rect 19339 37352 19432 37380
rect 19426 37340 19432 37352
rect 19484 37380 19490 37392
rect 21085 37383 21143 37389
rect 21085 37380 21097 37383
rect 19484 37352 21097 37380
rect 19484 37340 19490 37352
rect 21085 37349 21097 37352
rect 21131 37380 21143 37383
rect 21726 37380 21732 37392
rect 21131 37352 21732 37380
rect 21131 37349 21143 37352
rect 21085 37343 21143 37349
rect 21726 37340 21732 37352
rect 21784 37340 21790 37392
rect 22756 37324 22784 37420
rect 23492 37420 23664 37448
rect 23492 37389 23520 37420
rect 23658 37408 23664 37420
rect 23716 37448 23722 37460
rect 23753 37451 23811 37457
rect 23753 37448 23765 37451
rect 23716 37420 23765 37448
rect 23716 37408 23722 37420
rect 23753 37417 23765 37420
rect 23799 37417 23811 37451
rect 24946 37448 24952 37460
rect 24907 37420 24952 37448
rect 23753 37411 23811 37417
rect 24946 37408 24952 37420
rect 25004 37408 25010 37460
rect 27709 37451 27767 37457
rect 27709 37417 27721 37451
rect 27755 37448 27767 37451
rect 28166 37448 28172 37460
rect 27755 37420 28172 37448
rect 27755 37417 27767 37420
rect 27709 37411 27767 37417
rect 28166 37408 28172 37420
rect 28224 37408 28230 37460
rect 28534 37408 28540 37460
rect 28592 37448 28598 37460
rect 29181 37451 29239 37457
rect 29181 37448 29193 37451
rect 28592 37420 29193 37448
rect 28592 37408 28598 37420
rect 29181 37417 29193 37420
rect 29227 37417 29239 37451
rect 29181 37411 29239 37417
rect 29270 37408 29276 37460
rect 29328 37448 29334 37460
rect 30929 37451 30987 37457
rect 30929 37448 30941 37451
rect 29328 37420 30941 37448
rect 29328 37408 29334 37420
rect 30929 37417 30941 37420
rect 30975 37448 30987 37451
rect 31294 37448 31300 37460
rect 30975 37420 31300 37448
rect 30975 37417 30987 37420
rect 30929 37411 30987 37417
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 32769 37451 32827 37457
rect 32769 37417 32781 37451
rect 32815 37448 32827 37451
rect 33042 37448 33048 37460
rect 32815 37420 33048 37448
rect 32815 37417 32827 37420
rect 32769 37411 32827 37417
rect 33042 37408 33048 37420
rect 33100 37408 33106 37460
rect 33612 37420 37780 37448
rect 23477 37383 23535 37389
rect 23477 37349 23489 37383
rect 23523 37349 23535 37383
rect 23477 37343 23535 37349
rect 28353 37383 28411 37389
rect 28353 37349 28365 37383
rect 28399 37380 28411 37383
rect 28442 37380 28448 37392
rect 28399 37352 28448 37380
rect 28399 37349 28411 37352
rect 28353 37343 28411 37349
rect 28442 37340 28448 37352
rect 28500 37340 28506 37392
rect 33612 37380 33640 37420
rect 29840 37352 33640 37380
rect 33689 37383 33747 37389
rect 29840 37324 29868 37352
rect 33689 37349 33701 37383
rect 33735 37380 33747 37383
rect 33778 37380 33784 37392
rect 33735 37352 33784 37380
rect 33735 37349 33747 37352
rect 33689 37343 33747 37349
rect 33778 37340 33784 37352
rect 33836 37340 33842 37392
rect 35805 37383 35863 37389
rect 35805 37349 35817 37383
rect 35851 37380 35863 37383
rect 35986 37380 35992 37392
rect 35851 37352 35992 37380
rect 35851 37349 35863 37352
rect 35805 37343 35863 37349
rect 35986 37340 35992 37352
rect 36044 37340 36050 37392
rect 13998 37272 14004 37324
rect 14056 37312 14062 37324
rect 14220 37315 14278 37321
rect 14220 37312 14232 37315
rect 14056 37284 14232 37312
rect 14056 37272 14062 37284
rect 14220 37281 14232 37284
rect 14266 37281 14278 37315
rect 22738 37312 22744 37324
rect 22651 37284 22744 37312
rect 14220 37275 14278 37281
rect 22738 37272 22744 37284
rect 22796 37272 22802 37324
rect 23198 37312 23204 37324
rect 23159 37284 23204 37312
rect 23198 37272 23204 37284
rect 23256 37272 23262 37324
rect 24356 37315 24414 37321
rect 24356 37281 24368 37315
rect 24402 37312 24414 37315
rect 24670 37312 24676 37324
rect 24402 37284 24676 37312
rect 24402 37281 24414 37284
rect 24356 37275 24414 37281
rect 24670 37272 24676 37284
rect 24728 37272 24734 37324
rect 25314 37312 25320 37324
rect 25275 37284 25320 37312
rect 25314 37272 25320 37284
rect 25372 37272 25378 37324
rect 26580 37315 26638 37321
rect 26580 37281 26592 37315
rect 26626 37312 26638 37315
rect 26786 37312 26792 37324
rect 26626 37284 26792 37312
rect 26626 37281 26638 37284
rect 26580 37275 26638 37281
rect 26786 37272 26792 37284
rect 26844 37272 26850 37324
rect 29822 37312 29828 37324
rect 29783 37284 29828 37312
rect 29822 37272 29828 37284
rect 29880 37272 29886 37324
rect 31018 37312 31024 37324
rect 30979 37284 31024 37312
rect 31018 37272 31024 37284
rect 31076 37272 31082 37324
rect 35342 37312 35348 37324
rect 35303 37284 35348 37312
rect 35342 37272 35348 37284
rect 35400 37272 35406 37324
rect 35434 37272 35440 37324
rect 35492 37312 35498 37324
rect 35529 37315 35587 37321
rect 35529 37312 35541 37315
rect 35492 37284 35541 37312
rect 35492 37272 35498 37284
rect 35529 37281 35541 37284
rect 35575 37281 35587 37315
rect 35529 37275 35587 37281
rect 36262 37272 36268 37324
rect 36320 37312 36326 37324
rect 37752 37321 37780 37420
rect 39114 37408 39120 37460
rect 39172 37448 39178 37460
rect 39209 37451 39267 37457
rect 39209 37448 39221 37451
rect 39172 37420 39221 37448
rect 39172 37408 39178 37420
rect 39209 37417 39221 37420
rect 39255 37417 39267 37451
rect 39758 37448 39764 37460
rect 39719 37420 39764 37448
rect 39209 37411 39267 37417
rect 39758 37408 39764 37420
rect 39816 37408 39822 37460
rect 41782 37448 41788 37460
rect 41743 37420 41788 37448
rect 41782 37408 41788 37420
rect 41840 37408 41846 37460
rect 42426 37448 42432 37460
rect 42387 37420 42432 37448
rect 42426 37408 42432 37420
rect 42484 37408 42490 37460
rect 43990 37448 43996 37460
rect 43951 37420 43996 37448
rect 43990 37408 43996 37420
rect 44048 37408 44054 37460
rect 40678 37340 40684 37392
rect 40736 37380 40742 37392
rect 40910 37383 40968 37389
rect 40910 37380 40922 37383
rect 40736 37352 40922 37380
rect 40736 37340 40742 37352
rect 40910 37349 40922 37352
rect 40956 37349 40968 37383
rect 40910 37343 40968 37349
rect 44453 37383 44511 37389
rect 44453 37349 44465 37383
rect 44499 37380 44511 37383
rect 45094 37380 45100 37392
rect 44499 37352 45100 37380
rect 44499 37349 44511 37352
rect 44453 37343 44511 37349
rect 45094 37340 45100 37352
rect 45152 37380 45158 37392
rect 46017 37383 46075 37389
rect 46017 37380 46029 37383
rect 45152 37352 46029 37380
rect 45152 37340 45158 37352
rect 46017 37349 46029 37352
rect 46063 37349 46075 37383
rect 46017 37343 46075 37349
rect 36633 37315 36691 37321
rect 36633 37312 36645 37315
rect 36320 37284 36645 37312
rect 36320 37272 36326 37284
rect 36633 37281 36645 37284
rect 36679 37281 36691 37315
rect 36633 37275 36691 37281
rect 37737 37315 37795 37321
rect 37737 37281 37749 37315
rect 37783 37312 37795 37315
rect 37826 37312 37832 37324
rect 37783 37284 37832 37312
rect 37783 37281 37795 37284
rect 37737 37275 37795 37281
rect 37826 37272 37832 37284
rect 37884 37272 37890 37324
rect 19334 37244 19340 37256
rect 19295 37216 19340 37244
rect 19334 37204 19340 37216
rect 19392 37204 19398 37256
rect 19610 37244 19616 37256
rect 19571 37216 19616 37244
rect 19610 37204 19616 37216
rect 19668 37204 19674 37256
rect 20990 37244 20996 37256
rect 20951 37216 20996 37244
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 21358 37244 21364 37256
rect 21319 37216 21364 37244
rect 21358 37204 21364 37216
rect 21416 37204 21422 37256
rect 24443 37247 24501 37253
rect 24443 37213 24455 37247
rect 24489 37244 24501 37247
rect 25682 37244 25688 37256
rect 24489 37216 25688 37244
rect 24489 37213 24501 37216
rect 24443 37207 24501 37213
rect 25682 37204 25688 37216
rect 25740 37244 25746 37256
rect 25777 37247 25835 37253
rect 25777 37244 25789 37247
rect 25740 37216 25789 37244
rect 25740 37204 25746 37216
rect 25777 37213 25789 37216
rect 25823 37213 25835 37247
rect 25777 37207 25835 37213
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 28261 37247 28319 37253
rect 28261 37244 28273 37247
rect 27764 37216 28273 37244
rect 27764 37204 27770 37216
rect 28261 37213 28273 37216
rect 28307 37213 28319 37247
rect 28261 37207 28319 37213
rect 28350 37204 28356 37256
rect 28408 37244 28414 37256
rect 28537 37247 28595 37253
rect 28537 37244 28549 37247
rect 28408 37216 28549 37244
rect 28408 37204 28414 37216
rect 28537 37213 28549 37216
rect 28583 37213 28595 37247
rect 32214 37244 32220 37256
rect 32175 37216 32220 37244
rect 28537 37207 28595 37213
rect 32214 37204 32220 37216
rect 32272 37204 32278 37256
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 34241 37247 34299 37253
rect 34241 37213 34253 37247
rect 34287 37244 34299 37247
rect 34330 37244 34336 37256
rect 34287 37216 34336 37244
rect 34287 37213 34299 37216
rect 34241 37207 34299 37213
rect 16390 37136 16396 37188
rect 16448 37176 16454 37188
rect 16577 37179 16635 37185
rect 16577 37176 16589 37179
rect 16448 37148 16589 37176
rect 16448 37136 16454 37148
rect 16577 37145 16589 37148
rect 16623 37176 16635 37179
rect 18325 37179 18383 37185
rect 18325 37176 18337 37179
rect 16623 37148 18337 37176
rect 16623 37145 16635 37148
rect 16577 37139 16635 37145
rect 18325 37145 18337 37148
rect 18371 37176 18383 37179
rect 19886 37176 19892 37188
rect 18371 37148 19892 37176
rect 18371 37145 18383 37148
rect 18325 37139 18383 37145
rect 19886 37136 19892 37148
rect 19944 37136 19950 37188
rect 25222 37136 25228 37188
rect 25280 37176 25286 37188
rect 26651 37179 26709 37185
rect 26651 37176 26663 37179
rect 25280 37148 26663 37176
rect 25280 37136 25286 37148
rect 26651 37145 26663 37148
rect 26697 37145 26709 37179
rect 26651 37139 26709 37145
rect 31110 37136 31116 37188
rect 31168 37176 31174 37188
rect 31168 37148 32489 37176
rect 31168 37136 31174 37148
rect 32461 37120 32489 37148
rect 32674 37136 32680 37188
rect 32732 37176 32738 37188
rect 33137 37179 33195 37185
rect 33137 37176 33149 37179
rect 32732 37148 33149 37176
rect 32732 37136 32738 37148
rect 33137 37145 33149 37148
rect 33183 37176 33195 37179
rect 34256 37176 34284 37207
rect 34330 37204 34336 37216
rect 34388 37204 34394 37256
rect 38841 37247 38899 37253
rect 38841 37213 38853 37247
rect 38887 37244 38899 37247
rect 38930 37244 38936 37256
rect 38887 37216 38936 37244
rect 38887 37213 38899 37216
rect 38841 37207 38899 37213
rect 38930 37204 38936 37216
rect 38988 37204 38994 37256
rect 40586 37244 40592 37256
rect 40547 37216 40592 37244
rect 40586 37204 40592 37216
rect 40644 37204 40650 37256
rect 44358 37244 44364 37256
rect 44319 37216 44364 37244
rect 44358 37204 44364 37216
rect 44416 37204 44422 37256
rect 44726 37244 44732 37256
rect 44687 37216 44732 37244
rect 44726 37204 44732 37216
rect 44784 37204 44790 37256
rect 45922 37244 45928 37256
rect 45883 37216 45928 37244
rect 45922 37204 45928 37216
rect 45980 37204 45986 37256
rect 46198 37244 46204 37256
rect 46159 37216 46204 37244
rect 46198 37204 46204 37216
rect 46256 37204 46262 37256
rect 33183 37148 34284 37176
rect 33183 37145 33195 37148
rect 33137 37139 33195 37145
rect 41046 37136 41052 37188
rect 41104 37176 41110 37188
rect 41509 37179 41567 37185
rect 41509 37176 41521 37179
rect 41104 37148 41521 37176
rect 41104 37136 41110 37148
rect 41509 37145 41521 37148
rect 41555 37176 41567 37179
rect 44266 37176 44272 37188
rect 41555 37148 44272 37176
rect 41555 37145 41567 37148
rect 41509 37139 41567 37145
rect 44266 37136 44272 37148
rect 44324 37136 44330 37188
rect 14323 37111 14381 37117
rect 14323 37077 14335 37111
rect 14369 37108 14381 37111
rect 15378 37108 15384 37120
rect 14369 37080 15384 37108
rect 14369 37077 14381 37080
rect 14323 37071 14381 37077
rect 15378 37068 15384 37080
rect 15436 37068 15442 37120
rect 16022 37068 16028 37120
rect 16080 37108 16086 37120
rect 21818 37108 21824 37120
rect 16080 37080 21824 37108
rect 16080 37068 16086 37080
rect 21818 37068 21824 37080
rect 21876 37068 21882 37120
rect 22002 37108 22008 37120
rect 21963 37080 22008 37108
rect 22002 37068 22008 37080
rect 22060 37068 22066 37120
rect 24118 37108 24124 37120
rect 24079 37080 24124 37108
rect 24118 37068 24124 37080
rect 24176 37068 24182 37120
rect 25455 37111 25513 37117
rect 25455 37077 25467 37111
rect 25501 37108 25513 37111
rect 26326 37108 26332 37120
rect 25501 37080 26332 37108
rect 25501 37077 25513 37080
rect 25455 37071 25513 37077
rect 26326 37068 26332 37080
rect 26384 37068 26390 37120
rect 29362 37068 29368 37120
rect 29420 37108 29426 37120
rect 29549 37111 29607 37117
rect 29549 37108 29561 37111
rect 29420 37080 29561 37108
rect 29420 37068 29426 37080
rect 29549 37077 29561 37080
rect 29595 37077 29607 37111
rect 29549 37071 29607 37077
rect 30055 37111 30113 37117
rect 30055 37077 30067 37111
rect 30101 37108 30113 37111
rect 30282 37108 30288 37120
rect 30101 37080 30288 37108
rect 30101 37077 30113 37080
rect 30055 37071 30113 37077
rect 30282 37068 30288 37080
rect 30340 37068 30346 37120
rect 30466 37108 30472 37120
rect 30427 37080 30472 37108
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 31205 37111 31263 37117
rect 31205 37077 31217 37111
rect 31251 37108 31263 37111
rect 31294 37108 31300 37120
rect 31251 37080 31300 37108
rect 31251 37077 31263 37080
rect 31205 37071 31263 37077
rect 31294 37068 31300 37080
rect 31352 37068 31358 37120
rect 32398 37108 32404 37120
rect 32356 37080 32404 37108
rect 32398 37068 32404 37080
rect 32456 37108 32489 37120
rect 36817 37111 36875 37117
rect 36817 37108 36829 37111
rect 32456 37080 36829 37108
rect 32456 37068 32462 37080
rect 36817 37077 36829 37080
rect 36863 37077 36875 37111
rect 37090 37108 37096 37120
rect 37051 37080 37096 37108
rect 36817 37071 36875 37077
rect 37090 37068 37096 37080
rect 37148 37068 37154 37120
rect 37967 37111 38025 37117
rect 37967 37077 37979 37111
rect 38013 37108 38025 37111
rect 38194 37108 38200 37120
rect 38013 37080 38200 37108
rect 38013 37077 38025 37080
rect 37967 37071 38025 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 38381 37111 38439 37117
rect 38381 37077 38393 37111
rect 38427 37108 38439 37111
rect 38470 37108 38476 37120
rect 38427 37080 38476 37108
rect 38427 37077 38439 37080
rect 38381 37071 38439 37077
rect 38470 37068 38476 37080
rect 38528 37108 38534 37120
rect 39022 37108 39028 37120
rect 38528 37080 39028 37108
rect 38528 37068 38534 37080
rect 39022 37068 39028 37080
rect 39080 37068 39086 37120
rect 43898 37068 43904 37120
rect 43956 37108 43962 37120
rect 45738 37108 45744 37120
rect 43956 37080 45744 37108
rect 43956 37068 43962 37080
rect 45738 37068 45744 37080
rect 45796 37068 45802 37120
rect 1104 37018 48852 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 48852 37018
rect 1104 36944 48852 36966
rect 15473 36907 15531 36913
rect 15473 36873 15485 36907
rect 15519 36904 15531 36907
rect 16025 36907 16083 36913
rect 16025 36904 16037 36907
rect 15519 36876 16037 36904
rect 15519 36873 15531 36876
rect 15473 36867 15531 36873
rect 16025 36873 16037 36876
rect 16071 36904 16083 36907
rect 16114 36904 16120 36916
rect 16071 36876 16120 36904
rect 16071 36873 16083 36876
rect 16025 36867 16083 36873
rect 16114 36864 16120 36876
rect 16172 36864 16178 36916
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19705 36907 19763 36913
rect 19705 36904 19717 36907
rect 19392 36876 19717 36904
rect 19392 36864 19398 36876
rect 19705 36873 19717 36876
rect 19751 36873 19763 36907
rect 19705 36867 19763 36873
rect 20165 36907 20223 36913
rect 20165 36873 20177 36907
rect 20211 36904 20223 36907
rect 20990 36904 20996 36916
rect 20211 36876 20996 36904
rect 20211 36873 20223 36876
rect 20165 36867 20223 36873
rect 20990 36864 20996 36876
rect 21048 36904 21054 36916
rect 22327 36907 22385 36913
rect 22327 36904 22339 36907
rect 21048 36876 22339 36904
rect 21048 36864 21054 36876
rect 22327 36873 22339 36876
rect 22373 36873 22385 36907
rect 22327 36867 22385 36873
rect 22738 36864 22744 36916
rect 22796 36904 22802 36916
rect 23385 36907 23443 36913
rect 23385 36904 23397 36907
rect 22796 36876 23397 36904
rect 22796 36864 22802 36876
rect 23385 36873 23397 36876
rect 23431 36873 23443 36907
rect 24670 36904 24676 36916
rect 24631 36876 24676 36904
rect 23385 36867 23443 36873
rect 24670 36864 24676 36876
rect 24728 36864 24734 36916
rect 25314 36904 25320 36916
rect 25275 36876 25320 36904
rect 25314 36864 25320 36876
rect 25372 36864 25378 36916
rect 26786 36904 26792 36916
rect 26747 36876 26792 36904
rect 26786 36864 26792 36876
rect 26844 36864 26850 36916
rect 28074 36864 28080 36916
rect 28132 36904 28138 36916
rect 28353 36907 28411 36913
rect 28353 36904 28365 36907
rect 28132 36876 28365 36904
rect 28132 36864 28138 36876
rect 28353 36873 28365 36876
rect 28399 36873 28411 36907
rect 28353 36867 28411 36873
rect 29822 36864 29828 36916
rect 29880 36904 29886 36916
rect 30653 36907 30711 36913
rect 30653 36904 30665 36907
rect 29880 36876 30665 36904
rect 29880 36864 29886 36876
rect 30653 36873 30665 36876
rect 30699 36873 30711 36907
rect 32214 36904 32220 36916
rect 32175 36876 32220 36904
rect 30653 36867 30711 36873
rect 32214 36864 32220 36876
rect 32272 36864 32278 36916
rect 35161 36907 35219 36913
rect 35161 36873 35173 36907
rect 35207 36904 35219 36907
rect 35434 36904 35440 36916
rect 35207 36876 35440 36904
rect 35207 36873 35219 36876
rect 35161 36867 35219 36873
rect 35434 36864 35440 36876
rect 35492 36904 35498 36916
rect 35805 36907 35863 36913
rect 35805 36904 35817 36907
rect 35492 36876 35817 36904
rect 35492 36864 35498 36876
rect 35805 36873 35817 36876
rect 35851 36873 35863 36907
rect 36630 36904 36636 36916
rect 36591 36876 36636 36904
rect 35805 36867 35863 36873
rect 36630 36864 36636 36876
rect 36688 36864 36694 36916
rect 37737 36907 37795 36913
rect 37737 36873 37749 36907
rect 37783 36904 37795 36907
rect 41138 36904 41144 36916
rect 37783 36876 41144 36904
rect 37783 36873 37795 36876
rect 37737 36867 37795 36873
rect 41138 36864 41144 36876
rect 41196 36864 41202 36916
rect 42426 36864 42432 36916
rect 42484 36904 42490 36916
rect 42567 36907 42625 36913
rect 42567 36904 42579 36907
rect 42484 36876 42579 36904
rect 42484 36864 42490 36876
rect 42567 36873 42579 36876
rect 42613 36873 42625 36907
rect 42567 36867 42625 36873
rect 43349 36907 43407 36913
rect 43349 36873 43361 36907
rect 43395 36904 43407 36907
rect 43579 36907 43637 36913
rect 43579 36904 43591 36907
rect 43395 36876 43591 36904
rect 43395 36873 43407 36876
rect 43349 36867 43407 36873
rect 43579 36873 43591 36876
rect 43625 36904 43637 36907
rect 44358 36904 44364 36916
rect 43625 36876 44364 36904
rect 43625 36873 43637 36876
rect 43579 36867 43637 36873
rect 44358 36864 44364 36876
rect 44416 36864 44422 36916
rect 16945 36839 17003 36845
rect 16945 36805 16957 36839
rect 16991 36836 17003 36839
rect 17678 36836 17684 36848
rect 16991 36808 17684 36836
rect 16991 36805 17003 36808
rect 16945 36799 17003 36805
rect 17678 36796 17684 36808
rect 17736 36836 17742 36848
rect 19426 36836 19432 36848
rect 17736 36808 19104 36836
rect 19387 36808 19432 36836
rect 17736 36796 17742 36808
rect 15378 36728 15384 36780
rect 15436 36768 15442 36780
rect 16393 36771 16451 36777
rect 16393 36768 16405 36771
rect 15436 36740 16405 36768
rect 15436 36728 15442 36740
rect 16393 36737 16405 36740
rect 16439 36768 16451 36771
rect 16666 36768 16672 36780
rect 16439 36740 16672 36768
rect 16439 36737 16451 36740
rect 16393 36731 16451 36737
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 18414 36768 18420 36780
rect 18375 36740 18420 36768
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 19076 36777 19104 36808
rect 19426 36796 19432 36808
rect 19484 36796 19490 36848
rect 21818 36796 21824 36848
rect 21876 36836 21882 36848
rect 23017 36839 23075 36845
rect 23017 36836 23029 36839
rect 21876 36808 23029 36836
rect 21876 36796 21882 36808
rect 23017 36805 23029 36808
rect 23063 36836 23075 36839
rect 23198 36836 23204 36848
rect 23063 36808 23204 36836
rect 23063 36805 23075 36808
rect 23017 36799 23075 36805
rect 23198 36796 23204 36808
rect 23256 36796 23262 36848
rect 24486 36796 24492 36848
rect 24544 36836 24550 36848
rect 24544 36808 30788 36836
rect 24544 36796 24550 36808
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36768 19119 36771
rect 19610 36768 19616 36780
rect 19107 36740 19616 36768
rect 19107 36737 19119 36740
rect 19061 36731 19119 36737
rect 19610 36728 19616 36740
rect 19668 36768 19674 36780
rect 19886 36768 19892 36780
rect 19668 36740 19892 36768
rect 19668 36728 19674 36740
rect 19886 36728 19892 36740
rect 19944 36728 19950 36780
rect 20714 36768 20720 36780
rect 20675 36740 20720 36768
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 23753 36771 23811 36777
rect 23753 36737 23765 36771
rect 23799 36768 23811 36771
rect 24118 36768 24124 36780
rect 23799 36740 24124 36768
rect 23799 36737 23811 36740
rect 23753 36731 23811 36737
rect 24118 36728 24124 36740
rect 24176 36728 24182 36780
rect 24210 36728 24216 36780
rect 24268 36768 24274 36780
rect 25869 36771 25927 36777
rect 24268 36740 24313 36768
rect 24268 36728 24274 36740
rect 25869 36737 25881 36771
rect 25915 36768 25927 36771
rect 26142 36768 26148 36780
rect 25915 36740 26148 36768
rect 25915 36737 25927 36740
rect 25869 36731 25927 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 26234 36728 26240 36780
rect 26292 36768 26298 36780
rect 26292 36740 26337 36768
rect 26292 36728 26298 36740
rect 26878 36728 26884 36780
rect 26936 36768 26942 36780
rect 30009 36771 30067 36777
rect 30009 36768 30021 36771
rect 26936 36740 30021 36768
rect 26936 36728 26942 36740
rect 30009 36737 30021 36740
rect 30055 36768 30067 36771
rect 30466 36768 30472 36780
rect 30055 36740 30472 36768
rect 30055 36737 30067 36740
rect 30009 36731 30067 36737
rect 30466 36728 30472 36740
rect 30524 36728 30530 36780
rect 14550 36700 14556 36712
rect 14511 36672 14556 36700
rect 14550 36660 14556 36672
rect 14608 36660 14614 36712
rect 22256 36703 22314 36709
rect 22256 36669 22268 36703
rect 22302 36700 22314 36703
rect 22646 36700 22652 36712
rect 22302 36672 22652 36700
rect 22302 36669 22314 36672
rect 22256 36663 22314 36669
rect 22646 36660 22652 36672
rect 22704 36660 22710 36712
rect 27960 36703 28018 36709
rect 27960 36669 27972 36703
rect 28006 36700 28018 36703
rect 28074 36700 28080 36712
rect 28006 36672 28080 36700
rect 28006 36669 28018 36672
rect 27960 36663 28018 36669
rect 28074 36660 28080 36672
rect 28132 36660 28138 36712
rect 30760 36700 30788 36808
rect 32232 36768 32260 36864
rect 34146 36796 34152 36848
rect 34204 36836 34210 36848
rect 34701 36839 34759 36845
rect 34701 36836 34713 36839
rect 34204 36808 34713 36836
rect 34204 36796 34210 36808
rect 34701 36805 34713 36808
rect 34747 36836 34759 36839
rect 35342 36836 35348 36848
rect 34747 36808 35348 36836
rect 34747 36805 34759 36808
rect 34701 36799 34759 36805
rect 35342 36796 35348 36808
rect 35400 36796 35406 36848
rect 37826 36796 37832 36848
rect 37884 36836 37890 36848
rect 38013 36839 38071 36845
rect 38013 36836 38025 36839
rect 37884 36808 38025 36836
rect 37884 36796 37890 36808
rect 38013 36805 38025 36808
rect 38059 36805 38071 36839
rect 38013 36799 38071 36805
rect 39114 36796 39120 36848
rect 39172 36836 39178 36848
rect 39577 36839 39635 36845
rect 39577 36836 39589 36839
rect 39172 36808 39589 36836
rect 39172 36796 39178 36808
rect 39577 36805 39589 36808
rect 39623 36836 39635 36839
rect 40129 36839 40187 36845
rect 40129 36836 40141 36839
rect 39623 36808 40141 36836
rect 39623 36805 39635 36808
rect 39577 36799 39635 36805
rect 40129 36805 40141 36808
rect 40175 36805 40187 36839
rect 40129 36799 40187 36805
rect 40313 36839 40371 36845
rect 40313 36805 40325 36839
rect 40359 36836 40371 36839
rect 41046 36836 41052 36848
rect 40359 36808 41052 36836
rect 40359 36805 40371 36808
rect 40313 36799 40371 36805
rect 41046 36796 41052 36808
rect 41104 36796 41110 36848
rect 41506 36836 41512 36848
rect 41467 36808 41512 36836
rect 41506 36796 41512 36808
rect 41564 36796 41570 36848
rect 45094 36796 45100 36848
rect 45152 36836 45158 36848
rect 45833 36839 45891 36845
rect 45833 36836 45845 36839
rect 45152 36808 45845 36836
rect 45152 36796 45158 36808
rect 45833 36805 45845 36808
rect 45879 36805 45891 36839
rect 45833 36799 45891 36805
rect 32401 36771 32459 36777
rect 32401 36768 32413 36771
rect 32232 36740 32413 36768
rect 32401 36737 32413 36740
rect 32447 36737 32459 36771
rect 32674 36768 32680 36780
rect 32635 36740 32680 36768
rect 32401 36731 32459 36737
rect 32674 36728 32680 36740
rect 32732 36728 32738 36780
rect 36817 36771 36875 36777
rect 36817 36737 36829 36771
rect 36863 36768 36875 36771
rect 37090 36768 37096 36780
rect 36863 36740 37096 36768
rect 36863 36737 36875 36740
rect 36817 36731 36875 36737
rect 37090 36728 37096 36740
rect 37148 36728 37154 36780
rect 38194 36728 38200 36780
rect 38252 36768 38258 36780
rect 40957 36771 41015 36777
rect 40957 36768 40969 36771
rect 38252 36740 40969 36768
rect 38252 36728 38258 36740
rect 40957 36737 40969 36740
rect 41003 36768 41015 36771
rect 41877 36771 41935 36777
rect 41877 36768 41889 36771
rect 41003 36740 41889 36768
rect 41003 36737 41015 36740
rect 40957 36731 41015 36737
rect 41877 36737 41889 36740
rect 41923 36737 41935 36771
rect 41877 36731 41935 36737
rect 42334 36728 42340 36780
rect 42392 36768 42398 36780
rect 44361 36771 44419 36777
rect 42392 36740 43551 36768
rect 42392 36728 42398 36740
rect 31348 36703 31406 36709
rect 31348 36700 31360 36703
rect 30760 36672 31360 36700
rect 31348 36669 31360 36672
rect 31394 36700 31406 36703
rect 34977 36703 35035 36709
rect 31394 36669 31407 36700
rect 31348 36663 31407 36669
rect 34977 36669 34989 36703
rect 35023 36700 35035 36703
rect 38562 36700 38568 36712
rect 35023 36672 35572 36700
rect 35023 36669 35035 36672
rect 34977 36663 35035 36669
rect 14461 36635 14519 36641
rect 14461 36601 14473 36635
rect 14507 36632 14519 36635
rect 14642 36632 14648 36644
rect 14507 36604 14648 36632
rect 14507 36601 14519 36604
rect 14461 36595 14519 36601
rect 14642 36592 14648 36604
rect 14700 36632 14706 36644
rect 14874 36635 14932 36641
rect 14874 36632 14886 36635
rect 14700 36604 14886 36632
rect 14700 36592 14706 36604
rect 14874 36601 14886 36604
rect 14920 36601 14932 36635
rect 14874 36595 14932 36601
rect 16485 36635 16543 36641
rect 16485 36601 16497 36635
rect 16531 36601 16543 36635
rect 16485 36595 16543 36601
rect 17497 36635 17555 36641
rect 17497 36601 17509 36635
rect 17543 36632 17555 36635
rect 17865 36635 17923 36641
rect 17865 36632 17877 36635
rect 17543 36604 17877 36632
rect 17543 36601 17555 36604
rect 17497 36595 17555 36601
rect 17865 36601 17877 36604
rect 17911 36632 17923 36635
rect 17954 36632 17960 36644
rect 17911 36604 17960 36632
rect 17911 36601 17923 36604
rect 17865 36595 17923 36601
rect 13998 36564 14004 36576
rect 13959 36536 14004 36564
rect 13998 36524 14004 36536
rect 14056 36524 14062 36576
rect 16114 36524 16120 36576
rect 16172 36564 16178 36576
rect 16500 36564 16528 36595
rect 17954 36592 17960 36604
rect 18012 36632 18018 36644
rect 18509 36635 18567 36641
rect 18509 36632 18521 36635
rect 18012 36604 18521 36632
rect 18012 36592 18018 36604
rect 18509 36601 18521 36604
rect 18555 36632 18567 36635
rect 20533 36635 20591 36641
rect 20533 36632 20545 36635
rect 18555 36604 20545 36632
rect 18555 36601 18567 36604
rect 18509 36595 18567 36601
rect 20533 36601 20545 36604
rect 20579 36632 20591 36635
rect 20806 36632 20812 36644
rect 20579 36604 20812 36632
rect 20579 36601 20591 36604
rect 20533 36595 20591 36601
rect 20806 36592 20812 36604
rect 20864 36592 20870 36644
rect 21358 36632 21364 36644
rect 21271 36604 21364 36632
rect 21358 36592 21364 36604
rect 21416 36592 21422 36644
rect 21726 36632 21732 36644
rect 21639 36604 21732 36632
rect 21726 36592 21732 36604
rect 21784 36632 21790 36644
rect 23845 36635 23903 36641
rect 23845 36632 23857 36635
rect 21784 36604 23857 36632
rect 21784 36592 21790 36604
rect 23845 36601 23857 36604
rect 23891 36632 23903 36635
rect 23934 36632 23940 36644
rect 23891 36604 23940 36632
rect 23891 36601 23903 36604
rect 23845 36595 23903 36601
rect 23934 36592 23940 36604
rect 23992 36592 23998 36644
rect 25958 36632 25964 36644
rect 25919 36604 25964 36632
rect 25958 36592 25964 36604
rect 26016 36592 26022 36644
rect 29730 36632 29736 36644
rect 29691 36604 29736 36632
rect 29730 36592 29736 36604
rect 29788 36592 29794 36644
rect 29825 36635 29883 36641
rect 29825 36601 29837 36635
rect 29871 36632 29883 36635
rect 30926 36632 30932 36644
rect 29871 36604 30932 36632
rect 29871 36601 29883 36604
rect 29825 36595 29883 36601
rect 16172 36536 16528 36564
rect 16172 36524 16178 36536
rect 16574 36524 16580 36576
rect 16632 36564 16638 36576
rect 21376 36564 21404 36592
rect 22646 36564 22652 36576
rect 16632 36536 21404 36564
rect 22607 36536 22652 36564
rect 16632 36524 16638 36536
rect 22646 36524 22652 36536
rect 22704 36524 22710 36576
rect 27706 36564 27712 36576
rect 27667 36536 27712 36564
rect 27706 36524 27712 36536
rect 27764 36524 27770 36576
rect 27798 36524 27804 36576
rect 27856 36564 27862 36576
rect 28031 36567 28089 36573
rect 28031 36564 28043 36567
rect 27856 36536 28043 36564
rect 27856 36524 27862 36536
rect 28031 36533 28043 36536
rect 28077 36533 28089 36567
rect 28031 36527 28089 36533
rect 28442 36524 28448 36576
rect 28500 36564 28506 36576
rect 28813 36567 28871 36573
rect 28813 36564 28825 36567
rect 28500 36536 28825 36564
rect 28500 36524 28506 36536
rect 28813 36533 28825 36536
rect 28859 36564 28871 36567
rect 29549 36567 29607 36573
rect 29549 36564 29561 36567
rect 28859 36536 29561 36564
rect 28859 36533 28871 36536
rect 28813 36527 28871 36533
rect 29549 36533 29561 36536
rect 29595 36564 29607 36567
rect 29840 36564 29868 36595
rect 30926 36592 30932 36604
rect 30984 36592 30990 36644
rect 31018 36564 31024 36576
rect 29595 36536 29868 36564
rect 30979 36536 31024 36564
rect 29595 36533 29607 36536
rect 29549 36527 29607 36533
rect 31018 36524 31024 36536
rect 31076 36524 31082 36576
rect 31379 36564 31407 36663
rect 31435 36635 31493 36641
rect 31435 36601 31447 36635
rect 31481 36632 31493 36635
rect 31481 36604 32444 36632
rect 31481 36601 31493 36604
rect 31435 36595 31493 36601
rect 31754 36564 31760 36576
rect 31379 36536 31760 36564
rect 31754 36524 31760 36536
rect 31812 36524 31818 36576
rect 32416 36564 32444 36604
rect 32490 36592 32496 36644
rect 32548 36632 32554 36644
rect 33594 36632 33600 36644
rect 32548 36604 32593 36632
rect 33106 36604 33600 36632
rect 32548 36592 32554 36604
rect 33106 36564 33134 36604
rect 33594 36592 33600 36604
rect 33652 36632 33658 36644
rect 33873 36635 33931 36641
rect 33873 36632 33885 36635
rect 33652 36604 33885 36632
rect 33652 36592 33658 36604
rect 33873 36601 33885 36604
rect 33919 36601 33931 36635
rect 33873 36595 33931 36601
rect 35544 36576 35572 36672
rect 38396 36672 38568 36700
rect 36630 36592 36636 36644
rect 36688 36632 36694 36644
rect 37138 36635 37196 36641
rect 37138 36632 37150 36635
rect 36688 36604 37150 36632
rect 36688 36592 36694 36604
rect 37138 36601 37150 36604
rect 37184 36601 37196 36635
rect 37138 36595 37196 36601
rect 32416 36536 33134 36564
rect 33505 36567 33563 36573
rect 33505 36533 33517 36567
rect 33551 36564 33563 36567
rect 33778 36564 33784 36576
rect 33551 36536 33784 36564
rect 33551 36533 33563 36536
rect 33505 36527 33563 36533
rect 33778 36524 33784 36536
rect 33836 36524 33842 36576
rect 35526 36564 35532 36576
rect 35487 36536 35532 36564
rect 35526 36524 35532 36536
rect 35584 36524 35590 36576
rect 36262 36564 36268 36576
rect 36223 36536 36268 36564
rect 36262 36524 36268 36536
rect 36320 36524 36326 36576
rect 37826 36524 37832 36576
rect 37884 36564 37890 36576
rect 38396 36573 38424 36672
rect 38562 36660 38568 36672
rect 38620 36660 38626 36712
rect 39022 36700 39028 36712
rect 38983 36672 39028 36700
rect 39022 36660 39028 36672
rect 39080 36660 39086 36712
rect 40129 36703 40187 36709
rect 40129 36669 40141 36703
rect 40175 36700 40187 36703
rect 40678 36700 40684 36712
rect 40175 36672 40684 36700
rect 40175 36669 40187 36672
rect 40129 36663 40187 36669
rect 40678 36660 40684 36672
rect 40736 36660 40742 36712
rect 42518 36709 42524 36712
rect 42496 36703 42524 36709
rect 42496 36700 42508 36703
rect 42431 36672 42508 36700
rect 42496 36669 42508 36672
rect 42576 36700 42582 36712
rect 43523 36709 43551 36740
rect 44361 36737 44373 36771
rect 44407 36768 44419 36771
rect 44545 36771 44603 36777
rect 44545 36768 44557 36771
rect 44407 36740 44557 36768
rect 44407 36737 44419 36740
rect 44361 36731 44419 36737
rect 44545 36737 44557 36740
rect 44591 36768 44603 36771
rect 46109 36771 46167 36777
rect 46109 36768 46121 36771
rect 44591 36740 46121 36768
rect 44591 36737 44603 36740
rect 44545 36731 44603 36737
rect 46109 36737 46121 36740
rect 46155 36737 46167 36771
rect 46109 36731 46167 36737
rect 42889 36703 42947 36709
rect 42889 36700 42901 36703
rect 42576 36672 42901 36700
rect 42496 36663 42524 36669
rect 42511 36660 42524 36663
rect 42576 36660 42582 36672
rect 42889 36669 42901 36672
rect 42935 36669 42947 36703
rect 42889 36663 42947 36669
rect 43508 36703 43566 36709
rect 43508 36669 43520 36703
rect 43554 36700 43566 36703
rect 43554 36672 43944 36700
rect 43554 36669 43566 36672
rect 43508 36663 43566 36669
rect 39301 36635 39359 36641
rect 39301 36601 39313 36635
rect 39347 36632 39359 36635
rect 40586 36632 40592 36644
rect 39347 36604 40592 36632
rect 39347 36601 39359 36604
rect 39301 36595 39359 36601
rect 40586 36592 40592 36604
rect 40644 36592 40650 36644
rect 41046 36592 41052 36644
rect 41104 36632 41110 36644
rect 41104 36604 41149 36632
rect 41104 36592 41110 36604
rect 38381 36567 38439 36573
rect 38381 36564 38393 36567
rect 37884 36536 38393 36564
rect 37884 36524 37890 36536
rect 38381 36533 38393 36536
rect 38427 36533 38439 36567
rect 38381 36527 38439 36533
rect 40034 36524 40040 36576
rect 40092 36564 40098 36576
rect 42511 36564 42539 36660
rect 43916 36576 43944 36672
rect 44266 36592 44272 36644
rect 44324 36632 44330 36644
rect 44637 36635 44695 36641
rect 44637 36632 44649 36635
rect 44324 36604 44649 36632
rect 44324 36592 44330 36604
rect 44637 36601 44649 36604
rect 44683 36601 44695 36635
rect 45186 36632 45192 36644
rect 45147 36604 45192 36632
rect 44637 36595 44695 36601
rect 43898 36564 43904 36576
rect 40092 36536 42539 36564
rect 43859 36536 43904 36564
rect 40092 36524 40098 36536
rect 43898 36524 43904 36536
rect 43956 36524 43962 36576
rect 44652 36564 44680 36595
rect 45186 36592 45192 36604
rect 45244 36592 45250 36644
rect 45465 36567 45523 36573
rect 45465 36564 45477 36567
rect 44652 36536 45477 36564
rect 45465 36533 45477 36536
rect 45511 36533 45523 36567
rect 46566 36564 46572 36576
rect 46527 36536 46572 36564
rect 45465 36527 45523 36533
rect 46566 36524 46572 36536
rect 46624 36524 46630 36576
rect 1104 36474 48852 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 48852 36474
rect 1104 36400 48852 36422
rect 15105 36363 15163 36369
rect 15105 36329 15117 36363
rect 15151 36360 15163 36363
rect 15286 36360 15292 36372
rect 15151 36332 15292 36360
rect 15151 36329 15163 36332
rect 15105 36323 15163 36329
rect 15286 36320 15292 36332
rect 15344 36320 15350 36372
rect 15470 36360 15476 36372
rect 15431 36332 15476 36360
rect 15470 36320 15476 36332
rect 15528 36320 15534 36372
rect 16025 36363 16083 36369
rect 16025 36329 16037 36363
rect 16071 36360 16083 36363
rect 16114 36360 16120 36372
rect 16071 36332 16120 36360
rect 16071 36329 16083 36332
rect 16025 36323 16083 36329
rect 16114 36320 16120 36332
rect 16172 36320 16178 36372
rect 17770 36360 17776 36372
rect 17731 36332 17776 36360
rect 17770 36320 17776 36332
rect 17828 36320 17834 36372
rect 19334 36320 19340 36372
rect 19392 36360 19398 36372
rect 19567 36363 19625 36369
rect 19567 36360 19579 36363
rect 19392 36332 19579 36360
rect 19392 36320 19398 36332
rect 19567 36329 19579 36332
rect 19613 36329 19625 36363
rect 20714 36360 20720 36372
rect 20675 36332 20720 36360
rect 19567 36323 19625 36329
rect 20714 36320 20720 36332
rect 20772 36320 20778 36372
rect 23934 36320 23940 36372
rect 23992 36360 23998 36372
rect 24029 36363 24087 36369
rect 24029 36360 24041 36363
rect 23992 36332 24041 36360
rect 23992 36320 23998 36332
rect 24029 36329 24041 36332
rect 24075 36329 24087 36363
rect 24029 36323 24087 36329
rect 25869 36363 25927 36369
rect 25869 36329 25881 36363
rect 25915 36360 25927 36363
rect 25958 36360 25964 36372
rect 25915 36332 25964 36360
rect 25915 36329 25927 36332
rect 25869 36323 25927 36329
rect 25958 36320 25964 36332
rect 26016 36360 26022 36372
rect 27709 36363 27767 36369
rect 26016 36332 26740 36360
rect 26016 36320 26022 36332
rect 14369 36295 14427 36301
rect 14369 36261 14381 36295
rect 14415 36292 14427 36295
rect 14550 36292 14556 36304
rect 14415 36264 14556 36292
rect 14415 36261 14427 36264
rect 14369 36255 14427 36261
rect 14550 36252 14556 36264
rect 14608 36292 14614 36304
rect 14645 36295 14703 36301
rect 14645 36292 14657 36295
rect 14608 36264 14657 36292
rect 14608 36252 14614 36264
rect 14645 36261 14657 36264
rect 14691 36261 14703 36295
rect 16482 36292 16488 36304
rect 16443 36264 16488 36292
rect 14645 36255 14703 36261
rect 16482 36252 16488 36264
rect 16540 36252 16546 36304
rect 20806 36252 20812 36304
rect 20864 36292 20870 36304
rect 23106 36292 23112 36304
rect 20864 36264 23112 36292
rect 20864 36252 20870 36264
rect 23106 36252 23112 36264
rect 23164 36292 23170 36304
rect 23201 36295 23259 36301
rect 23201 36292 23213 36295
rect 23164 36264 23213 36292
rect 23164 36252 23170 36264
rect 23201 36261 23213 36264
rect 23247 36292 23259 36295
rect 23842 36292 23848 36304
rect 23247 36264 23848 36292
rect 23247 36261 23259 36264
rect 23201 36255 23259 36261
rect 23842 36252 23848 36264
rect 23900 36252 23906 36304
rect 26326 36252 26332 36304
rect 26384 36292 26390 36304
rect 26712 36301 26740 36332
rect 27709 36329 27721 36363
rect 27755 36360 27767 36363
rect 27798 36360 27804 36372
rect 27755 36332 27804 36360
rect 27755 36329 27767 36332
rect 27709 36323 27767 36329
rect 27798 36320 27804 36332
rect 27856 36320 27862 36372
rect 29730 36360 29736 36372
rect 29691 36332 29736 36360
rect 29730 36320 29736 36332
rect 29788 36320 29794 36372
rect 32401 36363 32459 36369
rect 32401 36329 32413 36363
rect 32447 36360 32459 36363
rect 32490 36360 32496 36372
rect 32447 36332 32496 36360
rect 32447 36329 32459 36332
rect 32401 36323 32459 36329
rect 26605 36295 26663 36301
rect 26605 36292 26617 36295
rect 26384 36264 26617 36292
rect 26384 36252 26390 36264
rect 26605 36261 26617 36264
rect 26651 36261 26663 36295
rect 26605 36255 26663 36261
rect 26697 36295 26755 36301
rect 26697 36261 26709 36295
rect 26743 36292 26755 36295
rect 26786 36292 26792 36304
rect 26743 36264 26792 36292
rect 26743 36261 26755 36264
rect 26697 36255 26755 36261
rect 26786 36252 26792 36264
rect 26844 36252 26850 36304
rect 28534 36292 28540 36304
rect 28495 36264 28540 36292
rect 28534 36252 28540 36264
rect 28592 36252 28598 36304
rect 30282 36292 30288 36304
rect 30243 36264 30288 36292
rect 30282 36252 30288 36264
rect 30340 36252 30346 36304
rect 30374 36252 30380 36304
rect 30432 36292 30438 36304
rect 32416 36292 32444 36323
rect 32490 36320 32496 36332
rect 32548 36320 32554 36372
rect 33134 36320 33140 36372
rect 33192 36360 33198 36372
rect 38930 36360 38936 36372
rect 33192 36332 37780 36360
rect 38891 36332 38936 36360
rect 33192 36320 33198 36332
rect 33781 36295 33839 36301
rect 33781 36292 33793 36295
rect 30432 36264 32444 36292
rect 32508 36264 33793 36292
rect 30432 36252 30438 36264
rect 13630 36224 13636 36236
rect 13591 36196 13636 36224
rect 13630 36184 13636 36196
rect 13688 36184 13694 36236
rect 14182 36224 14188 36236
rect 14143 36196 14188 36224
rect 14182 36184 14188 36196
rect 14240 36184 14246 36236
rect 14918 36184 14924 36236
rect 14976 36224 14982 36236
rect 15324 36227 15382 36233
rect 15324 36224 15336 36227
rect 14976 36196 15336 36224
rect 14976 36184 14982 36196
rect 15324 36193 15336 36196
rect 15370 36193 15382 36227
rect 17862 36224 17868 36236
rect 17823 36196 17868 36224
rect 15324 36187 15382 36193
rect 17862 36184 17868 36196
rect 17920 36184 17926 36236
rect 18414 36224 18420 36236
rect 18375 36196 18420 36224
rect 18414 36184 18420 36196
rect 18472 36184 18478 36236
rect 19496 36227 19554 36233
rect 19496 36193 19508 36227
rect 19542 36224 19554 36227
rect 20254 36224 20260 36236
rect 19542 36196 20260 36224
rect 19542 36193 19554 36196
rect 19496 36187 19554 36193
rect 20254 36184 20260 36196
rect 20312 36184 20318 36236
rect 21726 36224 21732 36236
rect 21687 36196 21732 36224
rect 21726 36184 21732 36196
rect 21784 36184 21790 36236
rect 21910 36224 21916 36236
rect 21871 36196 21916 36224
rect 21910 36184 21916 36196
rect 21968 36184 21974 36236
rect 23753 36227 23811 36233
rect 23753 36193 23765 36227
rect 23799 36224 23811 36227
rect 24210 36224 24216 36236
rect 23799 36196 24216 36224
rect 23799 36193 23811 36196
rect 23753 36187 23811 36193
rect 24210 36184 24216 36196
rect 24268 36184 24274 36236
rect 24486 36184 24492 36236
rect 24544 36224 24550 36236
rect 24616 36227 24674 36233
rect 24616 36224 24628 36227
rect 24544 36196 24628 36224
rect 24544 36184 24550 36196
rect 24616 36193 24628 36196
rect 24662 36193 24674 36227
rect 24616 36187 24674 36193
rect 30926 36184 30932 36236
rect 30984 36224 30990 36236
rect 32508 36224 32536 36264
rect 33781 36261 33793 36264
rect 33827 36292 33839 36295
rect 34054 36292 34060 36304
rect 33827 36264 34060 36292
rect 33827 36261 33839 36264
rect 33781 36255 33839 36261
rect 34054 36252 34060 36264
rect 34112 36252 34118 36304
rect 34330 36292 34336 36304
rect 34291 36264 34336 36292
rect 34330 36252 34336 36264
rect 34388 36252 34394 36304
rect 36817 36295 36875 36301
rect 36817 36261 36829 36295
rect 36863 36292 36875 36295
rect 37090 36292 37096 36304
rect 36863 36264 37096 36292
rect 36863 36261 36875 36264
rect 36817 36255 36875 36261
rect 37090 36252 37096 36264
rect 37148 36252 37154 36304
rect 30984 36196 32536 36224
rect 36357 36227 36415 36233
rect 30984 36184 30990 36196
rect 36357 36193 36369 36227
rect 36403 36224 36415 36227
rect 36538 36224 36544 36236
rect 36403 36196 36544 36224
rect 36403 36193 36415 36196
rect 36357 36187 36415 36193
rect 36538 36184 36544 36196
rect 36596 36184 36602 36236
rect 36633 36227 36691 36233
rect 36633 36193 36645 36227
rect 36679 36224 36691 36227
rect 36722 36224 36728 36236
rect 36679 36196 36728 36224
rect 36679 36193 36691 36196
rect 36633 36187 36691 36193
rect 16390 36156 16396 36168
rect 16351 36128 16396 36156
rect 16390 36116 16396 36128
rect 16448 36116 16454 36168
rect 17034 36156 17040 36168
rect 16995 36128 17040 36156
rect 17034 36116 17040 36128
rect 17092 36116 17098 36168
rect 18506 36156 18512 36168
rect 18467 36128 18512 36156
rect 18506 36116 18512 36128
rect 18564 36116 18570 36168
rect 18782 36116 18788 36168
rect 18840 36156 18846 36168
rect 22186 36156 22192 36168
rect 18840 36128 19334 36156
rect 22147 36128 22192 36156
rect 18840 36116 18846 36128
rect 19306 36088 19334 36128
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 23109 36159 23167 36165
rect 23109 36125 23121 36159
rect 23155 36156 23167 36159
rect 23474 36156 23480 36168
rect 23155 36128 23480 36156
rect 23155 36125 23167 36128
rect 23109 36119 23167 36125
rect 23474 36116 23480 36128
rect 23532 36156 23538 36168
rect 24719 36159 24777 36165
rect 24719 36156 24731 36159
rect 23532 36128 24731 36156
rect 23532 36116 23538 36128
rect 24719 36125 24731 36128
rect 24765 36125 24777 36159
rect 26878 36156 26884 36168
rect 26839 36128 26884 36156
rect 24719 36119 24777 36125
rect 26878 36116 26884 36128
rect 26936 36116 26942 36168
rect 28445 36159 28503 36165
rect 28445 36125 28457 36159
rect 28491 36156 28503 36159
rect 28902 36156 28908 36168
rect 28491 36128 28908 36156
rect 28491 36125 28503 36128
rect 28445 36119 28503 36125
rect 28902 36116 28908 36128
rect 28960 36116 28966 36168
rect 30466 36116 30472 36168
rect 30524 36156 30530 36168
rect 30561 36159 30619 36165
rect 30561 36156 30573 36159
rect 30524 36128 30573 36156
rect 30524 36116 30530 36128
rect 30561 36125 30573 36128
rect 30607 36125 30619 36159
rect 30561 36119 30619 36125
rect 32306 36116 32312 36168
rect 32364 36156 32370 36168
rect 32493 36159 32551 36165
rect 32493 36156 32505 36159
rect 32364 36128 32505 36156
rect 32364 36116 32370 36128
rect 32493 36125 32505 36128
rect 32539 36125 32551 36159
rect 32493 36119 32551 36125
rect 32723 36159 32781 36165
rect 32723 36125 32735 36159
rect 32769 36156 32781 36159
rect 33686 36156 33692 36168
rect 32769 36128 33692 36156
rect 32769 36125 32781 36128
rect 32723 36119 32781 36125
rect 33686 36116 33692 36128
rect 33744 36116 33750 36168
rect 35897 36159 35955 36165
rect 34164 36128 34928 36156
rect 21726 36088 21732 36100
rect 19306 36060 21732 36088
rect 21726 36048 21732 36060
rect 21784 36048 21790 36100
rect 26234 36048 26240 36100
rect 26292 36088 26298 36100
rect 28997 36091 29055 36097
rect 28997 36088 29009 36091
rect 26292 36060 29009 36088
rect 26292 36048 26298 36060
rect 28997 36057 29009 36060
rect 29043 36088 29055 36091
rect 29362 36088 29368 36100
rect 29043 36060 29368 36088
rect 29043 36057 29055 36060
rect 28997 36051 29055 36057
rect 29362 36048 29368 36060
rect 29420 36048 29426 36100
rect 31386 36048 31392 36100
rect 31444 36088 31450 36100
rect 34164 36088 34192 36128
rect 31444 36060 34192 36088
rect 34900 36088 34928 36128
rect 35897 36125 35909 36159
rect 35943 36156 35955 36159
rect 36648 36156 36676 36187
rect 36722 36184 36728 36196
rect 36780 36184 36786 36236
rect 37752 36233 37780 36332
rect 38930 36320 38936 36332
rect 38988 36320 38994 36372
rect 40586 36360 40592 36372
rect 40547 36332 40592 36360
rect 40586 36320 40592 36332
rect 40644 36320 40650 36372
rect 43763 36363 43821 36369
rect 43763 36329 43775 36363
rect 43809 36360 43821 36363
rect 45922 36360 45928 36372
rect 43809 36332 45928 36360
rect 43809 36329 43821 36332
rect 43763 36323 43821 36329
rect 45922 36320 45928 36332
rect 45980 36360 45986 36372
rect 46566 36360 46572 36372
rect 45980 36332 46572 36360
rect 45980 36320 45986 36332
rect 46566 36320 46572 36332
rect 46624 36320 46630 36372
rect 40862 36252 40868 36304
rect 40920 36292 40926 36304
rect 41049 36295 41107 36301
rect 41049 36292 41061 36295
rect 40920 36264 41061 36292
rect 40920 36252 40926 36264
rect 41049 36261 41061 36264
rect 41095 36261 41107 36295
rect 41049 36255 41107 36261
rect 41138 36252 41144 36304
rect 41196 36292 41202 36304
rect 44545 36295 44603 36301
rect 44545 36292 44557 36295
rect 41196 36264 44557 36292
rect 41196 36252 41202 36264
rect 44545 36261 44557 36264
rect 44591 36292 44603 36295
rect 45005 36295 45063 36301
rect 45005 36292 45017 36295
rect 44591 36264 45017 36292
rect 44591 36261 44603 36264
rect 44545 36255 44603 36261
rect 45005 36261 45017 36264
rect 45051 36292 45063 36295
rect 45094 36292 45100 36304
rect 45051 36264 45100 36292
rect 45051 36261 45063 36264
rect 45005 36255 45063 36261
rect 45094 36252 45100 36264
rect 45152 36252 45158 36304
rect 37737 36227 37795 36233
rect 37737 36193 37749 36227
rect 37783 36224 37795 36227
rect 38197 36227 38255 36233
rect 38197 36224 38209 36227
rect 37783 36196 38209 36224
rect 37783 36193 37795 36196
rect 37737 36187 37795 36193
rect 38197 36193 38209 36196
rect 38243 36193 38255 36227
rect 38197 36187 38255 36193
rect 38838 36184 38844 36236
rect 38896 36224 38902 36236
rect 39117 36227 39175 36233
rect 39117 36224 39129 36227
rect 38896 36196 39129 36224
rect 38896 36184 38902 36196
rect 39117 36193 39129 36196
rect 39163 36193 39175 36227
rect 39117 36187 39175 36193
rect 39577 36227 39635 36233
rect 39577 36193 39589 36227
rect 39623 36193 39635 36227
rect 39577 36187 39635 36193
rect 43625 36227 43683 36233
rect 43625 36193 43637 36227
rect 43671 36224 43683 36227
rect 43714 36224 43720 36236
rect 43671 36196 43720 36224
rect 43671 36193 43683 36196
rect 43625 36187 43683 36193
rect 39022 36156 39028 36168
rect 35943 36128 36676 36156
rect 38580 36128 39028 36156
rect 35943 36125 35955 36128
rect 35897 36119 35955 36125
rect 37921 36091 37979 36097
rect 37921 36088 37933 36091
rect 34900 36060 37933 36088
rect 31444 36048 31450 36060
rect 37921 36057 37933 36060
rect 37967 36057 37979 36091
rect 37921 36051 37979 36057
rect 38580 36032 38608 36128
rect 39022 36116 39028 36128
rect 39080 36156 39086 36168
rect 39592 36156 39620 36187
rect 43714 36184 43720 36196
rect 43772 36184 43778 36236
rect 46382 36224 46388 36236
rect 46343 36196 46388 36224
rect 46382 36184 46388 36196
rect 46440 36184 46446 36236
rect 39850 36156 39856 36168
rect 39080 36128 39620 36156
rect 39811 36128 39856 36156
rect 39080 36116 39086 36128
rect 39850 36116 39856 36128
rect 39908 36116 39914 36168
rect 41506 36156 41512 36168
rect 41467 36128 41512 36156
rect 41506 36116 41512 36128
rect 41564 36156 41570 36168
rect 41969 36159 42027 36165
rect 41969 36156 41981 36159
rect 41564 36128 41981 36156
rect 41564 36116 41570 36128
rect 41969 36125 41981 36128
rect 42015 36125 42027 36159
rect 41969 36119 42027 36125
rect 44913 36159 44971 36165
rect 44913 36125 44925 36159
rect 44959 36125 44971 36159
rect 45186 36156 45192 36168
rect 45147 36128 45192 36156
rect 44913 36119 44971 36125
rect 19242 36020 19248 36032
rect 19203 35992 19248 36020
rect 19242 35980 19248 35992
rect 19300 35980 19306 36032
rect 21266 36020 21272 36032
rect 21227 35992 21272 36020
rect 21266 35980 21272 35992
rect 21324 35980 21330 36032
rect 26142 36020 26148 36032
rect 26103 35992 26148 36020
rect 26142 35980 26148 35992
rect 26200 35980 26206 36032
rect 27154 35980 27160 36032
rect 27212 36020 27218 36032
rect 29822 36020 29828 36032
rect 27212 35992 29828 36020
rect 27212 35980 27218 35992
rect 29822 35980 29828 35992
rect 29880 35980 29886 36032
rect 32858 35980 32864 36032
rect 32916 36020 32922 36032
rect 33045 36023 33103 36029
rect 33045 36020 33057 36023
rect 32916 35992 33057 36020
rect 32916 35980 32922 35992
rect 33045 35989 33057 35992
rect 33091 35989 33103 36023
rect 37090 36020 37096 36032
rect 37051 35992 37096 36020
rect 33045 35983 33103 35989
rect 37090 35980 37096 35992
rect 37148 35980 37154 36032
rect 38562 36020 38568 36032
rect 38523 35992 38568 36020
rect 38562 35980 38568 35992
rect 38620 35980 38626 36032
rect 44269 36023 44327 36029
rect 44269 35989 44281 36023
rect 44315 36020 44327 36023
rect 44358 36020 44364 36032
rect 44315 35992 44364 36020
rect 44315 35989 44327 35992
rect 44269 35983 44327 35989
rect 44358 35980 44364 35992
rect 44416 35980 44422 36032
rect 44928 36020 44956 36119
rect 45186 36116 45192 36128
rect 45244 36116 45250 36168
rect 45646 36020 45652 36032
rect 44928 35992 45652 36020
rect 45646 35980 45652 35992
rect 45704 36020 45710 36032
rect 46523 36023 46581 36029
rect 46523 36020 46535 36023
rect 45704 35992 46535 36020
rect 45704 35980 45710 35992
rect 46523 35989 46535 35992
rect 46569 35989 46581 36023
rect 46523 35983 46581 35989
rect 1104 35930 48852 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 48852 35930
rect 1104 35856 48852 35878
rect 14642 35816 14648 35828
rect 14603 35788 14648 35816
rect 14642 35776 14648 35788
rect 14700 35776 14706 35828
rect 15657 35819 15715 35825
rect 15657 35785 15669 35819
rect 15703 35816 15715 35819
rect 16393 35819 16451 35825
rect 16393 35816 16405 35819
rect 15703 35788 16405 35816
rect 15703 35785 15715 35788
rect 15657 35779 15715 35785
rect 16393 35785 16405 35788
rect 16439 35816 16451 35819
rect 16482 35816 16488 35828
rect 16439 35788 16488 35816
rect 16439 35785 16451 35788
rect 16393 35779 16451 35785
rect 16482 35776 16488 35788
rect 16540 35776 16546 35828
rect 16666 35816 16672 35828
rect 16627 35788 16672 35816
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 18598 35816 18604 35828
rect 18559 35788 18604 35816
rect 18598 35776 18604 35788
rect 18656 35776 18662 35828
rect 20254 35816 20260 35828
rect 20215 35788 20260 35816
rect 20254 35776 20260 35788
rect 20312 35776 20318 35828
rect 23106 35816 23112 35828
rect 23067 35788 23112 35816
rect 23106 35776 23112 35788
rect 23164 35776 23170 35828
rect 23474 35776 23480 35828
rect 23532 35816 23538 35828
rect 23799 35819 23857 35825
rect 23532 35788 23577 35816
rect 23532 35776 23538 35788
rect 23799 35785 23811 35819
rect 23845 35816 23857 35819
rect 24118 35816 24124 35828
rect 23845 35788 24124 35816
rect 23845 35785 23857 35788
rect 23799 35779 23857 35785
rect 24118 35776 24124 35788
rect 24176 35776 24182 35828
rect 24486 35776 24492 35828
rect 24544 35816 24550 35828
rect 24581 35819 24639 35825
rect 24581 35816 24593 35819
rect 24544 35788 24593 35816
rect 24544 35776 24550 35788
rect 24581 35785 24593 35788
rect 24627 35785 24639 35819
rect 24581 35779 24639 35785
rect 24903 35819 24961 35825
rect 24903 35785 24915 35819
rect 24949 35816 24961 35819
rect 26142 35816 26148 35828
rect 24949 35788 26148 35816
rect 24949 35785 24961 35788
rect 24903 35779 24961 35785
rect 26142 35776 26148 35788
rect 26200 35776 26206 35828
rect 26878 35816 26884 35828
rect 26839 35788 26884 35816
rect 26878 35776 26884 35788
rect 26936 35776 26942 35828
rect 28445 35819 28503 35825
rect 28445 35816 28457 35819
rect 27448 35788 28457 35816
rect 13262 35708 13268 35760
rect 13320 35748 13326 35760
rect 15746 35748 15752 35760
rect 13320 35720 15752 35748
rect 13320 35708 13326 35720
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 15838 35708 15844 35760
rect 15896 35748 15902 35760
rect 17865 35751 17923 35757
rect 17865 35748 17877 35751
rect 15896 35720 17877 35748
rect 15896 35708 15902 35720
rect 17865 35717 17877 35720
rect 17911 35748 17923 35751
rect 18414 35748 18420 35760
rect 17911 35720 18420 35748
rect 17911 35717 17923 35720
rect 17865 35711 17923 35717
rect 18414 35708 18420 35720
rect 18472 35748 18478 35760
rect 21085 35751 21143 35757
rect 21085 35748 21097 35751
rect 18472 35720 21097 35748
rect 18472 35708 18478 35720
rect 21085 35717 21097 35720
rect 21131 35748 21143 35751
rect 21910 35748 21916 35760
rect 21131 35720 21916 35748
rect 21131 35717 21143 35720
rect 21085 35711 21143 35717
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 24213 35751 24271 35757
rect 24213 35717 24225 35751
rect 24259 35748 24271 35751
rect 24302 35748 24308 35760
rect 24259 35720 24308 35748
rect 24259 35717 24271 35720
rect 24213 35711 24271 35717
rect 13081 35683 13139 35689
rect 13081 35649 13093 35683
rect 13127 35680 13139 35683
rect 14182 35680 14188 35692
rect 13127 35652 13676 35680
rect 13127 35649 13139 35652
rect 13081 35643 13139 35649
rect 13262 35612 13268 35624
rect 13223 35584 13268 35612
rect 13262 35572 13268 35584
rect 13320 35572 13326 35624
rect 13648 35621 13676 35652
rect 13786 35652 14188 35680
rect 13786 35624 13814 35652
rect 14182 35640 14188 35652
rect 14240 35680 14246 35692
rect 14277 35683 14335 35689
rect 14277 35680 14289 35683
rect 14240 35652 14289 35680
rect 14240 35640 14246 35652
rect 14277 35649 14289 35652
rect 14323 35680 14335 35683
rect 15856 35680 15884 35708
rect 14323 35652 15884 35680
rect 17083 35683 17141 35689
rect 14323 35649 14335 35652
rect 14277 35643 14335 35649
rect 17083 35649 17095 35683
rect 17129 35680 17141 35683
rect 19242 35680 19248 35692
rect 17129 35652 19248 35680
rect 17129 35649 17141 35652
rect 17083 35643 17141 35649
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 19889 35683 19947 35689
rect 19889 35649 19901 35683
rect 19935 35680 19947 35683
rect 19978 35680 19984 35692
rect 19935 35652 19984 35680
rect 19935 35649 19947 35652
rect 19889 35643 19947 35649
rect 19978 35640 19984 35652
rect 20036 35640 20042 35692
rect 21266 35680 21272 35692
rect 21227 35652 21272 35680
rect 21266 35640 21272 35652
rect 21324 35640 21330 35692
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 21784 35652 22324 35680
rect 21784 35640 21790 35652
rect 13633 35615 13691 35621
rect 13633 35581 13645 35615
rect 13679 35612 13691 35615
rect 13786 35612 13820 35624
rect 13679 35584 13820 35612
rect 13679 35581 13691 35584
rect 13633 35575 13691 35581
rect 13814 35572 13820 35584
rect 13872 35572 13878 35624
rect 13909 35615 13967 35621
rect 13909 35581 13921 35615
rect 13955 35612 13967 35615
rect 14734 35612 14740 35624
rect 13955 35584 14740 35612
rect 13955 35581 13967 35584
rect 13909 35575 13967 35581
rect 14734 35572 14740 35584
rect 14792 35572 14798 35624
rect 16996 35615 17054 35621
rect 16996 35581 17008 35615
rect 17042 35612 17054 35615
rect 17494 35612 17500 35624
rect 17042 35584 17500 35612
rect 17042 35581 17054 35584
rect 16996 35575 17054 35581
rect 17494 35572 17500 35584
rect 17552 35572 17558 35624
rect 18208 35615 18266 35621
rect 18208 35581 18220 35615
rect 18254 35612 18266 35615
rect 18598 35612 18604 35624
rect 18254 35584 18604 35612
rect 18254 35581 18266 35584
rect 18208 35575 18266 35581
rect 18598 35572 18604 35584
rect 18656 35572 18662 35624
rect 22296 35621 22324 35652
rect 22281 35615 22339 35621
rect 22281 35581 22293 35615
rect 22327 35612 22339 35615
rect 22925 35615 22983 35621
rect 22925 35612 22937 35615
rect 22327 35584 22937 35612
rect 22327 35581 22339 35584
rect 22281 35575 22339 35581
rect 22925 35581 22937 35584
rect 22971 35581 22983 35615
rect 22925 35575 22983 35581
rect 23728 35615 23786 35621
rect 23728 35581 23740 35615
rect 23774 35612 23786 35615
rect 24228 35612 24256 35711
rect 24302 35708 24308 35720
rect 24360 35748 24366 35760
rect 27448 35748 27476 35788
rect 28445 35785 28457 35788
rect 28491 35785 28503 35819
rect 28445 35779 28503 35785
rect 29411 35819 29469 35825
rect 29411 35785 29423 35819
rect 29457 35816 29469 35819
rect 29730 35816 29736 35828
rect 29457 35788 29736 35816
rect 29457 35785 29469 35788
rect 29411 35779 29469 35785
rect 29730 35776 29736 35788
rect 29788 35776 29794 35828
rect 30285 35819 30343 35825
rect 30285 35785 30297 35819
rect 30331 35816 30343 35819
rect 30374 35816 30380 35828
rect 30331 35788 30380 35816
rect 30331 35785 30343 35788
rect 30285 35779 30343 35785
rect 24360 35720 27476 35748
rect 27525 35751 27583 35757
rect 24360 35708 24366 35720
rect 27525 35717 27537 35751
rect 27571 35748 27583 35751
rect 28534 35748 28540 35760
rect 27571 35720 28540 35748
rect 27571 35717 27583 35720
rect 27525 35711 27583 35717
rect 23774 35584 24256 35612
rect 23774 35581 23786 35584
rect 23728 35575 23786 35581
rect 24578 35572 24584 35624
rect 24636 35612 24642 35624
rect 24800 35615 24858 35621
rect 24800 35612 24812 35615
rect 24636 35584 24812 35612
rect 24636 35572 24642 35584
rect 24800 35581 24812 35584
rect 24846 35612 24858 35615
rect 25225 35615 25283 35621
rect 25225 35612 25237 35615
rect 24846 35584 25237 35612
rect 24846 35581 24858 35584
rect 24800 35575 24858 35581
rect 25225 35581 25237 35584
rect 25271 35581 25283 35615
rect 25225 35575 25283 35581
rect 14642 35504 14648 35556
rect 14700 35544 14706 35556
rect 15058 35547 15116 35553
rect 15058 35544 15070 35547
rect 14700 35516 15070 35544
rect 14700 35504 14706 35516
rect 15058 35513 15070 35516
rect 15104 35513 15116 35547
rect 15058 35507 15116 35513
rect 14918 35436 14924 35488
rect 14976 35476 14982 35488
rect 15933 35479 15991 35485
rect 15933 35476 15945 35479
rect 14976 35448 15945 35476
rect 14976 35436 14982 35448
rect 15933 35445 15945 35448
rect 15979 35445 15991 35479
rect 17494 35476 17500 35488
rect 17455 35448 17500 35476
rect 15933 35439 15991 35445
rect 17494 35436 17500 35448
rect 17552 35436 17558 35488
rect 18279 35479 18337 35485
rect 18279 35445 18291 35479
rect 18325 35476 18337 35479
rect 18414 35476 18420 35488
rect 18325 35448 18420 35476
rect 18325 35445 18337 35448
rect 18279 35439 18337 35445
rect 18414 35436 18420 35448
rect 18472 35436 18478 35488
rect 18616 35476 18644 35572
rect 19061 35547 19119 35553
rect 19061 35513 19073 35547
rect 19107 35544 19119 35547
rect 19334 35544 19340 35556
rect 19107 35516 19340 35544
rect 19107 35513 19119 35516
rect 19061 35507 19119 35513
rect 19334 35504 19340 35516
rect 19392 35504 19398 35556
rect 20622 35504 20628 35556
rect 20680 35544 20686 35556
rect 20717 35547 20775 35553
rect 20717 35544 20729 35547
rect 20680 35516 20729 35544
rect 20680 35504 20686 35516
rect 20717 35513 20729 35516
rect 20763 35544 20775 35547
rect 21361 35547 21419 35553
rect 21361 35544 21373 35547
rect 20763 35516 21373 35544
rect 20763 35513 20775 35516
rect 20717 35507 20775 35513
rect 21361 35513 21373 35516
rect 21407 35513 21419 35547
rect 21361 35507 21419 35513
rect 21913 35547 21971 35553
rect 21913 35513 21925 35547
rect 21959 35544 21971 35547
rect 24026 35544 24032 35556
rect 21959 35516 24032 35544
rect 21959 35513 21971 35516
rect 21913 35507 21971 35513
rect 24026 35504 24032 35516
rect 24084 35544 24090 35556
rect 24210 35544 24216 35556
rect 24084 35516 24216 35544
rect 24084 35504 24090 35516
rect 24210 35504 24216 35516
rect 24268 35504 24274 35556
rect 25866 35544 25872 35556
rect 25827 35516 25872 35544
rect 25866 35504 25872 35516
rect 25924 35504 25930 35556
rect 25958 35504 25964 35556
rect 26016 35544 26022 35556
rect 26513 35547 26571 35553
rect 26016 35516 26061 35544
rect 26016 35504 26022 35516
rect 26513 35513 26525 35547
rect 26559 35544 26571 35547
rect 27540 35544 27568 35711
rect 28534 35708 28540 35720
rect 28592 35748 28598 35760
rect 28721 35751 28779 35757
rect 28721 35748 28733 35751
rect 28592 35720 28733 35748
rect 28592 35708 28598 35720
rect 28721 35717 28733 35720
rect 28767 35748 28779 35751
rect 30300 35748 30328 35779
rect 30374 35776 30380 35788
rect 30432 35776 30438 35828
rect 32033 35819 32091 35825
rect 32033 35785 32045 35819
rect 32079 35816 32091 35819
rect 32490 35816 32496 35828
rect 32079 35788 32496 35816
rect 32079 35785 32091 35788
rect 32033 35779 32091 35785
rect 32490 35776 32496 35788
rect 32548 35776 32554 35828
rect 33686 35776 33692 35828
rect 33744 35816 33750 35828
rect 34425 35819 34483 35825
rect 34425 35816 34437 35819
rect 33744 35788 34437 35816
rect 33744 35776 33750 35788
rect 34425 35785 34437 35788
rect 34471 35785 34483 35819
rect 36630 35816 36636 35828
rect 36591 35788 36636 35816
rect 34425 35779 34483 35785
rect 36630 35776 36636 35788
rect 36688 35776 36694 35828
rect 37642 35776 37648 35828
rect 37700 35816 37706 35828
rect 38838 35816 38844 35828
rect 37700 35788 38844 35816
rect 37700 35776 37706 35788
rect 38838 35776 38844 35788
rect 38896 35816 38902 35828
rect 39853 35819 39911 35825
rect 39853 35816 39865 35819
rect 38896 35788 39865 35816
rect 38896 35776 38902 35788
rect 39853 35785 39865 35788
rect 39899 35785 39911 35819
rect 39853 35779 39911 35785
rect 40313 35819 40371 35825
rect 40313 35785 40325 35819
rect 40359 35816 40371 35819
rect 40862 35816 40868 35828
rect 40359 35788 40868 35816
rect 40359 35785 40371 35788
rect 40313 35779 40371 35785
rect 40862 35776 40868 35788
rect 40920 35776 40926 35828
rect 41138 35776 41144 35828
rect 41196 35816 41202 35828
rect 41325 35819 41383 35825
rect 41325 35816 41337 35819
rect 41196 35788 41337 35816
rect 41196 35776 41202 35788
rect 41325 35785 41337 35788
rect 41371 35785 41383 35819
rect 41325 35779 41383 35785
rect 45094 35776 45100 35828
rect 45152 35816 45158 35828
rect 45189 35819 45247 35825
rect 45189 35816 45201 35819
rect 45152 35788 45201 35816
rect 45152 35776 45158 35788
rect 45189 35785 45201 35788
rect 45235 35785 45247 35819
rect 45646 35816 45652 35828
rect 45607 35788 45652 35816
rect 45189 35779 45247 35785
rect 45646 35776 45652 35788
rect 45704 35776 45710 35828
rect 28767 35720 30328 35748
rect 28767 35717 28779 35720
rect 28721 35711 28779 35717
rect 30466 35708 30472 35760
rect 30524 35748 30530 35760
rect 31021 35751 31079 35757
rect 31021 35748 31033 35751
rect 30524 35720 31033 35748
rect 30524 35708 30530 35720
rect 31021 35717 31033 35720
rect 31067 35748 31079 35751
rect 32122 35748 32128 35760
rect 31067 35720 32128 35748
rect 31067 35717 31079 35720
rect 31021 35711 31079 35717
rect 27709 35683 27767 35689
rect 27709 35649 27721 35683
rect 27755 35680 27767 35683
rect 27798 35680 27804 35692
rect 27755 35652 27804 35680
rect 27755 35649 27767 35652
rect 27709 35643 27767 35649
rect 27798 35640 27804 35652
rect 27856 35640 27862 35692
rect 29340 35615 29398 35621
rect 29340 35581 29352 35615
rect 29386 35612 29398 35615
rect 29730 35612 29736 35624
rect 29386 35584 29736 35612
rect 29386 35581 29398 35584
rect 29340 35575 29398 35581
rect 29730 35572 29736 35584
rect 29788 35572 29794 35624
rect 30653 35615 30711 35621
rect 30653 35581 30665 35615
rect 30699 35612 30711 35615
rect 30742 35612 30748 35624
rect 30699 35584 30748 35612
rect 30699 35581 30711 35584
rect 30653 35575 30711 35581
rect 30742 35572 30748 35584
rect 30800 35612 30806 35624
rect 31113 35615 31171 35621
rect 31113 35612 31125 35615
rect 30800 35584 31125 35612
rect 30800 35572 30806 35584
rect 31113 35581 31125 35584
rect 31159 35581 31171 35615
rect 31113 35575 31171 35581
rect 27801 35547 27859 35553
rect 27801 35544 27813 35547
rect 26559 35516 27476 35544
rect 27540 35516 27813 35544
rect 26559 35513 26571 35516
rect 26513 35507 26571 35513
rect 18966 35476 18972 35488
rect 18616 35448 18972 35476
rect 18966 35436 18972 35448
rect 19024 35476 19030 35488
rect 22830 35476 22836 35488
rect 19024 35448 22836 35476
rect 19024 35436 19030 35448
rect 22830 35436 22836 35448
rect 22888 35436 22894 35488
rect 22925 35479 22983 35485
rect 22925 35445 22937 35479
rect 22971 35476 22983 35479
rect 24946 35476 24952 35488
rect 22971 35448 24952 35476
rect 22971 35445 22983 35448
rect 22925 35439 22983 35445
rect 24946 35436 24952 35448
rect 25004 35436 25010 35488
rect 25685 35479 25743 35485
rect 25685 35445 25697 35479
rect 25731 35476 25743 35479
rect 25976 35476 26004 35504
rect 25731 35448 26004 35476
rect 27448 35476 27476 35516
rect 27801 35513 27813 35516
rect 27847 35513 27859 35547
rect 28350 35544 28356 35556
rect 28263 35516 28356 35544
rect 27801 35507 27859 35513
rect 28350 35504 28356 35516
rect 28408 35504 28414 35556
rect 31449 35553 31477 35720
rect 32122 35708 32128 35720
rect 32180 35748 32186 35760
rect 32677 35751 32735 35757
rect 32677 35748 32689 35751
rect 32180 35720 32689 35748
rect 32180 35708 32186 35720
rect 32677 35717 32689 35720
rect 32723 35717 32735 35751
rect 34054 35748 34060 35760
rect 34015 35720 34060 35748
rect 32677 35711 32735 35717
rect 28445 35547 28503 35553
rect 28445 35513 28457 35547
rect 28491 35544 28503 35547
rect 31434 35547 31492 35553
rect 28491 35516 29132 35544
rect 28491 35513 28503 35516
rect 28445 35507 28503 35513
rect 28368 35476 28396 35504
rect 28994 35476 29000 35488
rect 27448 35448 28396 35476
rect 28955 35448 29000 35476
rect 25731 35445 25743 35448
rect 25685 35439 25743 35445
rect 28994 35436 29000 35448
rect 29052 35436 29058 35488
rect 29104 35476 29132 35516
rect 31434 35513 31446 35547
rect 31480 35513 31492 35547
rect 32692 35544 32720 35711
rect 34054 35708 34060 35720
rect 34112 35708 34118 35760
rect 35989 35751 36047 35757
rect 35989 35717 36001 35751
rect 36035 35748 36047 35751
rect 37182 35748 37188 35760
rect 36035 35720 37188 35748
rect 36035 35717 36047 35720
rect 35989 35711 36047 35717
rect 37182 35708 37188 35720
rect 37240 35708 37246 35760
rect 38654 35748 38660 35760
rect 38615 35720 38660 35748
rect 38654 35708 38660 35720
rect 38712 35708 38718 35760
rect 39482 35708 39488 35760
rect 39540 35748 39546 35760
rect 45002 35748 45008 35760
rect 39540 35720 45008 35748
rect 39540 35708 39546 35720
rect 45002 35708 45008 35720
rect 45060 35748 45066 35760
rect 46382 35748 46388 35760
rect 45060 35720 46388 35748
rect 45060 35708 45066 35720
rect 46382 35708 46388 35720
rect 46440 35708 46446 35760
rect 36817 35683 36875 35689
rect 36817 35649 36829 35683
rect 36863 35680 36875 35683
rect 37090 35680 37096 35692
rect 36863 35652 37096 35680
rect 36863 35649 36875 35652
rect 36817 35643 36875 35649
rect 37090 35640 37096 35652
rect 37148 35640 37154 35692
rect 32858 35612 32864 35624
rect 32819 35584 32864 35612
rect 32858 35572 32864 35584
rect 32916 35572 32922 35624
rect 33778 35612 33784 35624
rect 33739 35584 33784 35612
rect 33778 35572 33784 35584
rect 33836 35572 33842 35624
rect 35713 35615 35771 35621
rect 35713 35581 35725 35615
rect 35759 35612 35771 35615
rect 35805 35615 35863 35621
rect 35805 35612 35817 35615
rect 35759 35584 35817 35612
rect 35759 35581 35771 35584
rect 35713 35575 35771 35581
rect 35805 35581 35817 35584
rect 35851 35612 35863 35615
rect 36722 35612 36728 35624
rect 35851 35584 36728 35612
rect 35851 35581 35863 35584
rect 35805 35575 35863 35581
rect 36722 35572 36728 35584
rect 36780 35572 36786 35624
rect 38102 35572 38108 35624
rect 38160 35612 38166 35624
rect 38672 35612 38700 35708
rect 41506 35640 41512 35692
rect 41564 35680 41570 35692
rect 41693 35683 41751 35689
rect 41693 35680 41705 35683
rect 41564 35652 41705 35680
rect 41564 35640 41570 35652
rect 41693 35649 41705 35652
rect 41739 35649 41751 35683
rect 41693 35643 41751 35649
rect 44913 35683 44971 35689
rect 44913 35649 44925 35683
rect 44959 35680 44971 35683
rect 45186 35680 45192 35692
rect 44959 35652 45192 35680
rect 44959 35649 44971 35652
rect 44913 35643 44971 35649
rect 45186 35640 45192 35652
rect 45244 35640 45250 35692
rect 38841 35615 38899 35621
rect 38841 35612 38853 35615
rect 38160 35584 38853 35612
rect 38160 35572 38166 35584
rect 38841 35581 38853 35584
rect 38887 35581 38899 35615
rect 38841 35575 38899 35581
rect 39301 35615 39359 35621
rect 39301 35581 39313 35615
rect 39347 35581 39359 35615
rect 39301 35575 39359 35581
rect 33182 35547 33240 35553
rect 33182 35544 33194 35547
rect 32692 35516 33194 35544
rect 31434 35507 31492 35513
rect 33182 35513 33194 35516
rect 33228 35544 33240 35547
rect 33318 35544 33324 35556
rect 33228 35516 33324 35544
rect 33228 35513 33240 35516
rect 33182 35507 33240 35513
rect 33318 35504 33324 35516
rect 33376 35504 33382 35556
rect 36630 35504 36636 35556
rect 36688 35544 36694 35556
rect 37138 35547 37196 35553
rect 37138 35544 37150 35547
rect 36688 35516 37150 35544
rect 36688 35504 36694 35516
rect 37138 35513 37150 35516
rect 37184 35544 37196 35547
rect 38010 35544 38016 35556
rect 37184 35516 38016 35544
rect 37184 35513 37196 35516
rect 37138 35507 37196 35513
rect 38010 35504 38016 35516
rect 38068 35504 38074 35556
rect 39316 35544 39344 35575
rect 39942 35572 39948 35624
rect 40000 35612 40006 35624
rect 40532 35615 40590 35621
rect 40532 35612 40544 35615
rect 40000 35584 40544 35612
rect 40000 35572 40006 35584
rect 40532 35581 40544 35584
rect 40578 35612 40590 35615
rect 40957 35615 41015 35621
rect 40957 35612 40969 35615
rect 40578 35584 40969 35612
rect 40578 35581 40590 35584
rect 40532 35575 40590 35581
rect 40957 35581 40969 35584
rect 41003 35581 41015 35615
rect 40957 35575 41015 35581
rect 42610 35572 42616 35624
rect 42668 35612 42674 35624
rect 43254 35621 43260 35624
rect 43232 35615 43260 35621
rect 43232 35612 43244 35615
rect 42668 35584 43244 35612
rect 42668 35572 42674 35584
rect 43232 35581 43244 35584
rect 43312 35612 43318 35624
rect 43993 35615 44051 35621
rect 43993 35612 44005 35615
rect 43312 35584 44005 35612
rect 43232 35575 43260 35581
rect 43254 35572 43260 35575
rect 43312 35572 43318 35584
rect 43993 35581 44005 35584
rect 44039 35581 44051 35615
rect 43993 35575 44051 35581
rect 38580 35516 39344 35544
rect 39577 35547 39635 35553
rect 38580 35488 38608 35516
rect 39577 35513 39589 35547
rect 39623 35544 39635 35547
rect 40402 35544 40408 35556
rect 39623 35516 40408 35544
rect 39623 35513 39635 35516
rect 39577 35507 39635 35513
rect 40402 35504 40408 35516
rect 40460 35504 40466 35556
rect 41782 35504 41788 35556
rect 41840 35544 41846 35556
rect 42337 35547 42395 35553
rect 41840 35516 41885 35544
rect 41840 35504 41846 35516
rect 42337 35513 42349 35547
rect 42383 35544 42395 35547
rect 42794 35544 42800 35556
rect 42383 35516 42800 35544
rect 42383 35513 42395 35516
rect 42337 35507 42395 35513
rect 42794 35504 42800 35516
rect 42852 35504 42858 35556
rect 44266 35544 44272 35556
rect 44227 35516 44272 35544
rect 44266 35504 44272 35516
rect 44324 35504 44330 35556
rect 44358 35504 44364 35556
rect 44416 35544 44422 35556
rect 44416 35516 44461 35544
rect 44416 35504 44422 35516
rect 32122 35476 32128 35488
rect 29104 35448 32128 35476
rect 32122 35436 32128 35448
rect 32180 35476 32186 35488
rect 32306 35476 32312 35488
rect 32180 35448 32312 35476
rect 32180 35436 32186 35448
rect 32306 35436 32312 35448
rect 32364 35436 32370 35488
rect 36357 35479 36415 35485
rect 36357 35445 36369 35479
rect 36403 35476 36415 35479
rect 36538 35476 36544 35488
rect 36403 35448 36544 35476
rect 36403 35445 36415 35448
rect 36357 35439 36415 35445
rect 36538 35436 36544 35448
rect 36596 35436 36602 35488
rect 37737 35479 37795 35485
rect 37737 35445 37749 35479
rect 37783 35476 37795 35479
rect 38194 35476 38200 35488
rect 37783 35448 38200 35476
rect 37783 35445 37795 35448
rect 37737 35439 37795 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 38381 35479 38439 35485
rect 38381 35445 38393 35479
rect 38427 35476 38439 35479
rect 38562 35476 38568 35488
rect 38427 35448 38568 35476
rect 38427 35445 38439 35448
rect 38381 35439 38439 35445
rect 38562 35436 38568 35448
rect 38620 35436 38626 35488
rect 40635 35479 40693 35485
rect 40635 35445 40647 35479
rect 40681 35476 40693 35479
rect 40862 35476 40868 35488
rect 40681 35448 40868 35476
rect 40681 35445 40693 35448
rect 40635 35439 40693 35445
rect 40862 35436 40868 35448
rect 40920 35436 40926 35488
rect 43303 35479 43361 35485
rect 43303 35445 43315 35479
rect 43349 35476 43361 35479
rect 43438 35476 43444 35488
rect 43349 35448 43444 35476
rect 43349 35445 43361 35448
rect 43303 35439 43361 35445
rect 43438 35436 43444 35448
rect 43496 35436 43502 35488
rect 43714 35476 43720 35488
rect 43675 35448 43720 35476
rect 43714 35436 43720 35448
rect 43772 35436 43778 35488
rect 1104 35386 48852 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 48852 35386
rect 1104 35312 48852 35334
rect 14734 35272 14740 35284
rect 14695 35244 14740 35272
rect 14734 35232 14740 35244
rect 14792 35232 14798 35284
rect 15473 35275 15531 35281
rect 15473 35241 15485 35275
rect 15519 35272 15531 35275
rect 15838 35272 15844 35284
rect 15519 35244 15844 35272
rect 15519 35241 15531 35244
rect 15473 35235 15531 35241
rect 15838 35232 15844 35244
rect 15896 35232 15902 35284
rect 16209 35275 16267 35281
rect 16209 35241 16221 35275
rect 16255 35272 16267 35275
rect 16390 35272 16396 35284
rect 16255 35244 16396 35272
rect 16255 35241 16267 35244
rect 16209 35235 16267 35241
rect 16390 35232 16396 35244
rect 16448 35232 16454 35284
rect 18874 35272 18880 35284
rect 18835 35244 18880 35272
rect 18874 35232 18880 35244
rect 18932 35232 18938 35284
rect 20993 35275 21051 35281
rect 20993 35241 21005 35275
rect 21039 35272 21051 35275
rect 21266 35272 21272 35284
rect 21039 35244 21272 35272
rect 21039 35241 21051 35244
rect 20993 35235 21051 35241
rect 21266 35232 21272 35244
rect 21324 35232 21330 35284
rect 22554 35272 22560 35284
rect 22515 35244 22560 35272
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 23109 35275 23167 35281
rect 23109 35241 23121 35275
rect 23155 35272 23167 35275
rect 23155 35244 23474 35272
rect 23155 35241 23167 35244
rect 23109 35235 23167 35241
rect 16482 35204 16488 35216
rect 16443 35176 16488 35204
rect 16482 35164 16488 35176
rect 16540 35164 16546 35216
rect 23446 35204 23474 35244
rect 26326 35232 26332 35284
rect 26384 35272 26390 35284
rect 26697 35275 26755 35281
rect 26697 35272 26709 35275
rect 26384 35244 26709 35272
rect 26384 35232 26390 35244
rect 26697 35241 26709 35244
rect 26743 35241 26755 35275
rect 30282 35272 30288 35284
rect 30243 35244 30288 35272
rect 26697 35235 26755 35241
rect 30282 35232 30288 35244
rect 30340 35232 30346 35284
rect 30742 35272 30748 35284
rect 30703 35244 30748 35272
rect 30742 35232 30748 35244
rect 30800 35232 30806 35284
rect 32398 35272 32404 35284
rect 32359 35244 32404 35272
rect 32398 35232 32404 35244
rect 32456 35232 32462 35284
rect 33318 35272 33324 35284
rect 33279 35244 33324 35272
rect 33318 35232 33324 35244
rect 33376 35232 33382 35284
rect 33873 35275 33931 35281
rect 33873 35241 33885 35275
rect 33919 35272 33931 35275
rect 34054 35272 34060 35284
rect 33919 35244 34060 35272
rect 33919 35241 33931 35244
rect 33873 35235 33931 35241
rect 34054 35232 34060 35244
rect 34112 35232 34118 35284
rect 38562 35232 38568 35284
rect 38620 35272 38626 35284
rect 39209 35275 39267 35281
rect 39209 35272 39221 35275
rect 38620 35244 39221 35272
rect 38620 35232 38626 35244
rect 39209 35241 39221 35244
rect 39255 35241 39267 35275
rect 39209 35235 39267 35241
rect 41509 35275 41567 35281
rect 41509 35241 41521 35275
rect 41555 35272 41567 35275
rect 41555 35244 43576 35272
rect 41555 35241 41567 35244
rect 41509 35235 41567 35241
rect 43548 35216 43576 35244
rect 44266 35232 44272 35284
rect 44324 35272 44330 35284
rect 44453 35275 44511 35281
rect 44453 35272 44465 35275
rect 44324 35244 44465 35272
rect 44324 35232 44330 35244
rect 44453 35241 44465 35244
rect 44499 35272 44511 35275
rect 46615 35275 46673 35281
rect 46615 35272 46627 35275
rect 44499 35244 46627 35272
rect 44499 35241 44511 35244
rect 44453 35235 44511 35241
rect 46615 35241 46627 35244
rect 46661 35241 46673 35275
rect 46615 35235 46673 35241
rect 24118 35204 24124 35216
rect 23446 35176 24124 35204
rect 24118 35164 24124 35176
rect 24176 35164 24182 35216
rect 28442 35204 28448 35216
rect 28403 35176 28448 35204
rect 28442 35164 28448 35176
rect 28500 35164 28506 35216
rect 28997 35207 29055 35213
rect 28997 35173 29009 35207
rect 29043 35204 29055 35207
rect 29362 35204 29368 35216
rect 29043 35176 29368 35204
rect 29043 35173 29055 35176
rect 28997 35167 29055 35173
rect 29362 35164 29368 35176
rect 29420 35164 29426 35216
rect 34701 35207 34759 35213
rect 34701 35173 34713 35207
rect 34747 35204 34759 35207
rect 35618 35204 35624 35216
rect 34747 35176 35624 35204
rect 34747 35173 34759 35176
rect 34701 35167 34759 35173
rect 35618 35164 35624 35176
rect 35676 35164 35682 35216
rect 36817 35207 36875 35213
rect 36817 35173 36829 35207
rect 36863 35204 36875 35207
rect 37090 35204 37096 35216
rect 36863 35176 37096 35204
rect 36863 35173 36875 35176
rect 36817 35167 36875 35173
rect 37090 35164 37096 35176
rect 37148 35164 37154 35216
rect 38010 35164 38016 35216
rect 38068 35204 38074 35216
rect 38334 35207 38392 35213
rect 38334 35204 38346 35207
rect 38068 35176 38346 35204
rect 38068 35164 38074 35176
rect 38334 35173 38346 35176
rect 38380 35173 38392 35207
rect 38334 35167 38392 35173
rect 40678 35164 40684 35216
rect 40736 35204 40742 35216
rect 40910 35207 40968 35213
rect 40910 35204 40922 35207
rect 40736 35176 40922 35204
rect 40736 35164 40742 35176
rect 40910 35173 40922 35176
rect 40956 35173 40968 35207
rect 43530 35204 43536 35216
rect 43443 35176 43536 35204
rect 40910 35167 40968 35173
rect 43530 35164 43536 35176
rect 43588 35164 43594 35216
rect 45094 35204 45100 35216
rect 45055 35176 45100 35204
rect 45094 35164 45100 35176
rect 45152 35164 45158 35216
rect 15289 35139 15347 35145
rect 15289 35105 15301 35139
rect 15335 35136 15347 35139
rect 16022 35136 16028 35148
rect 15335 35108 16028 35136
rect 15335 35105 15347 35108
rect 15289 35099 15347 35105
rect 16022 35096 16028 35108
rect 16080 35096 16086 35148
rect 18506 35136 18512 35148
rect 18467 35108 18512 35136
rect 18506 35096 18512 35108
rect 18564 35096 18570 35148
rect 22186 35136 22192 35148
rect 22147 35108 22192 35136
rect 22186 35096 22192 35108
rect 22244 35096 22250 35148
rect 27246 35136 27252 35148
rect 27207 35108 27252 35136
rect 27246 35096 27252 35108
rect 27304 35096 27310 35148
rect 30742 35136 30748 35148
rect 30703 35108 30748 35136
rect 30742 35096 30748 35108
rect 30800 35096 30806 35148
rect 31021 35139 31079 35145
rect 31021 35105 31033 35139
rect 31067 35136 31079 35139
rect 31202 35136 31208 35148
rect 31067 35108 31208 35136
rect 31067 35105 31079 35108
rect 31021 35099 31079 35105
rect 31202 35096 31208 35108
rect 31260 35096 31266 35148
rect 32214 35096 32220 35148
rect 32272 35136 32278 35148
rect 34146 35136 34152 35148
rect 32272 35108 34152 35136
rect 32272 35096 32278 35108
rect 34146 35096 34152 35108
rect 34204 35096 34210 35148
rect 34790 35096 34796 35148
rect 34848 35136 34854 35148
rect 34885 35139 34943 35145
rect 34885 35136 34897 35139
rect 34848 35108 34897 35136
rect 34848 35096 34854 35108
rect 34885 35105 34897 35108
rect 34931 35105 34943 35139
rect 36078 35136 36084 35148
rect 34885 35099 34943 35105
rect 35176 35108 36084 35136
rect 16393 35071 16451 35077
rect 16393 35037 16405 35071
rect 16439 35068 16451 35071
rect 16574 35068 16580 35080
rect 16439 35040 16580 35068
rect 16439 35037 16451 35040
rect 16393 35031 16451 35037
rect 16574 35028 16580 35040
rect 16632 35028 16638 35080
rect 17034 35068 17040 35080
rect 16947 35040 17040 35068
rect 17034 35028 17040 35040
rect 17092 35068 17098 35080
rect 18598 35068 18604 35080
rect 17092 35040 18604 35068
rect 17092 35028 17098 35040
rect 18598 35028 18604 35040
rect 18656 35028 18662 35080
rect 24026 35068 24032 35080
rect 23987 35040 24032 35068
rect 24026 35028 24032 35040
rect 24084 35028 24090 35080
rect 24302 35068 24308 35080
rect 24263 35040 24308 35068
rect 24302 35028 24308 35040
rect 24360 35028 24366 35080
rect 28353 35071 28411 35077
rect 28353 35068 28365 35071
rect 27816 35040 28365 35068
rect 27816 34944 27844 35040
rect 28353 35037 28365 35040
rect 28399 35037 28411 35071
rect 32950 35068 32956 35080
rect 32911 35040 32956 35068
rect 28353 35031 28411 35037
rect 32950 35028 32956 35040
rect 33008 35028 33014 35080
rect 34164 35068 34192 35096
rect 35176 35068 35204 35108
rect 36078 35096 36084 35108
rect 36136 35096 36142 35148
rect 36633 35139 36691 35145
rect 36633 35105 36645 35139
rect 36679 35136 36691 35139
rect 36722 35136 36728 35148
rect 36679 35108 36728 35136
rect 36679 35105 36691 35108
rect 36633 35099 36691 35105
rect 36722 35096 36728 35108
rect 36780 35096 36786 35148
rect 39850 35096 39856 35148
rect 39908 35136 39914 35148
rect 40589 35139 40647 35145
rect 40589 35136 40601 35139
rect 39908 35108 40601 35136
rect 39908 35096 39914 35108
rect 40589 35105 40601 35108
rect 40635 35105 40647 35139
rect 40589 35099 40647 35105
rect 46544 35139 46602 35145
rect 46544 35105 46556 35139
rect 46590 35136 46602 35139
rect 46934 35136 46940 35148
rect 46590 35108 46940 35136
rect 46590 35105 46602 35108
rect 46544 35099 46602 35105
rect 46934 35096 46940 35108
rect 46992 35096 46998 35148
rect 34164 35040 35204 35068
rect 35253 35071 35311 35077
rect 35253 35037 35265 35071
rect 35299 35068 35311 35071
rect 36170 35068 36176 35080
rect 35299 35040 36176 35068
rect 35299 35037 35311 35040
rect 35253 35031 35311 35037
rect 36170 35028 36176 35040
rect 36228 35028 36234 35080
rect 38010 35068 38016 35080
rect 37971 35040 38016 35068
rect 38010 35028 38016 35040
rect 38068 35028 38074 35080
rect 43162 35028 43168 35080
rect 43220 35068 43226 35080
rect 43441 35071 43499 35077
rect 43441 35068 43453 35071
rect 43220 35040 43453 35068
rect 43220 35028 43226 35040
rect 43441 35037 43453 35040
rect 43487 35068 43499 35071
rect 43622 35068 43628 35080
rect 43487 35040 43628 35068
rect 43487 35037 43499 35040
rect 43441 35031 43499 35037
rect 43622 35028 43628 35040
rect 43680 35028 43686 35080
rect 43717 35071 43775 35077
rect 43717 35037 43729 35071
rect 43763 35037 43775 35071
rect 43717 35031 43775 35037
rect 45005 35071 45063 35077
rect 45005 35037 45017 35071
rect 45051 35068 45063 35071
rect 45186 35068 45192 35080
rect 45051 35040 45192 35068
rect 45051 35037 45063 35040
rect 45005 35031 45063 35037
rect 29822 34960 29828 35012
rect 29880 35000 29886 35012
rect 35802 35000 35808 35012
rect 29880 34972 35808 35000
rect 29880 34960 29886 34972
rect 35802 34960 35808 34972
rect 35860 34960 35866 35012
rect 38933 35003 38991 35009
rect 38933 34969 38945 35003
rect 38979 35000 38991 35003
rect 41782 35000 41788 35012
rect 38979 34972 41788 35000
rect 38979 34969 38991 34972
rect 38933 34963 38991 34969
rect 41782 34960 41788 34972
rect 41840 34960 41846 35012
rect 42794 34960 42800 35012
rect 42852 35000 42858 35012
rect 43732 35000 43760 35031
rect 45186 35028 45192 35040
rect 45244 35028 45250 35080
rect 45373 35071 45431 35077
rect 45373 35037 45385 35071
rect 45419 35037 45431 35071
rect 45373 35031 45431 35037
rect 42852 34972 43760 35000
rect 42852 34960 42858 34972
rect 13262 34932 13268 34944
rect 13223 34904 13268 34932
rect 13262 34892 13268 34904
rect 13320 34892 13326 34944
rect 13630 34932 13636 34944
rect 13591 34904 13636 34932
rect 13630 34892 13636 34904
rect 13688 34892 13694 34944
rect 17218 34892 17224 34944
rect 17276 34932 17282 34944
rect 17862 34932 17868 34944
rect 17276 34904 17868 34932
rect 17276 34892 17282 34904
rect 17862 34892 17868 34904
rect 17920 34892 17926 34944
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 19429 34935 19487 34941
rect 19429 34932 19441 34935
rect 19392 34904 19441 34932
rect 19392 34892 19398 34904
rect 19429 34901 19441 34904
rect 19475 34932 19487 34935
rect 20622 34932 20628 34944
rect 19475 34904 20628 34932
rect 19475 34901 19487 34904
rect 19429 34895 19487 34901
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 25590 34932 25596 34944
rect 25551 34904 25596 34932
rect 25590 34892 25596 34904
rect 25648 34892 25654 34944
rect 25866 34932 25872 34944
rect 25827 34904 25872 34932
rect 25866 34892 25872 34904
rect 25924 34892 25930 34944
rect 27387 34935 27445 34941
rect 27387 34901 27399 34935
rect 27433 34932 27445 34935
rect 27798 34932 27804 34944
rect 27433 34904 27804 34932
rect 27433 34901 27445 34904
rect 27387 34895 27445 34901
rect 27798 34892 27804 34904
rect 27856 34892 27862 34944
rect 35342 34892 35348 34944
rect 35400 34932 35406 34944
rect 35529 34935 35587 34941
rect 35529 34932 35541 34935
rect 35400 34904 35541 34932
rect 35400 34892 35406 34904
rect 35529 34901 35541 34904
rect 35575 34901 35587 34935
rect 37182 34932 37188 34944
rect 37143 34904 37188 34932
rect 35529 34895 35587 34901
rect 37182 34892 37188 34904
rect 37240 34892 37246 34944
rect 43732 34932 43760 34972
rect 45388 34944 45416 35031
rect 45370 34932 45376 34944
rect 43732 34904 45376 34932
rect 45370 34892 45376 34904
rect 45428 34892 45434 34944
rect 1104 34842 48852 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 48852 34842
rect 1104 34768 48852 34790
rect 14642 34728 14648 34740
rect 14603 34700 14648 34728
rect 14642 34688 14648 34700
rect 14700 34688 14706 34740
rect 15749 34731 15807 34737
rect 15749 34697 15761 34731
rect 15795 34728 15807 34731
rect 16482 34728 16488 34740
rect 15795 34700 16488 34728
rect 15795 34697 15807 34700
rect 15749 34691 15807 34697
rect 16482 34688 16488 34700
rect 16540 34688 16546 34740
rect 16574 34688 16580 34740
rect 16632 34728 16638 34740
rect 16761 34731 16819 34737
rect 16761 34728 16773 34731
rect 16632 34700 16773 34728
rect 16632 34688 16638 34700
rect 16761 34697 16773 34700
rect 16807 34697 16819 34731
rect 16761 34691 16819 34697
rect 17865 34731 17923 34737
rect 17865 34697 17877 34731
rect 17911 34728 17923 34731
rect 18506 34728 18512 34740
rect 17911 34700 18512 34728
rect 17911 34697 17923 34700
rect 17865 34691 17923 34697
rect 18506 34688 18512 34700
rect 18564 34688 18570 34740
rect 20622 34728 20628 34740
rect 20583 34700 20628 34728
rect 20622 34688 20628 34700
rect 20680 34688 20686 34740
rect 21913 34731 21971 34737
rect 21913 34697 21925 34731
rect 21959 34728 21971 34731
rect 22186 34728 22192 34740
rect 21959 34700 22192 34728
rect 21959 34697 21971 34700
rect 21913 34691 21971 34697
rect 22186 34688 22192 34700
rect 22244 34688 22250 34740
rect 22830 34688 22836 34740
rect 22888 34728 22894 34740
rect 23017 34731 23075 34737
rect 23017 34728 23029 34731
rect 22888 34700 23029 34728
rect 22888 34688 22894 34700
rect 23017 34697 23029 34700
rect 23063 34697 23075 34731
rect 24118 34728 24124 34740
rect 24079 34700 24124 34728
rect 23017 34691 23075 34697
rect 24118 34688 24124 34700
rect 24176 34688 24182 34740
rect 27798 34728 27804 34740
rect 27759 34700 27804 34728
rect 27798 34688 27804 34700
rect 27856 34688 27862 34740
rect 28123 34731 28181 34737
rect 28123 34697 28135 34731
rect 28169 34728 28181 34731
rect 28994 34728 29000 34740
rect 28169 34700 29000 34728
rect 28169 34697 28181 34700
rect 28123 34691 28181 34697
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 29822 34728 29828 34740
rect 29783 34700 29828 34728
rect 29822 34688 29828 34700
rect 29880 34688 29886 34740
rect 30742 34688 30748 34740
rect 30800 34728 30806 34740
rect 31205 34731 31263 34737
rect 31205 34728 31217 34731
rect 30800 34700 31217 34728
rect 30800 34688 30806 34700
rect 31205 34697 31217 34700
rect 31251 34728 31263 34731
rect 33410 34728 33416 34740
rect 31251 34700 33416 34728
rect 31251 34697 31263 34700
rect 31205 34691 31263 34697
rect 33410 34688 33416 34700
rect 33468 34688 33474 34740
rect 33502 34688 33508 34740
rect 33560 34728 33566 34740
rect 36078 34728 36084 34740
rect 33560 34700 35985 34728
rect 36039 34700 36084 34728
rect 33560 34688 33566 34700
rect 16022 34660 16028 34672
rect 15983 34632 16028 34660
rect 16022 34620 16028 34632
rect 16080 34620 16086 34672
rect 16390 34620 16396 34672
rect 16448 34660 16454 34672
rect 18601 34663 18659 34669
rect 18601 34660 18613 34663
rect 16448 34632 18613 34660
rect 16448 34620 16454 34632
rect 18601 34629 18613 34632
rect 18647 34660 18659 34663
rect 18874 34660 18880 34672
rect 18647 34632 18880 34660
rect 18647 34629 18659 34632
rect 18601 34623 18659 34629
rect 18874 34620 18880 34632
rect 18932 34620 18938 34672
rect 21358 34660 21364 34672
rect 21319 34632 21364 34660
rect 21358 34620 21364 34632
rect 21416 34620 21422 34672
rect 22281 34663 22339 34669
rect 22281 34629 22293 34663
rect 22327 34660 22339 34663
rect 22554 34660 22560 34672
rect 22327 34632 22560 34660
rect 22327 34629 22339 34632
rect 22281 34623 22339 34629
rect 22554 34620 22560 34632
rect 22612 34660 22618 34672
rect 23106 34660 23112 34672
rect 22612 34632 23112 34660
rect 22612 34620 22618 34632
rect 23106 34620 23112 34632
rect 23164 34620 23170 34672
rect 23477 34663 23535 34669
rect 23477 34629 23489 34663
rect 23523 34660 23535 34663
rect 24026 34660 24032 34672
rect 23523 34632 24032 34660
rect 23523 34629 23535 34632
rect 23477 34623 23535 34629
rect 24026 34620 24032 34632
rect 24084 34620 24090 34672
rect 27706 34620 27712 34672
rect 27764 34660 27770 34672
rect 29411 34663 29469 34669
rect 29411 34660 29423 34663
rect 27764 34632 29423 34660
rect 27764 34620 27770 34632
rect 29411 34629 29423 34632
rect 29457 34629 29469 34663
rect 29411 34623 29469 34629
rect 29546 34620 29552 34672
rect 29604 34660 29610 34672
rect 33318 34660 33324 34672
rect 29604 34632 31375 34660
rect 33279 34632 33324 34660
rect 29604 34620 29610 34632
rect 17420 34564 18368 34592
rect 13538 34524 13544 34536
rect 13499 34496 13544 34524
rect 13538 34484 13544 34496
rect 13596 34484 13602 34536
rect 13814 34524 13820 34536
rect 13786 34484 13820 34524
rect 13872 34524 13878 34536
rect 14001 34527 14059 34533
rect 13872 34496 13917 34524
rect 13872 34484 13878 34496
rect 14001 34493 14013 34527
rect 14047 34524 14059 34527
rect 14826 34524 14832 34536
rect 14047 34496 14832 34524
rect 14047 34493 14059 34496
rect 14001 34487 14059 34493
rect 14826 34484 14832 34496
rect 14884 34484 14890 34536
rect 17420 34533 17448 34564
rect 16996 34527 17054 34533
rect 16996 34493 17008 34527
rect 17042 34524 17054 34527
rect 17405 34527 17463 34533
rect 17405 34524 17417 34527
rect 17042 34496 17417 34524
rect 17042 34493 17054 34496
rect 16996 34487 17054 34493
rect 17405 34493 17417 34496
rect 17451 34493 17463 34527
rect 18046 34524 18052 34536
rect 18007 34496 18052 34524
rect 17405 34487 17463 34493
rect 18046 34484 18052 34496
rect 18104 34484 18110 34536
rect 13173 34459 13231 34465
rect 13173 34425 13185 34459
rect 13219 34456 13231 34459
rect 13786 34456 13814 34484
rect 13219 34428 13814 34456
rect 13219 34425 13231 34428
rect 13173 34419 13231 34425
rect 14642 34416 14648 34468
rect 14700 34456 14706 34468
rect 15150 34459 15208 34465
rect 15150 34456 15162 34459
rect 14700 34428 15162 34456
rect 14700 34416 14706 34428
rect 15150 34425 15162 34428
rect 15196 34425 15208 34459
rect 15150 34419 15208 34425
rect 17083 34459 17141 34465
rect 17083 34425 17095 34459
rect 17129 34456 17141 34459
rect 18340 34456 18368 34564
rect 18414 34552 18420 34604
rect 18472 34592 18478 34604
rect 19245 34595 19303 34601
rect 19245 34592 19257 34595
rect 18472 34564 19257 34592
rect 18472 34552 18478 34564
rect 19245 34561 19257 34564
rect 19291 34592 19303 34595
rect 19426 34592 19432 34604
rect 19291 34564 19432 34592
rect 19291 34561 19303 34564
rect 19245 34555 19303 34561
rect 19426 34552 19432 34564
rect 19484 34552 19490 34604
rect 19886 34592 19892 34604
rect 19847 34564 19892 34592
rect 19886 34552 19892 34564
rect 19944 34552 19950 34604
rect 20254 34552 20260 34604
rect 20312 34592 20318 34604
rect 27246 34592 27252 34604
rect 20312 34564 27252 34592
rect 20312 34552 20318 34564
rect 27246 34552 27252 34564
rect 27304 34552 27310 34604
rect 28442 34592 28448 34604
rect 28403 34564 28448 34592
rect 28442 34552 28448 34564
rect 28500 34552 28506 34604
rect 28534 34552 28540 34604
rect 28592 34592 28598 34604
rect 28813 34595 28871 34601
rect 28813 34592 28825 34595
rect 28592 34564 28825 34592
rect 28592 34552 28598 34564
rect 28813 34561 28825 34564
rect 28859 34561 28871 34595
rect 28813 34555 28871 34561
rect 30193 34595 30251 34601
rect 30193 34561 30205 34595
rect 30239 34592 30251 34595
rect 31202 34592 31208 34604
rect 30239 34564 31208 34592
rect 30239 34561 30251 34564
rect 30193 34555 30251 34561
rect 31202 34552 31208 34564
rect 31260 34552 31266 34604
rect 31347 34592 31375 34632
rect 33318 34620 33324 34632
rect 33376 34620 33382 34672
rect 35957 34660 35985 34700
rect 36078 34688 36084 34700
rect 36136 34688 36142 34740
rect 37918 34688 37924 34740
rect 37976 34728 37982 34740
rect 38105 34731 38163 34737
rect 38105 34728 38117 34731
rect 37976 34700 38117 34728
rect 37976 34688 37982 34700
rect 38105 34697 38117 34700
rect 38151 34728 38163 34731
rect 38473 34731 38531 34737
rect 38473 34728 38485 34731
rect 38151 34700 38485 34728
rect 38151 34697 38163 34700
rect 38105 34691 38163 34697
rect 38473 34697 38485 34700
rect 38519 34697 38531 34731
rect 39850 34728 39856 34740
rect 39811 34700 39856 34728
rect 38473 34691 38531 34697
rect 36909 34663 36967 34669
rect 36909 34660 36921 34663
rect 35957 34632 36921 34660
rect 36909 34629 36921 34632
rect 36955 34629 36967 34663
rect 36909 34623 36967 34629
rect 31754 34592 31760 34604
rect 31347 34564 31760 34592
rect 22624 34527 22682 34533
rect 22624 34493 22636 34527
rect 22670 34524 22682 34527
rect 22830 34524 22836 34536
rect 22670 34496 22836 34524
rect 22670 34493 22682 34496
rect 22624 34487 22682 34493
rect 22830 34484 22836 34496
rect 22888 34484 22894 34536
rect 23566 34524 23572 34536
rect 23527 34496 23572 34524
rect 23566 34484 23572 34496
rect 23624 34524 23630 34536
rect 24302 34524 24308 34536
rect 23624 34496 24308 34524
rect 23624 34484 23630 34496
rect 24302 34484 24308 34496
rect 24360 34524 24366 34536
rect 24489 34527 24547 34533
rect 24489 34524 24501 34527
rect 24360 34496 24501 34524
rect 24360 34484 24366 34496
rect 24489 34493 24501 34496
rect 24535 34493 24547 34527
rect 24489 34487 24547 34493
rect 28052 34527 28110 34533
rect 28052 34493 28064 34527
rect 28098 34524 28110 34527
rect 28460 34524 28488 34552
rect 28098 34496 28488 34524
rect 28098 34493 28110 34496
rect 28052 34487 28110 34493
rect 28626 34484 28632 34536
rect 28684 34524 28690 34536
rect 29340 34527 29398 34533
rect 29340 34524 29352 34527
rect 28684 34496 29352 34524
rect 28684 34484 28690 34496
rect 29340 34493 29352 34496
rect 29386 34524 29398 34527
rect 29822 34524 29828 34536
rect 29386 34496 29828 34524
rect 29386 34493 29398 34496
rect 29340 34487 29398 34493
rect 29822 34484 29828 34496
rect 29880 34484 29886 34536
rect 31347 34533 31375 34564
rect 31754 34552 31760 34564
rect 31812 34552 31818 34604
rect 32950 34552 32956 34604
rect 33008 34592 33014 34604
rect 33045 34595 33103 34601
rect 33045 34592 33057 34595
rect 33008 34564 33057 34592
rect 33008 34552 33014 34564
rect 33045 34561 33057 34564
rect 33091 34592 33103 34595
rect 33689 34595 33747 34601
rect 33689 34592 33701 34595
rect 33091 34564 33701 34592
rect 33091 34561 33103 34564
rect 33045 34555 33103 34561
rect 33689 34561 33701 34564
rect 33735 34561 33747 34595
rect 33689 34555 33747 34561
rect 30336 34527 30394 34533
rect 30336 34493 30348 34527
rect 30382 34524 30394 34527
rect 31332 34527 31390 34533
rect 30382 34496 30598 34524
rect 30382 34493 30394 34496
rect 30336 34487 30394 34493
rect 19334 34456 19340 34468
rect 17129 34428 18184 34456
rect 18340 34428 19196 34456
rect 19295 34428 19340 34456
rect 17129 34425 17141 34428
rect 17083 34419 17141 34425
rect 18156 34400 18184 34428
rect 18138 34348 18144 34400
rect 18196 34348 18202 34400
rect 18279 34391 18337 34397
rect 18279 34357 18291 34391
rect 18325 34388 18337 34391
rect 18506 34388 18512 34400
rect 18325 34360 18512 34388
rect 18325 34357 18337 34360
rect 18279 34351 18337 34357
rect 18506 34348 18512 34360
rect 18564 34348 18570 34400
rect 19058 34388 19064 34400
rect 19019 34360 19064 34388
rect 19058 34348 19064 34360
rect 19116 34348 19122 34400
rect 19168 34388 19196 34428
rect 19334 34416 19340 34428
rect 19392 34416 19398 34468
rect 20257 34459 20315 34465
rect 20257 34425 20269 34459
rect 20303 34456 20315 34459
rect 20806 34456 20812 34468
rect 20303 34428 20812 34456
rect 20303 34425 20315 34428
rect 20257 34419 20315 34425
rect 20806 34416 20812 34428
rect 20864 34416 20870 34468
rect 20901 34459 20959 34465
rect 20901 34425 20913 34459
rect 20947 34425 20959 34459
rect 23799 34459 23857 34465
rect 23799 34456 23811 34459
rect 20901 34419 20959 34425
rect 22572 34428 23811 34456
rect 20346 34388 20352 34400
rect 19168 34360 20352 34388
rect 20346 34348 20352 34360
rect 20404 34348 20410 34400
rect 20622 34348 20628 34400
rect 20680 34388 20686 34400
rect 20916 34388 20944 34419
rect 22572 34400 22600 34428
rect 23799 34425 23811 34428
rect 23845 34425 23857 34459
rect 25590 34456 25596 34468
rect 25551 34428 25596 34456
rect 23799 34419 23857 34425
rect 25590 34416 25596 34428
rect 25648 34416 25654 34468
rect 25685 34459 25743 34465
rect 25685 34425 25697 34459
rect 25731 34425 25743 34459
rect 25685 34419 25743 34425
rect 26237 34459 26295 34465
rect 26237 34425 26249 34459
rect 26283 34456 26295 34459
rect 26878 34456 26884 34468
rect 26283 34428 26884 34456
rect 26283 34425 26295 34428
rect 26237 34419 26295 34425
rect 20680 34360 20944 34388
rect 20680 34348 20686 34360
rect 22554 34348 22560 34400
rect 22612 34348 22618 34400
rect 22695 34391 22753 34397
rect 22695 34357 22707 34391
rect 22741 34388 22753 34391
rect 22922 34388 22928 34400
rect 22741 34360 22928 34388
rect 22741 34357 22753 34360
rect 22695 34351 22753 34357
rect 22922 34348 22928 34360
rect 22980 34348 22986 34400
rect 25130 34348 25136 34400
rect 25188 34388 25194 34400
rect 25317 34391 25375 34397
rect 25317 34388 25329 34391
rect 25188 34360 25329 34388
rect 25188 34348 25194 34360
rect 25317 34357 25329 34360
rect 25363 34388 25375 34391
rect 25700 34388 25728 34419
rect 26878 34416 26884 34428
rect 26936 34416 26942 34468
rect 30423 34459 30481 34465
rect 30423 34456 30435 34459
rect 27448 34428 30435 34456
rect 25363 34360 25728 34388
rect 25363 34357 25375 34360
rect 25317 34351 25375 34357
rect 26694 34348 26700 34400
rect 26752 34388 26758 34400
rect 27448 34388 27476 34428
rect 30423 34425 30435 34428
rect 30469 34425 30481 34459
rect 30423 34419 30481 34425
rect 26752 34360 27476 34388
rect 26752 34348 26758 34360
rect 28074 34348 28080 34400
rect 28132 34388 28138 34400
rect 30570 34388 30598 34496
rect 31332 34493 31344 34527
rect 31378 34493 31390 34527
rect 31332 34487 31390 34493
rect 31478 34484 31484 34536
rect 31536 34524 31542 34536
rect 32125 34527 32183 34533
rect 32125 34524 32137 34527
rect 31536 34496 32137 34524
rect 31536 34484 31542 34496
rect 32125 34493 32137 34496
rect 32171 34524 32183 34527
rect 32309 34527 32367 34533
rect 32309 34524 32321 34527
rect 32171 34496 32321 34524
rect 32171 34493 32183 34496
rect 32125 34487 32183 34493
rect 32309 34493 32321 34496
rect 32355 34493 32367 34527
rect 32309 34487 32367 34493
rect 32398 34484 32404 34536
rect 32456 34524 32462 34536
rect 32769 34527 32827 34533
rect 32769 34524 32781 34527
rect 32456 34496 32781 34524
rect 32456 34484 32462 34496
rect 32769 34493 32781 34496
rect 32815 34493 32827 34527
rect 32769 34487 32827 34493
rect 34333 34527 34391 34533
rect 34333 34493 34345 34527
rect 34379 34524 34391 34527
rect 35618 34524 35624 34536
rect 34379 34496 35624 34524
rect 34379 34493 34391 34496
rect 34333 34487 34391 34493
rect 35618 34484 35624 34496
rect 35676 34484 35682 34536
rect 36924 34524 36952 34623
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34592 37887 34595
rect 38010 34592 38016 34604
rect 37875 34564 38016 34592
rect 37875 34561 37887 34564
rect 37829 34555 37887 34561
rect 38010 34552 38016 34564
rect 38068 34552 38074 34604
rect 38488 34592 38516 34691
rect 39850 34688 39856 34700
rect 39908 34688 39914 34740
rect 40313 34731 40371 34737
rect 40313 34697 40325 34731
rect 40359 34728 40371 34731
rect 40678 34728 40684 34740
rect 40359 34700 40684 34728
rect 40359 34697 40371 34700
rect 40313 34691 40371 34697
rect 40678 34688 40684 34700
rect 40736 34688 40742 34740
rect 43530 34728 43536 34740
rect 43491 34700 43536 34728
rect 43530 34688 43536 34700
rect 43588 34688 43594 34740
rect 45186 34688 45192 34740
rect 45244 34728 45250 34740
rect 45373 34731 45431 34737
rect 45373 34728 45385 34731
rect 45244 34700 45385 34728
rect 45244 34688 45250 34700
rect 45373 34697 45385 34700
rect 45419 34697 45431 34731
rect 45373 34691 45431 34697
rect 39577 34663 39635 34669
rect 39577 34629 39589 34663
rect 39623 34660 39635 34663
rect 45005 34663 45063 34669
rect 45005 34660 45017 34663
rect 39623 34632 45017 34660
rect 39623 34629 39635 34632
rect 39577 34623 39635 34629
rect 45005 34629 45017 34632
rect 45051 34660 45063 34663
rect 45094 34660 45100 34672
rect 45051 34632 45100 34660
rect 45051 34629 45063 34632
rect 45005 34623 45063 34629
rect 45094 34620 45100 34632
rect 45152 34620 45158 34672
rect 38488 34564 39021 34592
rect 36998 34524 37004 34536
rect 36911 34496 37004 34524
rect 36998 34484 37004 34496
rect 37056 34524 37062 34536
rect 37093 34527 37151 34533
rect 37093 34524 37105 34527
rect 37056 34496 37105 34524
rect 37056 34484 37062 34496
rect 37093 34493 37105 34496
rect 37139 34493 37151 34527
rect 37093 34487 37151 34493
rect 37182 34484 37188 34536
rect 37240 34524 37246 34536
rect 37645 34527 37703 34533
rect 37645 34524 37657 34527
rect 37240 34496 37657 34524
rect 37240 34484 37246 34496
rect 37645 34493 37657 34496
rect 37691 34493 37703 34527
rect 38654 34524 38660 34536
rect 38615 34496 38660 34524
rect 37645 34487 37703 34493
rect 34701 34459 34759 34465
rect 34701 34425 34713 34459
rect 34747 34456 34759 34459
rect 34790 34456 34796 34468
rect 34747 34428 34796 34456
rect 34747 34425 34759 34428
rect 34701 34419 34759 34425
rect 34790 34416 34796 34428
rect 34848 34456 34854 34468
rect 35158 34456 35164 34468
rect 34848 34428 35164 34456
rect 34848 34416 34854 34428
rect 35158 34416 35164 34428
rect 35216 34416 35222 34468
rect 37660 34456 37688 34487
rect 38654 34484 38660 34496
rect 38712 34484 38718 34536
rect 38562 34456 38568 34468
rect 37660 34428 38568 34456
rect 38562 34416 38568 34428
rect 38620 34416 38626 34468
rect 38993 34465 39021 34564
rect 40402 34552 40408 34604
rect 40460 34592 40466 34604
rect 40681 34595 40739 34601
rect 40681 34592 40693 34595
rect 40460 34564 40693 34592
rect 40460 34552 40466 34564
rect 40681 34561 40693 34564
rect 40727 34592 40739 34595
rect 41877 34595 41935 34601
rect 41877 34592 41889 34595
rect 40727 34564 41889 34592
rect 40727 34561 40739 34564
rect 40681 34555 40739 34561
rect 41877 34561 41889 34564
rect 41923 34561 41935 34595
rect 42794 34592 42800 34604
rect 42755 34564 42800 34592
rect 41877 34555 41935 34561
rect 42794 34552 42800 34564
rect 42852 34552 42858 34604
rect 43438 34552 43444 34604
rect 43496 34592 43502 34604
rect 44085 34595 44143 34601
rect 44085 34592 44097 34595
rect 43496 34564 44097 34592
rect 43496 34552 43502 34564
rect 44085 34561 44097 34564
rect 44131 34592 44143 34595
rect 44542 34592 44548 34604
rect 44131 34564 44548 34592
rect 44131 34561 44143 34564
rect 44085 34555 44143 34561
rect 44542 34552 44548 34564
rect 44600 34552 44606 34604
rect 41601 34527 41659 34533
rect 41601 34493 41613 34527
rect 41647 34524 41659 34527
rect 42245 34527 42303 34533
rect 42245 34524 42257 34527
rect 41647 34496 42257 34524
rect 41647 34493 41659 34496
rect 41601 34487 41659 34493
rect 42245 34493 42257 34496
rect 42291 34493 42303 34527
rect 42245 34487 42303 34493
rect 38978 34459 39036 34465
rect 38978 34425 38990 34459
rect 39024 34425 39036 34459
rect 38978 34419 39036 34425
rect 40678 34416 40684 34468
rect 40736 34456 40742 34468
rect 41002 34459 41060 34465
rect 41002 34456 41014 34459
rect 40736 34428 41014 34456
rect 40736 34416 40742 34428
rect 41002 34425 41014 34428
rect 41048 34425 41060 34459
rect 41002 34419 41060 34425
rect 30745 34391 30803 34397
rect 30745 34388 30757 34391
rect 28132 34360 30757 34388
rect 28132 34348 28138 34360
rect 30745 34357 30757 34360
rect 30791 34357 30803 34391
rect 30745 34351 30803 34357
rect 31202 34348 31208 34400
rect 31260 34388 31266 34400
rect 31435 34391 31493 34397
rect 31435 34388 31447 34391
rect 31260 34360 31447 34388
rect 31260 34348 31266 34360
rect 31435 34357 31447 34360
rect 31481 34357 31493 34391
rect 35250 34388 35256 34400
rect 35211 34360 35256 34388
rect 31435 34351 31493 34357
rect 35250 34348 35256 34360
rect 35308 34348 35314 34400
rect 36541 34391 36599 34397
rect 36541 34357 36553 34391
rect 36587 34388 36599 34391
rect 36722 34388 36728 34400
rect 36587 34360 36728 34388
rect 36587 34357 36599 34360
rect 36541 34351 36599 34357
rect 36722 34348 36728 34360
rect 36780 34348 36786 34400
rect 42260 34388 42288 34487
rect 44818 34484 44824 34536
rect 44876 34524 44882 34536
rect 46144 34527 46202 34533
rect 46144 34524 46156 34527
rect 44876 34496 46156 34524
rect 44876 34484 44882 34496
rect 46144 34493 46156 34496
rect 46190 34524 46202 34527
rect 46569 34527 46627 34533
rect 46569 34524 46581 34527
rect 46190 34496 46581 34524
rect 46190 34493 46202 34496
rect 46144 34487 46202 34493
rect 46569 34493 46581 34496
rect 46615 34493 46627 34527
rect 46569 34487 46627 34493
rect 42518 34456 42524 34468
rect 42479 34428 42524 34456
rect 42518 34416 42524 34428
rect 42576 34416 42582 34468
rect 42613 34459 42671 34465
rect 42613 34425 42625 34459
rect 42659 34425 42671 34459
rect 42613 34419 42671 34425
rect 42628 34388 42656 34419
rect 43806 34416 43812 34468
rect 43864 34456 43870 34468
rect 43901 34459 43959 34465
rect 43901 34456 43913 34459
rect 43864 34428 43913 34456
rect 43864 34416 43870 34428
rect 43901 34425 43913 34428
rect 43947 34456 43959 34459
rect 44177 34459 44235 34465
rect 44177 34456 44189 34459
rect 43947 34428 44189 34456
rect 43947 34425 43959 34428
rect 43901 34419 43959 34425
rect 44177 34425 44189 34428
rect 44223 34456 44235 34459
rect 44358 34456 44364 34468
rect 44223 34428 44364 34456
rect 44223 34425 44235 34428
rect 44177 34419 44235 34425
rect 44358 34416 44364 34428
rect 44416 34416 44422 34468
rect 44726 34456 44732 34468
rect 44639 34428 44732 34456
rect 44726 34416 44732 34428
rect 44784 34416 44790 34468
rect 42260 34360 42656 34388
rect 44266 34348 44272 34400
rect 44324 34388 44330 34400
rect 44744 34388 44772 34416
rect 44324 34360 44772 34388
rect 44324 34348 44330 34360
rect 45094 34348 45100 34400
rect 45152 34388 45158 34400
rect 46247 34391 46305 34397
rect 46247 34388 46259 34391
rect 45152 34360 46259 34388
rect 45152 34348 45158 34360
rect 46247 34357 46259 34360
rect 46293 34357 46305 34391
rect 46934 34388 46940 34400
rect 46895 34360 46940 34388
rect 46247 34351 46305 34357
rect 46934 34348 46940 34360
rect 46992 34348 46998 34400
rect 1104 34298 48852 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 48852 34298
rect 1104 34224 48852 34246
rect 13354 34184 13360 34196
rect 13267 34156 13360 34184
rect 13354 34144 13360 34156
rect 13412 34184 13418 34196
rect 13538 34184 13544 34196
rect 13412 34156 13544 34184
rect 13412 34144 13418 34156
rect 13538 34144 13544 34156
rect 13596 34144 13602 34196
rect 14826 34184 14832 34196
rect 14787 34156 14832 34184
rect 14826 34144 14832 34156
rect 14884 34144 14890 34196
rect 15565 34187 15623 34193
rect 15565 34153 15577 34187
rect 15611 34184 15623 34187
rect 15654 34184 15660 34196
rect 15611 34156 15660 34184
rect 15611 34153 15623 34156
rect 15565 34147 15623 34153
rect 15654 34144 15660 34156
rect 15712 34144 15718 34196
rect 16390 34184 16396 34196
rect 16351 34156 16396 34184
rect 16390 34144 16396 34156
rect 16448 34144 16454 34196
rect 16945 34187 17003 34193
rect 16945 34153 16957 34187
rect 16991 34184 17003 34187
rect 16991 34156 18000 34184
rect 16991 34153 17003 34156
rect 16945 34147 17003 34153
rect 17972 34128 18000 34156
rect 18046 34144 18052 34196
rect 18104 34184 18110 34196
rect 19058 34184 19064 34196
rect 18104 34156 19064 34184
rect 18104 34144 18110 34156
rect 19058 34144 19064 34156
rect 19116 34144 19122 34196
rect 19245 34187 19303 34193
rect 19245 34153 19257 34187
rect 19291 34184 19303 34187
rect 19334 34184 19340 34196
rect 19291 34156 19340 34184
rect 19291 34153 19303 34156
rect 19245 34147 19303 34153
rect 19334 34144 19340 34156
rect 19392 34144 19398 34196
rect 19426 34144 19432 34196
rect 19484 34184 19490 34196
rect 19521 34187 19579 34193
rect 19521 34184 19533 34187
rect 19484 34156 19533 34184
rect 19484 34144 19490 34156
rect 19521 34153 19533 34156
rect 19567 34153 19579 34187
rect 19521 34147 19579 34153
rect 20806 34144 20812 34196
rect 20864 34184 20870 34196
rect 21039 34187 21097 34193
rect 21039 34184 21051 34187
rect 20864 34156 21051 34184
rect 20864 34144 20870 34156
rect 21039 34153 21051 34156
rect 21085 34153 21097 34187
rect 21039 34147 21097 34153
rect 22922 34144 22928 34196
rect 22980 34184 22986 34196
rect 24029 34187 24087 34193
rect 24029 34184 24041 34187
rect 22980 34156 24041 34184
rect 22980 34144 22986 34156
rect 24029 34153 24041 34156
rect 24075 34184 24087 34187
rect 24118 34184 24124 34196
rect 24075 34156 24124 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 24118 34144 24124 34156
rect 24176 34144 24182 34196
rect 31481 34187 31539 34193
rect 31481 34153 31493 34187
rect 31527 34184 31539 34187
rect 32398 34184 32404 34196
rect 31527 34156 32404 34184
rect 31527 34153 31539 34156
rect 31481 34147 31539 34153
rect 32398 34144 32404 34156
rect 32456 34144 32462 34196
rect 34793 34187 34851 34193
rect 34793 34153 34805 34187
rect 34839 34184 34851 34187
rect 35618 34184 35624 34196
rect 34839 34156 35624 34184
rect 34839 34153 34851 34156
rect 34793 34147 34851 34153
rect 35618 34144 35624 34156
rect 35676 34144 35682 34196
rect 36722 34184 36728 34196
rect 36683 34156 36728 34184
rect 36722 34144 36728 34156
rect 36780 34144 36786 34196
rect 38010 34184 38016 34196
rect 37971 34156 38016 34184
rect 38010 34144 38016 34156
rect 38068 34144 38074 34196
rect 38194 34144 38200 34196
rect 38252 34184 38258 34196
rect 42518 34184 42524 34196
rect 38252 34156 41184 34184
rect 42479 34156 42524 34184
rect 38252 34144 38258 34156
rect 17678 34116 17684 34128
rect 17639 34088 17684 34116
rect 17678 34076 17684 34088
rect 17736 34076 17742 34128
rect 17954 34116 17960 34128
rect 17867 34088 17960 34116
rect 17954 34076 17960 34088
rect 18012 34076 18018 34128
rect 18509 34119 18567 34125
rect 18509 34085 18521 34119
rect 18555 34116 18567 34119
rect 18598 34116 18604 34128
rect 18555 34088 18604 34116
rect 18555 34085 18567 34088
rect 18509 34079 18567 34085
rect 18598 34076 18604 34088
rect 18656 34076 18662 34128
rect 19935 34119 19993 34125
rect 19935 34085 19947 34119
rect 19981 34116 19993 34119
rect 24765 34119 24823 34125
rect 19981 34088 23474 34116
rect 19981 34085 19993 34088
rect 19935 34079 19993 34085
rect 16022 33980 16028 33992
rect 15983 33952 16028 33980
rect 16022 33940 16028 33952
rect 16080 33940 16086 33992
rect 17696 33980 17724 34076
rect 19848 34051 19906 34057
rect 19848 34017 19860 34051
rect 19894 34048 19906 34051
rect 20162 34048 20168 34060
rect 19894 34020 20168 34048
rect 19894 34017 19906 34020
rect 19848 34011 19906 34017
rect 20162 34008 20168 34020
rect 20220 34008 20226 34060
rect 20714 34008 20720 34060
rect 20772 34048 20778 34060
rect 20936 34051 20994 34057
rect 20936 34048 20948 34051
rect 20772 34020 20948 34048
rect 20772 34008 20778 34020
rect 20936 34017 20948 34020
rect 20982 34017 20994 34051
rect 22738 34048 22744 34060
rect 22699 34020 22744 34048
rect 20936 34011 20994 34017
rect 22738 34008 22744 34020
rect 22796 34008 22802 34060
rect 23198 34048 23204 34060
rect 23159 34020 23204 34048
rect 23198 34008 23204 34020
rect 23256 34008 23262 34060
rect 17865 33983 17923 33989
rect 17865 33980 17877 33983
rect 17696 33952 17877 33980
rect 17865 33949 17877 33952
rect 17911 33949 17923 33983
rect 23290 33980 23296 33992
rect 23251 33952 23296 33980
rect 17865 33943 17923 33949
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 23446 33980 23474 34088
rect 24765 34085 24777 34119
rect 24811 34116 24823 34119
rect 25130 34116 25136 34128
rect 24811 34088 25136 34116
rect 24811 34085 24823 34088
rect 24765 34079 24823 34085
rect 25130 34076 25136 34088
rect 25188 34076 25194 34128
rect 26602 34076 26608 34128
rect 26660 34116 26666 34128
rect 26697 34119 26755 34125
rect 26697 34116 26709 34119
rect 26660 34088 26709 34116
rect 26660 34076 26666 34088
rect 26697 34085 26709 34088
rect 26743 34116 26755 34119
rect 28261 34119 28319 34125
rect 28261 34116 28273 34119
rect 26743 34088 28273 34116
rect 26743 34085 26755 34088
rect 26697 34079 26755 34085
rect 28261 34085 28273 34088
rect 28307 34085 28319 34119
rect 28261 34079 28319 34085
rect 29730 34076 29736 34128
rect 29788 34116 29794 34128
rect 29825 34119 29883 34125
rect 29825 34116 29837 34119
rect 29788 34088 29837 34116
rect 29788 34076 29794 34088
rect 29825 34085 29837 34088
rect 29871 34085 29883 34119
rect 29825 34079 29883 34085
rect 32214 34048 32220 34060
rect 32175 34020 32220 34048
rect 32214 34008 32220 34020
rect 32272 34008 32278 34060
rect 32416 34048 32444 34144
rect 32858 34116 32864 34128
rect 32819 34088 32864 34116
rect 32858 34076 32864 34088
rect 32916 34076 32922 34128
rect 34977 34119 35035 34125
rect 34977 34085 34989 34119
rect 35023 34116 35035 34119
rect 35342 34116 35348 34128
rect 35023 34088 35348 34116
rect 35023 34085 35035 34088
rect 34977 34079 35035 34085
rect 35342 34076 35348 34088
rect 35400 34116 35406 34128
rect 36446 34116 36452 34128
rect 35400 34088 36452 34116
rect 35400 34076 35406 34088
rect 36446 34076 36452 34088
rect 36504 34076 36510 34128
rect 38654 34076 38660 34128
rect 38712 34116 38718 34128
rect 38841 34119 38899 34125
rect 38841 34116 38853 34119
rect 38712 34088 38853 34116
rect 38712 34076 38718 34088
rect 38841 34085 38853 34088
rect 38887 34116 38899 34119
rect 39117 34119 39175 34125
rect 39117 34116 39129 34119
rect 38887 34088 39129 34116
rect 38887 34085 38899 34088
rect 38841 34079 38899 34085
rect 39117 34085 39129 34088
rect 39163 34085 39175 34119
rect 39117 34079 39175 34085
rect 40402 34076 40408 34128
rect 40460 34116 40466 34128
rect 40678 34116 40684 34128
rect 40460 34088 40684 34116
rect 40460 34076 40466 34088
rect 40678 34076 40684 34088
rect 40736 34076 40742 34128
rect 40862 34076 40868 34128
rect 40920 34116 40926 34128
rect 41156 34125 41184 34156
rect 42518 34144 42524 34156
rect 42576 34184 42582 34196
rect 44266 34184 44272 34196
rect 42576 34156 44272 34184
rect 42576 34144 42582 34156
rect 44266 34144 44272 34156
rect 44324 34144 44330 34196
rect 44542 34144 44548 34196
rect 44600 34184 44606 34196
rect 44637 34187 44695 34193
rect 44637 34184 44649 34187
rect 44600 34156 44649 34184
rect 44600 34144 44606 34156
rect 44637 34153 44649 34156
rect 44683 34153 44695 34187
rect 44637 34147 44695 34153
rect 41049 34119 41107 34125
rect 41049 34116 41061 34119
rect 40920 34088 41061 34116
rect 40920 34076 40926 34088
rect 41049 34085 41061 34088
rect 41095 34085 41107 34119
rect 41049 34079 41107 34085
rect 41141 34119 41199 34125
rect 41141 34085 41153 34119
rect 41187 34116 41199 34119
rect 41414 34116 41420 34128
rect 41187 34088 41420 34116
rect 41187 34085 41199 34088
rect 41141 34079 41199 34085
rect 41414 34076 41420 34088
rect 41472 34076 41478 34128
rect 43162 34116 43168 34128
rect 43123 34088 43168 34116
rect 43162 34076 43168 34088
rect 43220 34076 43226 34128
rect 43806 34116 43812 34128
rect 43767 34088 43812 34116
rect 43806 34076 43812 34088
rect 43864 34076 43870 34128
rect 32585 34051 32643 34057
rect 32585 34048 32597 34051
rect 32416 34020 32597 34048
rect 32585 34017 32597 34020
rect 32631 34017 32643 34051
rect 32585 34011 32643 34017
rect 33965 34051 34023 34057
rect 33965 34017 33977 34051
rect 34011 34048 34023 34051
rect 34606 34048 34612 34060
rect 34011 34020 34612 34048
rect 34011 34017 34023 34020
rect 33965 34011 34023 34017
rect 34606 34008 34612 34020
rect 34664 34008 34670 34060
rect 35713 34051 35771 34057
rect 35713 34017 35725 34051
rect 35759 34048 35771 34051
rect 36541 34051 36599 34057
rect 36541 34048 36553 34051
rect 35759 34020 36553 34048
rect 35759 34017 35771 34020
rect 35713 34011 35771 34017
rect 36541 34017 36553 34020
rect 36587 34048 36599 34051
rect 37001 34051 37059 34057
rect 37001 34048 37013 34051
rect 36587 34020 37013 34048
rect 36587 34017 36599 34020
rect 36541 34011 36599 34017
rect 37001 34017 37013 34020
rect 37047 34017 37059 34051
rect 37001 34011 37059 34017
rect 37458 34008 37464 34060
rect 37516 34048 37522 34060
rect 38105 34051 38163 34057
rect 38105 34048 38117 34051
rect 37516 34020 38117 34048
rect 37516 34008 37522 34020
rect 38105 34017 38117 34020
rect 38151 34048 38163 34051
rect 38470 34048 38476 34060
rect 38151 34020 38476 34048
rect 38151 34017 38163 34020
rect 38105 34011 38163 34017
rect 38470 34008 38476 34020
rect 38528 34008 38534 34060
rect 38562 34008 38568 34060
rect 38620 34048 38626 34060
rect 39850 34048 39856 34060
rect 38620 34020 38665 34048
rect 39811 34020 39856 34048
rect 38620 34008 38626 34020
rect 39850 34008 39856 34020
rect 39908 34008 39914 34060
rect 45370 34008 45376 34060
rect 45428 34048 45434 34060
rect 45592 34051 45650 34057
rect 45592 34048 45604 34051
rect 45428 34020 45604 34048
rect 45428 34008 45434 34020
rect 45592 34017 45604 34020
rect 45638 34017 45650 34051
rect 45592 34011 45650 34017
rect 24670 33980 24676 33992
rect 23446 33952 24676 33980
rect 24670 33940 24676 33952
rect 24728 33940 24734 33992
rect 24762 33940 24768 33992
rect 24820 33980 24826 33992
rect 24949 33983 25007 33989
rect 24949 33980 24961 33983
rect 24820 33952 24961 33980
rect 24820 33940 24826 33952
rect 24949 33949 24961 33952
rect 24995 33949 25007 33983
rect 24949 33943 25007 33949
rect 26605 33983 26663 33989
rect 26605 33949 26617 33983
rect 26651 33980 26663 33983
rect 26694 33980 26700 33992
rect 26651 33952 26700 33980
rect 26651 33949 26663 33952
rect 26605 33943 26663 33949
rect 26694 33940 26700 33952
rect 26752 33940 26758 33992
rect 26878 33980 26884 33992
rect 26839 33952 26884 33980
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 28166 33980 28172 33992
rect 28127 33952 28172 33980
rect 28166 33940 28172 33952
rect 28224 33940 28230 33992
rect 29549 33983 29607 33989
rect 29549 33949 29561 33983
rect 29595 33980 29607 33983
rect 29733 33983 29791 33989
rect 29733 33980 29745 33983
rect 29595 33952 29745 33980
rect 29595 33949 29607 33952
rect 29549 33943 29607 33949
rect 29733 33949 29745 33952
rect 29779 33980 29791 33983
rect 31202 33980 31208 33992
rect 29779 33952 31208 33980
rect 29779 33949 29791 33952
rect 29733 33943 29791 33949
rect 31202 33940 31208 33952
rect 31260 33940 31266 33992
rect 33870 33980 33876 33992
rect 33783 33952 33876 33980
rect 33870 33940 33876 33952
rect 33928 33980 33934 33992
rect 33928 33952 35106 33980
rect 33928 33940 33934 33952
rect 28721 33915 28779 33921
rect 28721 33881 28733 33915
rect 28767 33912 28779 33915
rect 29086 33912 29092 33924
rect 28767 33884 29092 33912
rect 28767 33881 28779 33884
rect 28721 33875 28779 33881
rect 29086 33872 29092 33884
rect 29144 33912 29150 33924
rect 30285 33915 30343 33921
rect 30285 33912 30297 33915
rect 29144 33884 30297 33912
rect 29144 33872 29150 33884
rect 30285 33881 30297 33884
rect 30331 33881 30343 33915
rect 30285 33875 30343 33881
rect 32950 33872 32956 33924
rect 33008 33912 33014 33924
rect 33505 33915 33563 33921
rect 33505 33912 33517 33915
rect 33008 33884 33517 33912
rect 33008 33872 33014 33884
rect 33505 33881 33517 33884
rect 33551 33912 33563 33915
rect 34698 33912 34704 33924
rect 33551 33884 34704 33912
rect 33551 33881 33563 33884
rect 33505 33875 33563 33881
rect 34698 33872 34704 33884
rect 34756 33872 34762 33924
rect 19794 33804 19800 33856
rect 19852 33844 19858 33856
rect 21453 33847 21511 33853
rect 21453 33844 21465 33847
rect 19852 33816 21465 33844
rect 19852 33804 19858 33816
rect 21453 33813 21465 33816
rect 21499 33844 21511 33847
rect 21910 33844 21916 33856
rect 21499 33816 21916 33844
rect 21499 33813 21511 33816
rect 21453 33807 21511 33813
rect 21910 33804 21916 33816
rect 21968 33804 21974 33856
rect 27522 33844 27528 33856
rect 27483 33816 27528 33844
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 31110 33844 31116 33856
rect 31071 33816 31116 33844
rect 31110 33804 31116 33816
rect 31168 33804 31174 33856
rect 31849 33847 31907 33853
rect 31849 33813 31861 33847
rect 31895 33844 31907 33847
rect 32398 33844 32404 33856
rect 31895 33816 32404 33844
rect 31895 33813 31907 33816
rect 31849 33807 31907 33813
rect 32398 33804 32404 33816
rect 32456 33804 32462 33856
rect 34146 33844 34152 33856
rect 34107 33816 34152 33844
rect 34146 33804 34152 33816
rect 34204 33804 34210 33856
rect 35078 33844 35106 33952
rect 35158 33940 35164 33992
rect 35216 33980 35222 33992
rect 35345 33983 35403 33989
rect 35345 33980 35357 33983
rect 35216 33952 35357 33980
rect 35216 33940 35222 33952
rect 35345 33949 35357 33952
rect 35391 33980 35403 33983
rect 35802 33980 35808 33992
rect 35391 33952 35808 33980
rect 35391 33949 35403 33952
rect 35345 33943 35403 33949
rect 35802 33940 35808 33952
rect 35860 33940 35866 33992
rect 41506 33980 41512 33992
rect 41467 33952 41512 33980
rect 41506 33940 41512 33952
rect 41564 33940 41570 33992
rect 43717 33983 43775 33989
rect 43717 33949 43729 33983
rect 43763 33980 43775 33983
rect 44082 33980 44088 33992
rect 43763 33952 44088 33980
rect 43763 33949 43775 33952
rect 43717 33943 43775 33949
rect 44082 33940 44088 33952
rect 44140 33980 44146 33992
rect 45094 33980 45100 33992
rect 44140 33952 45100 33980
rect 44140 33940 44146 33952
rect 45094 33940 45100 33952
rect 45152 33940 45158 33992
rect 35250 33912 35256 33924
rect 35211 33884 35256 33912
rect 35250 33872 35256 33884
rect 35308 33912 35314 33924
rect 35989 33915 36047 33921
rect 35989 33912 36001 33915
rect 35308 33884 36001 33912
rect 35308 33872 35314 33884
rect 35989 33881 36001 33884
rect 36035 33912 36047 33915
rect 36357 33915 36415 33921
rect 36357 33912 36369 33915
rect 36035 33884 36369 33912
rect 36035 33881 36047 33884
rect 35989 33875 36047 33881
rect 36357 33881 36369 33884
rect 36403 33912 36415 33915
rect 36722 33912 36728 33924
rect 36403 33884 36728 33912
rect 36403 33881 36415 33884
rect 36357 33875 36415 33881
rect 36722 33872 36728 33884
rect 36780 33872 36786 33924
rect 43162 33872 43168 33924
rect 43220 33912 43226 33924
rect 44269 33915 44327 33921
rect 44269 33912 44281 33915
rect 43220 33884 44281 33912
rect 43220 33872 43226 33884
rect 44269 33881 44281 33884
rect 44315 33881 44327 33915
rect 44269 33875 44327 33881
rect 35142 33847 35200 33853
rect 35142 33844 35154 33847
rect 35078 33816 35154 33844
rect 35142 33813 35154 33816
rect 35188 33844 35200 33847
rect 35618 33844 35624 33856
rect 35188 33816 35624 33844
rect 35188 33813 35200 33816
rect 35142 33807 35200 33813
rect 35618 33804 35624 33816
rect 35676 33804 35682 33856
rect 40083 33847 40141 33853
rect 40083 33813 40095 33847
rect 40129 33844 40141 33847
rect 40494 33844 40500 33856
rect 40129 33816 40500 33844
rect 40129 33813 40141 33816
rect 40083 33807 40141 33813
rect 40494 33804 40500 33816
rect 40552 33804 40558 33856
rect 43622 33804 43628 33856
rect 43680 33844 43686 33856
rect 44818 33844 44824 33856
rect 43680 33816 44824 33844
rect 43680 33804 43686 33816
rect 44818 33804 44824 33816
rect 44876 33804 44882 33856
rect 45695 33847 45753 33853
rect 45695 33813 45707 33847
rect 45741 33844 45753 33847
rect 46014 33844 46020 33856
rect 45741 33816 46020 33844
rect 45741 33813 45753 33816
rect 45695 33807 45753 33813
rect 46014 33804 46020 33816
rect 46072 33804 46078 33856
rect 1104 33754 48852 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 48852 33754
rect 1104 33680 48852 33702
rect 14642 33600 14648 33652
rect 14700 33640 14706 33652
rect 16301 33643 16359 33649
rect 16301 33640 16313 33643
rect 14700 33612 16313 33640
rect 14700 33600 14706 33612
rect 16301 33609 16313 33612
rect 16347 33640 16359 33643
rect 16390 33640 16396 33652
rect 16347 33612 16396 33640
rect 16347 33609 16359 33612
rect 16301 33603 16359 33609
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 17494 33640 17500 33652
rect 17455 33612 17500 33640
rect 17494 33600 17500 33612
rect 17552 33600 17558 33652
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 19797 33643 19855 33649
rect 19797 33640 19809 33643
rect 19484 33612 19809 33640
rect 19484 33600 19490 33612
rect 19797 33609 19809 33612
rect 19843 33640 19855 33643
rect 20162 33640 20168 33652
rect 19843 33612 20168 33640
rect 19843 33609 19855 33612
rect 19797 33603 19855 33609
rect 20162 33600 20168 33612
rect 20220 33600 20226 33652
rect 22738 33640 22744 33652
rect 22699 33612 22744 33640
rect 22738 33600 22744 33612
rect 22796 33600 22802 33652
rect 23198 33640 23204 33652
rect 23159 33612 23204 33640
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 24670 33600 24676 33652
rect 24728 33640 24734 33652
rect 25409 33643 25467 33649
rect 25409 33640 25421 33643
rect 24728 33612 25421 33640
rect 24728 33600 24734 33612
rect 25409 33609 25421 33612
rect 25455 33609 25467 33643
rect 25409 33603 25467 33609
rect 25731 33643 25789 33649
rect 25731 33609 25743 33643
rect 25777 33640 25789 33643
rect 25866 33640 25872 33652
rect 25777 33612 25872 33640
rect 25777 33609 25789 33612
rect 25731 33603 25789 33609
rect 25866 33600 25872 33612
rect 25924 33600 25930 33652
rect 28166 33640 28172 33652
rect 28127 33612 28172 33640
rect 28166 33600 28172 33612
rect 28224 33600 28230 33652
rect 31294 33640 31300 33652
rect 28276 33612 30880 33640
rect 31255 33612 31300 33640
rect 13814 33532 13820 33584
rect 13872 33572 13878 33584
rect 15105 33575 15163 33581
rect 15105 33572 15117 33575
rect 13872 33544 15117 33572
rect 13872 33532 13878 33544
rect 15105 33541 15117 33544
rect 15151 33541 15163 33575
rect 20180 33572 20208 33600
rect 24578 33572 24584 33584
rect 20180 33544 24584 33572
rect 15105 33535 15163 33541
rect 15120 33504 15148 33535
rect 24578 33532 24584 33544
rect 24636 33532 24642 33584
rect 24854 33532 24860 33584
rect 24912 33572 24918 33584
rect 28276 33572 28304 33612
rect 24912 33544 28304 33572
rect 24912 33532 24918 33544
rect 29638 33532 29644 33584
rect 29696 33572 29702 33584
rect 30653 33575 30711 33581
rect 30653 33572 30665 33575
rect 29696 33544 30665 33572
rect 29696 33532 29702 33544
rect 30653 33541 30665 33544
rect 30699 33541 30711 33575
rect 30852 33572 30880 33612
rect 31294 33600 31300 33612
rect 31352 33640 31358 33652
rect 31895 33643 31953 33649
rect 31895 33640 31907 33643
rect 31352 33612 31907 33640
rect 31352 33600 31358 33612
rect 31895 33609 31907 33612
rect 31941 33609 31953 33643
rect 31895 33603 31953 33609
rect 32033 33643 32091 33649
rect 32033 33609 32045 33643
rect 32079 33640 32091 33643
rect 32398 33640 32404 33652
rect 32079 33612 32404 33640
rect 32079 33609 32091 33612
rect 32033 33603 32091 33609
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 35161 33643 35219 33649
rect 35161 33609 35173 33643
rect 35207 33640 35219 33643
rect 35250 33640 35256 33652
rect 35207 33612 35256 33640
rect 35207 33609 35219 33612
rect 35161 33603 35219 33609
rect 35250 33600 35256 33612
rect 35308 33600 35314 33652
rect 35526 33640 35532 33652
rect 35487 33612 35532 33640
rect 35526 33600 35532 33612
rect 35584 33600 35590 33652
rect 36354 33600 36360 33652
rect 36412 33640 36418 33652
rect 36587 33643 36645 33649
rect 36587 33640 36599 33643
rect 36412 33612 36599 33640
rect 36412 33600 36418 33612
rect 36587 33609 36599 33612
rect 36633 33609 36645 33643
rect 36722 33640 36728 33652
rect 36683 33612 36728 33640
rect 36587 33603 36645 33609
rect 36722 33600 36728 33612
rect 36780 33600 36786 33652
rect 36906 33640 36912 33652
rect 36867 33612 36912 33640
rect 36906 33600 36912 33612
rect 36964 33600 36970 33652
rect 38470 33640 38476 33652
rect 38431 33612 38476 33640
rect 38470 33600 38476 33612
rect 38528 33600 38534 33652
rect 39945 33643 40003 33649
rect 39945 33609 39957 33643
rect 39991 33640 40003 33643
rect 40034 33640 40040 33652
rect 39991 33612 40040 33640
rect 39991 33609 40003 33612
rect 39945 33603 40003 33609
rect 40034 33600 40040 33612
rect 40092 33600 40098 33652
rect 40862 33600 40868 33652
rect 40920 33640 40926 33652
rect 42613 33643 42671 33649
rect 42613 33640 42625 33643
rect 40920 33612 42625 33640
rect 40920 33600 40926 33612
rect 42613 33609 42625 33612
rect 42659 33609 42671 33643
rect 43717 33643 43775 33649
rect 43717 33640 43729 33643
rect 42613 33603 42671 33609
rect 42766 33612 43729 33640
rect 32217 33575 32275 33581
rect 32217 33572 32229 33575
rect 30852 33544 32229 33572
rect 30653 33535 30711 33541
rect 32217 33541 32229 33544
rect 32263 33541 32275 33575
rect 32217 33535 32275 33541
rect 35050 33575 35108 33581
rect 35050 33541 35062 33575
rect 35096 33572 35108 33575
rect 35618 33572 35624 33584
rect 35096 33544 35624 33572
rect 35096 33541 35108 33544
rect 35050 33535 35108 33541
rect 35618 33532 35624 33544
rect 35676 33572 35682 33584
rect 37461 33575 37519 33581
rect 37461 33572 37473 33575
rect 35676 33544 37473 33572
rect 35676 33532 35682 33544
rect 37461 33541 37473 33544
rect 37507 33541 37519 33575
rect 37461 33535 37519 33541
rect 37921 33575 37979 33581
rect 37921 33541 37933 33575
rect 37967 33572 37979 33575
rect 38562 33572 38568 33584
rect 37967 33544 38568 33572
rect 37967 33541 37979 33544
rect 37921 33535 37979 33541
rect 38562 33532 38568 33544
rect 38620 33532 38626 33584
rect 39390 33532 39396 33584
rect 39448 33572 39454 33584
rect 41230 33572 41236 33584
rect 39448 33544 40356 33572
rect 41191 33544 41236 33572
rect 39448 33532 39454 33544
rect 16022 33504 16028 33516
rect 15120 33476 15792 33504
rect 15935 33476 16028 33504
rect 14328 33439 14386 33445
rect 14328 33405 14340 33439
rect 14374 33436 14386 33439
rect 14415 33439 14473 33445
rect 14374 33405 14387 33436
rect 14328 33399 14387 33405
rect 14415 33405 14427 33439
rect 14461 33436 14473 33439
rect 14734 33436 14740 33448
rect 14461 33408 14740 33436
rect 14461 33405 14473 33408
rect 14415 33399 14473 33405
rect 14359 33368 14387 33399
rect 14734 33396 14740 33408
rect 14792 33396 14798 33448
rect 15286 33396 15292 33448
rect 15344 33436 15350 33448
rect 15565 33439 15623 33445
rect 15565 33436 15577 33439
rect 15344 33408 15577 33436
rect 15344 33396 15350 33408
rect 15565 33405 15577 33408
rect 15611 33436 15623 33439
rect 15654 33436 15660 33448
rect 15611 33408 15660 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 15654 33396 15660 33408
rect 15712 33396 15718 33448
rect 15764 33445 15792 33476
rect 16022 33464 16028 33476
rect 16080 33504 16086 33516
rect 16669 33507 16727 33513
rect 16669 33504 16681 33507
rect 16080 33476 16681 33504
rect 16080 33464 16086 33476
rect 16669 33473 16681 33476
rect 16715 33473 16727 33507
rect 18046 33504 18052 33516
rect 16669 33467 16727 33473
rect 16776 33476 18052 33504
rect 15749 33439 15807 33445
rect 15749 33405 15761 33439
rect 15795 33405 15807 33439
rect 15749 33399 15807 33405
rect 14829 33371 14887 33377
rect 14829 33368 14841 33371
rect 14359 33340 14841 33368
rect 14829 33337 14841 33340
rect 14875 33368 14887 33371
rect 16776 33368 16804 33476
rect 18046 33464 18052 33476
rect 18104 33464 18110 33516
rect 19429 33507 19487 33513
rect 19429 33473 19441 33507
rect 19475 33504 19487 33507
rect 20070 33504 20076 33516
rect 19475 33476 20076 33504
rect 19475 33473 19487 33476
rect 19429 33467 19487 33473
rect 20070 33464 20076 33476
rect 20128 33464 20134 33516
rect 24118 33504 24124 33516
rect 24079 33476 24124 33504
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24762 33504 24768 33516
rect 24723 33476 24768 33504
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 26786 33504 26792 33516
rect 26699 33476 26792 33504
rect 26786 33464 26792 33476
rect 26844 33504 26850 33516
rect 27522 33504 27528 33516
rect 26844 33476 27528 33504
rect 26844 33464 26850 33476
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 31110 33464 31116 33516
rect 31168 33504 31174 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31168 33476 32137 33504
rect 31168 33464 31174 33476
rect 32125 33473 32137 33476
rect 32171 33504 32183 33507
rect 32306 33504 32312 33516
rect 32171 33476 32312 33504
rect 32171 33473 32183 33476
rect 32125 33467 32183 33473
rect 32306 33464 32312 33476
rect 32364 33464 32370 33516
rect 35253 33507 35311 33513
rect 35253 33473 35265 33507
rect 35299 33504 35311 33507
rect 35802 33504 35808 33516
rect 35299 33476 35808 33504
rect 35299 33473 35311 33476
rect 35253 33467 35311 33473
rect 35802 33464 35808 33476
rect 35860 33504 35866 33516
rect 35989 33507 36047 33513
rect 35989 33504 36001 33507
rect 35860 33476 36001 33504
rect 35860 33464 35866 33476
rect 35989 33473 36001 33476
rect 36035 33504 36047 33507
rect 36357 33507 36415 33513
rect 36357 33504 36369 33507
rect 36035 33476 36369 33504
rect 36035 33473 36047 33476
rect 35989 33467 36047 33473
rect 36357 33473 36369 33476
rect 36403 33504 36415 33507
rect 36814 33504 36820 33516
rect 36403 33476 36820 33504
rect 36403 33473 36415 33476
rect 36357 33467 36415 33473
rect 36814 33464 36820 33476
rect 36872 33464 36878 33516
rect 39206 33464 39212 33516
rect 39264 33504 39270 33516
rect 39850 33504 39856 33516
rect 39264 33476 39856 33504
rect 39264 33464 39270 33476
rect 39850 33464 39856 33476
rect 39908 33504 39914 33516
rect 40221 33507 40279 33513
rect 40221 33504 40233 33507
rect 39908 33476 40233 33504
rect 39908 33464 39914 33476
rect 40221 33473 40233 33476
rect 40267 33473 40279 33507
rect 40221 33467 40279 33473
rect 17012 33439 17070 33445
rect 17012 33405 17024 33439
rect 17058 33436 17070 33439
rect 17494 33436 17500 33448
rect 17058 33408 17500 33436
rect 17058 33405 17070 33408
rect 17012 33399 17070 33405
rect 17494 33396 17500 33408
rect 17552 33396 17558 33448
rect 18598 33436 18604 33448
rect 18559 33408 18604 33436
rect 18598 33396 18604 33408
rect 18656 33396 18662 33448
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33436 18843 33439
rect 19794 33436 19800 33448
rect 18831 33408 19800 33436
rect 18831 33405 18843 33408
rect 18785 33399 18843 33405
rect 14875 33340 16804 33368
rect 14875 33337 14887 33340
rect 14829 33331 14887 33337
rect 16850 33328 16856 33380
rect 16908 33368 16914 33380
rect 17773 33371 17831 33377
rect 17773 33368 17785 33371
rect 16908 33340 17785 33368
rect 16908 33328 16914 33340
rect 17773 33337 17785 33340
rect 17819 33368 17831 33371
rect 18800 33368 18828 33399
rect 19794 33396 19800 33408
rect 19852 33396 19858 33448
rect 21269 33439 21327 33445
rect 21269 33405 21281 33439
rect 21315 33436 21327 33439
rect 21729 33439 21787 33445
rect 21729 33436 21741 33439
rect 21315 33408 21741 33436
rect 21315 33405 21327 33408
rect 21269 33399 21327 33405
rect 21729 33405 21741 33408
rect 21775 33405 21787 33439
rect 21910 33436 21916 33448
rect 21871 33408 21916 33436
rect 21729 33399 21787 33405
rect 19058 33368 19064 33380
rect 17819 33340 18828 33368
rect 19019 33340 19064 33368
rect 17819 33337 17831 33340
rect 17773 33331 17831 33337
rect 19058 33328 19064 33340
rect 19116 33328 19122 33380
rect 19981 33371 20039 33377
rect 19981 33337 19993 33371
rect 20027 33337 20039 33371
rect 19981 33331 20039 33337
rect 17083 33303 17141 33309
rect 17083 33269 17095 33303
rect 17129 33300 17141 33303
rect 17310 33300 17316 33312
rect 17129 33272 17316 33300
rect 17129 33269 17141 33272
rect 17083 33263 17141 33269
rect 17310 33260 17316 33272
rect 17368 33260 17374 33312
rect 19996 33300 20024 33331
rect 20070 33328 20076 33380
rect 20128 33368 20134 33380
rect 20625 33371 20683 33377
rect 20128 33340 20173 33368
rect 20128 33328 20134 33340
rect 20625 33337 20637 33371
rect 20671 33368 20683 33371
rect 21358 33368 21364 33380
rect 20671 33340 21364 33368
rect 20671 33337 20683 33340
rect 20625 33331 20683 33337
rect 21358 33328 21364 33340
rect 21416 33328 21422 33380
rect 21744 33368 21772 33399
rect 21910 33396 21916 33408
rect 21968 33436 21974 33448
rect 22370 33436 22376 33448
rect 21968 33408 22376 33436
rect 21968 33396 21974 33408
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 25660 33439 25718 33445
rect 25660 33405 25672 33439
rect 25706 33436 25718 33439
rect 26050 33436 26056 33448
rect 25706 33408 26056 33436
rect 25706 33405 25718 33408
rect 25660 33399 25718 33405
rect 26050 33396 26056 33408
rect 26108 33396 26114 33448
rect 29089 33439 29147 33445
rect 29089 33405 29101 33439
rect 29135 33436 29147 33439
rect 29730 33436 29736 33448
rect 29135 33408 29736 33436
rect 29135 33405 29147 33408
rect 29089 33399 29147 33405
rect 29730 33396 29736 33408
rect 29788 33396 29794 33448
rect 31386 33396 31392 33448
rect 31444 33436 31450 33448
rect 32214 33436 32220 33448
rect 31444 33408 32220 33436
rect 31444 33396 31450 33408
rect 32214 33396 32220 33408
rect 32272 33436 32278 33448
rect 32769 33439 32827 33445
rect 32769 33436 32781 33439
rect 32272 33408 32781 33436
rect 32272 33396 32278 33408
rect 32769 33405 32781 33408
rect 32815 33405 32827 33439
rect 32769 33399 32827 33405
rect 33597 33439 33655 33445
rect 33597 33405 33609 33439
rect 33643 33436 33655 33439
rect 34241 33439 34299 33445
rect 34241 33436 34253 33439
rect 33643 33408 34253 33436
rect 33643 33405 33655 33408
rect 33597 33399 33655 33405
rect 34241 33405 34253 33408
rect 34287 33436 34299 33439
rect 34330 33436 34336 33448
rect 34287 33408 34336 33436
rect 34287 33405 34299 33408
rect 34241 33399 34299 33405
rect 34330 33396 34336 33408
rect 34388 33396 34394 33448
rect 37274 33396 37280 33448
rect 37332 33436 37338 33448
rect 38013 33439 38071 33445
rect 38013 33436 38025 33439
rect 37332 33408 38025 33436
rect 37332 33396 37338 33408
rect 38013 33405 38025 33408
rect 38059 33436 38071 33439
rect 38841 33439 38899 33445
rect 38841 33436 38853 33439
rect 38059 33408 38853 33436
rect 38059 33405 38071 33408
rect 38013 33399 38071 33405
rect 38841 33405 38853 33408
rect 38887 33405 38899 33439
rect 38841 33399 38899 33405
rect 39444 33439 39502 33445
rect 39444 33405 39456 33439
rect 39490 33436 39502 33439
rect 40034 33436 40040 33448
rect 39490 33408 40040 33436
rect 39490 33405 39502 33408
rect 39444 33399 39502 33405
rect 40034 33396 40040 33408
rect 40092 33396 40098 33448
rect 40328 33436 40356 33544
rect 41230 33532 41236 33544
rect 41288 33532 41294 33584
rect 41414 33532 41420 33584
rect 41472 33572 41478 33584
rect 41509 33575 41567 33581
rect 41509 33572 41521 33575
rect 41472 33544 41521 33572
rect 41472 33532 41478 33544
rect 41509 33541 41521 33544
rect 41555 33572 41567 33575
rect 42766 33572 42794 33612
rect 43717 33609 43729 33612
rect 43763 33640 43775 33643
rect 43806 33640 43812 33652
rect 43763 33612 43812 33640
rect 43763 33609 43775 33612
rect 43717 33603 43775 33609
rect 43806 33600 43812 33612
rect 43864 33600 43870 33652
rect 44082 33640 44088 33652
rect 44043 33612 44088 33640
rect 44082 33600 44088 33612
rect 44140 33600 44146 33652
rect 45002 33640 45008 33652
rect 44963 33612 45008 33640
rect 45002 33600 45008 33612
rect 45060 33600 45066 33652
rect 45370 33600 45376 33652
rect 45428 33640 45434 33652
rect 45557 33643 45615 33649
rect 45557 33640 45569 33643
rect 45428 33612 45569 33640
rect 45428 33600 45434 33612
rect 45557 33609 45569 33612
rect 45603 33609 45615 33643
rect 45557 33603 45615 33609
rect 41555 33544 42794 33572
rect 41555 33541 41567 33544
rect 41509 33535 41567 33541
rect 40748 33439 40806 33445
rect 40748 33436 40760 33439
rect 40328 33408 40760 33436
rect 40748 33405 40760 33408
rect 40794 33436 40806 33439
rect 41248 33436 41276 33532
rect 46934 33504 46940 33516
rect 43272 33476 46940 33504
rect 40794 33408 41276 33436
rect 41852 33439 41910 33445
rect 40794 33405 40806 33408
rect 40748 33399 40806 33405
rect 41852 33405 41864 33439
rect 41898 33405 41910 33439
rect 41852 33399 41910 33405
rect 42864 33439 42922 33445
rect 42864 33405 42876 33439
rect 42910 33436 42922 33439
rect 42978 33436 42984 33448
rect 42910 33408 42984 33436
rect 42910 33405 42922 33408
rect 42864 33399 42922 33405
rect 22002 33368 22008 33380
rect 21744 33340 22008 33368
rect 22002 33328 22008 33340
rect 22060 33368 22066 33380
rect 22830 33368 22836 33380
rect 22060 33340 22836 33368
rect 22060 33328 22066 33340
rect 22830 33328 22836 33340
rect 22888 33328 22894 33380
rect 23937 33371 23995 33377
rect 23937 33337 23949 33371
rect 23983 33368 23995 33371
rect 24118 33368 24124 33380
rect 23983 33340 24124 33368
rect 23983 33337 23995 33340
rect 23937 33331 23995 33337
rect 24118 33328 24124 33340
rect 24176 33368 24182 33380
rect 24213 33371 24271 33377
rect 24213 33368 24225 33371
rect 24176 33340 24225 33368
rect 24176 33328 24182 33340
rect 24213 33337 24225 33340
rect 24259 33368 24271 33371
rect 26513 33371 26571 33377
rect 26513 33368 26525 33371
rect 24259 33340 26525 33368
rect 24259 33337 24271 33340
rect 24213 33331 24271 33337
rect 26513 33337 26525 33340
rect 26559 33368 26571 33371
rect 26602 33368 26608 33380
rect 26559 33340 26608 33368
rect 26559 33337 26571 33340
rect 26513 33331 26571 33337
rect 26602 33328 26608 33340
rect 26660 33368 26666 33380
rect 26881 33371 26939 33377
rect 26881 33368 26893 33371
rect 26660 33340 26893 33368
rect 26660 33328 26666 33340
rect 26881 33337 26893 33340
rect 26927 33337 26939 33371
rect 27430 33368 27436 33380
rect 27391 33340 27436 33368
rect 26881 33331 26939 33337
rect 20254 33300 20260 33312
rect 19996 33272 20260 33300
rect 20254 33260 20260 33272
rect 20312 33260 20318 33312
rect 20714 33260 20720 33312
rect 20772 33300 20778 33312
rect 20901 33303 20959 33309
rect 20901 33300 20913 33303
rect 20772 33272 20913 33300
rect 20772 33260 20778 33272
rect 20901 33269 20913 33272
rect 20947 33269 20959 33303
rect 21726 33300 21732 33312
rect 21687 33272 21732 33300
rect 20901 33263 20959 33269
rect 21726 33260 21732 33272
rect 21784 33260 21790 33312
rect 25130 33300 25136 33312
rect 25091 33272 25136 33300
rect 25130 33260 25136 33272
rect 25188 33260 25194 33312
rect 26896 33300 26924 33331
rect 27430 33328 27436 33340
rect 27488 33328 27494 33380
rect 29641 33371 29699 33377
rect 29641 33337 29653 33371
rect 29687 33368 29699 33371
rect 29822 33368 29828 33380
rect 29687 33340 29828 33368
rect 29687 33337 29699 33340
rect 29641 33331 29699 33337
rect 29822 33328 29828 33340
rect 29880 33368 29886 33380
rect 30095 33371 30153 33377
rect 30095 33368 30107 33371
rect 29880 33340 30107 33368
rect 29880 33328 29886 33340
rect 30095 33337 30107 33340
rect 30141 33368 30153 33371
rect 30466 33368 30472 33380
rect 30141 33340 30472 33368
rect 30141 33337 30153 33340
rect 30095 33331 30153 33337
rect 30466 33328 30472 33340
rect 30524 33328 30530 33380
rect 31665 33371 31723 33377
rect 31665 33337 31677 33371
rect 31711 33368 31723 33371
rect 31754 33368 31760 33380
rect 31711 33340 31760 33368
rect 31711 33337 31723 33340
rect 31665 33331 31723 33337
rect 31754 33328 31760 33340
rect 31812 33328 31818 33380
rect 33321 33371 33379 33377
rect 33321 33337 33333 33371
rect 33367 33368 33379 33371
rect 33413 33371 33471 33377
rect 33413 33368 33425 33371
rect 33367 33340 33425 33368
rect 33367 33337 33379 33340
rect 33321 33331 33379 33337
rect 33413 33337 33425 33340
rect 33459 33337 33471 33371
rect 33962 33368 33968 33380
rect 33923 33340 33968 33368
rect 33413 33331 33471 33337
rect 27709 33303 27767 33309
rect 27709 33300 27721 33303
rect 26896 33272 27721 33300
rect 27709 33269 27721 33272
rect 27755 33300 27767 33303
rect 28445 33303 28503 33309
rect 28445 33300 28457 33303
rect 27755 33272 28457 33300
rect 27755 33269 27767 33272
rect 27709 33263 27767 33269
rect 28445 33269 28457 33272
rect 28491 33269 28503 33303
rect 33428 33300 33456 33331
rect 33962 33328 33968 33340
rect 34020 33328 34026 33380
rect 34606 33368 34612 33380
rect 34567 33340 34612 33368
rect 34606 33328 34612 33340
rect 34664 33328 34670 33380
rect 34698 33328 34704 33380
rect 34756 33368 34762 33380
rect 34885 33371 34943 33377
rect 34885 33368 34897 33371
rect 34756 33340 34897 33368
rect 34756 33328 34762 33340
rect 34885 33337 34897 33340
rect 34931 33368 34943 33371
rect 35250 33368 35256 33380
rect 34931 33340 35256 33368
rect 34931 33337 34943 33340
rect 34885 33331 34943 33337
rect 35250 33328 35256 33340
rect 35308 33328 35314 33380
rect 36446 33368 36452 33380
rect 36407 33340 36452 33368
rect 36446 33328 36452 33340
rect 36504 33328 36510 33380
rect 39531 33371 39589 33377
rect 39531 33337 39543 33371
rect 39577 33368 39589 33371
rect 40586 33368 40592 33380
rect 39577 33340 40592 33368
rect 39577 33337 39589 33340
rect 39531 33331 39589 33337
rect 40586 33328 40592 33340
rect 40644 33328 40650 33380
rect 41867 33368 41895 33399
rect 42978 33396 42984 33408
rect 43036 33436 43042 33448
rect 43272 33445 43300 33476
rect 46934 33464 46940 33476
rect 46992 33464 46998 33516
rect 43257 33439 43315 33445
rect 43257 33436 43269 33439
rect 43036 33408 43269 33436
rect 43036 33396 43042 33408
rect 43257 33405 43269 33408
rect 43303 33405 43315 33439
rect 43257 33399 43315 33405
rect 44520 33439 44578 33445
rect 44520 33405 44532 33439
rect 44566 33436 44578 33439
rect 45002 33436 45008 33448
rect 44566 33408 45008 33436
rect 44566 33405 44578 33408
rect 44520 33399 44578 33405
rect 45002 33396 45008 33408
rect 45060 33396 45066 33448
rect 42337 33371 42395 33377
rect 42337 33368 42349 33371
rect 41867 33340 42349 33368
rect 42337 33337 42349 33340
rect 42383 33368 42395 33371
rect 43622 33368 43628 33380
rect 42383 33340 43628 33368
rect 42383 33337 42395 33340
rect 42337 33331 42395 33337
rect 43622 33328 43628 33340
rect 43680 33328 43686 33380
rect 34624 33300 34652 33328
rect 38194 33300 38200 33312
rect 33428 33272 34652 33300
rect 38155 33272 38200 33300
rect 28445 33263 28503 33269
rect 38194 33260 38200 33272
rect 38252 33260 38258 33312
rect 40819 33303 40877 33309
rect 40819 33269 40831 33303
rect 40865 33300 40877 33303
rect 40954 33300 40960 33312
rect 40865 33272 40960 33300
rect 40865 33269 40877 33272
rect 40819 33263 40877 33269
rect 40954 33260 40960 33272
rect 41012 33260 41018 33312
rect 41923 33303 41981 33309
rect 41923 33269 41935 33303
rect 41969 33300 41981 33303
rect 42150 33300 42156 33312
rect 41969 33272 42156 33300
rect 41969 33269 41981 33272
rect 41923 33263 41981 33269
rect 42150 33260 42156 33272
rect 42208 33260 42214 33312
rect 42935 33303 42993 33309
rect 42935 33269 42947 33303
rect 42981 33300 42993 33303
rect 43162 33300 43168 33312
rect 42981 33272 43168 33300
rect 42981 33269 42993 33272
rect 42935 33263 42993 33269
rect 43162 33260 43168 33272
rect 43220 33260 43226 33312
rect 44591 33303 44649 33309
rect 44591 33269 44603 33303
rect 44637 33300 44649 33303
rect 44726 33300 44732 33312
rect 44637 33272 44732 33300
rect 44637 33269 44649 33272
rect 44591 33263 44649 33269
rect 44726 33260 44732 33272
rect 44784 33260 44790 33312
rect 1104 33210 48852 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 48852 33210
rect 1104 33136 48852 33158
rect 17954 33096 17960 33108
rect 17915 33068 17960 33096
rect 17954 33056 17960 33068
rect 18012 33056 18018 33108
rect 20806 33056 20812 33108
rect 20864 33096 20870 33108
rect 22646 33096 22652 33108
rect 20864 33068 22652 33096
rect 20864 33056 20870 33068
rect 22646 33056 22652 33068
rect 22704 33056 22710 33108
rect 23569 33099 23627 33105
rect 23569 33096 23581 33099
rect 23446 33068 23581 33096
rect 13814 32988 13820 33040
rect 13872 33028 13878 33040
rect 15378 33028 15384 33040
rect 13872 33000 15384 33028
rect 13872 32988 13878 33000
rect 15378 32988 15384 33000
rect 15436 32988 15442 33040
rect 15473 33031 15531 33037
rect 15473 32997 15485 33031
rect 15519 33028 15531 33031
rect 15562 33028 15568 33040
rect 15519 33000 15568 33028
rect 15519 32997 15531 33000
rect 15473 32991 15531 32997
rect 15562 32988 15568 33000
rect 15620 32988 15626 33040
rect 17218 33028 17224 33040
rect 17052 33000 17224 33028
rect 13630 32960 13636 32972
rect 13591 32932 13636 32960
rect 13630 32920 13636 32932
rect 13688 32920 13694 32972
rect 13906 32920 13912 32972
rect 13964 32960 13970 32972
rect 17052 32969 17080 33000
rect 17218 32988 17224 33000
rect 17276 32988 17282 33040
rect 19334 33028 19340 33040
rect 19295 33000 19340 33028
rect 19334 32988 19340 33000
rect 19392 32988 19398 33040
rect 21082 33028 21088 33040
rect 21043 33000 21088 33028
rect 21082 32988 21088 33000
rect 21140 32988 21146 33040
rect 23106 32988 23112 33040
rect 23164 33028 23170 33040
rect 23446 33028 23474 33068
rect 23569 33065 23581 33068
rect 23615 33065 23627 33099
rect 24118 33096 24124 33108
rect 24079 33068 24124 33096
rect 23569 33059 23627 33065
rect 24118 33056 24124 33068
rect 24176 33056 24182 33108
rect 26329 33099 26387 33105
rect 26329 33065 26341 33099
rect 26375 33096 26387 33099
rect 26602 33096 26608 33108
rect 26375 33068 26608 33096
rect 26375 33065 26387 33068
rect 26329 33059 26387 33065
rect 26602 33056 26608 33068
rect 26660 33056 26666 33108
rect 29638 33096 29644 33108
rect 27080 33068 29644 33096
rect 27080 33040 27108 33068
rect 29638 33056 29644 33068
rect 29696 33056 29702 33108
rect 29730 33056 29736 33108
rect 29788 33096 29794 33108
rect 30101 33099 30159 33105
rect 30101 33096 30113 33099
rect 29788 33068 30113 33096
rect 29788 33056 29794 33068
rect 30101 33065 30113 33068
rect 30147 33065 30159 33099
rect 30101 33059 30159 33065
rect 35161 33099 35219 33105
rect 35161 33065 35173 33099
rect 35207 33096 35219 33099
rect 35434 33096 35440 33108
rect 35207 33068 35440 33096
rect 35207 33065 35219 33068
rect 35161 33059 35219 33065
rect 35434 33056 35440 33068
rect 35492 33096 35498 33108
rect 36449 33099 36507 33105
rect 36449 33096 36461 33099
rect 35492 33068 36461 33096
rect 35492 33056 35498 33068
rect 36449 33065 36461 33068
rect 36495 33065 36507 33099
rect 36449 33059 36507 33065
rect 36538 33056 36544 33108
rect 36596 33096 36602 33108
rect 36817 33099 36875 33105
rect 36817 33096 36829 33099
rect 36596 33068 36829 33096
rect 36596 33056 36602 33068
rect 36817 33065 36829 33068
rect 36863 33065 36875 33099
rect 36817 33059 36875 33065
rect 38102 33056 38108 33108
rect 38160 33096 38166 33108
rect 38930 33096 38936 33108
rect 38160 33068 38936 33096
rect 38160 33056 38166 33068
rect 38930 33056 38936 33068
rect 38988 33056 38994 33108
rect 23164 33000 23474 33028
rect 23164 32988 23170 33000
rect 25130 32988 25136 33040
rect 25188 33028 25194 33040
rect 26697 33031 26755 33037
rect 26697 33028 26709 33031
rect 25188 33000 26709 33028
rect 25188 32988 25194 33000
rect 26697 32997 26709 33000
rect 26743 33028 26755 33031
rect 27062 33028 27068 33040
rect 26743 33000 27068 33028
rect 26743 32997 26755 33000
rect 26697 32991 26755 32997
rect 27062 32988 27068 33000
rect 27120 32988 27126 33040
rect 28626 33028 28632 33040
rect 28587 33000 28632 33028
rect 28626 32988 28632 33000
rect 28684 32988 28690 33040
rect 32125 33031 32183 33037
rect 32125 32997 32137 33031
rect 32171 33028 32183 33031
rect 32950 33028 32956 33040
rect 32171 33000 32956 33028
rect 32171 32997 32183 33000
rect 32125 32991 32183 32997
rect 32950 32988 32956 33000
rect 33008 32988 33014 33040
rect 41046 33028 41052 33040
rect 41007 33000 41052 33028
rect 41046 32988 41052 33000
rect 41104 32988 41110 33040
rect 44818 33028 44824 33040
rect 44779 33000 44824 33028
rect 44818 32988 44824 33000
rect 44876 32988 44882 33040
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 13964 32932 14105 32960
rect 13964 32920 13970 32932
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 14093 32923 14151 32929
rect 17037 32963 17095 32969
rect 17037 32929 17049 32963
rect 17083 32929 17095 32963
rect 17037 32923 17095 32929
rect 17126 32920 17132 32972
rect 17184 32960 17190 32972
rect 17313 32963 17371 32969
rect 17313 32960 17325 32963
rect 17184 32932 17325 32960
rect 17184 32920 17190 32932
rect 17313 32929 17325 32932
rect 17359 32929 17371 32963
rect 17313 32923 17371 32929
rect 18138 32920 18144 32972
rect 18196 32960 18202 32972
rect 18196 32932 19840 32960
rect 18196 32920 18202 32932
rect 14366 32892 14372 32904
rect 14327 32864 14372 32892
rect 14366 32852 14372 32864
rect 14424 32852 14430 32904
rect 15838 32892 15844 32904
rect 15799 32864 15844 32892
rect 15838 32852 15844 32864
rect 15896 32852 15902 32904
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32892 17647 32895
rect 18046 32892 18052 32904
rect 17635 32864 18052 32892
rect 17635 32861 17647 32864
rect 17589 32855 17647 32861
rect 18046 32852 18052 32864
rect 18104 32892 18110 32904
rect 18693 32895 18751 32901
rect 18693 32892 18705 32895
rect 18104 32864 18705 32892
rect 18104 32852 18110 32864
rect 18693 32861 18705 32864
rect 18739 32861 18751 32895
rect 19058 32892 19064 32904
rect 19019 32864 19064 32892
rect 18693 32855 18751 32861
rect 19058 32852 19064 32864
rect 19116 32852 19122 32904
rect 19812 32892 19840 32932
rect 19886 32920 19892 32972
rect 19944 32960 19950 32972
rect 19981 32963 20039 32969
rect 19981 32960 19993 32963
rect 19944 32932 19993 32960
rect 19944 32920 19950 32932
rect 19981 32929 19993 32932
rect 20027 32960 20039 32963
rect 20070 32960 20076 32972
rect 20027 32932 20076 32960
rect 20027 32929 20039 32932
rect 19981 32923 20039 32929
rect 20070 32920 20076 32932
rect 20128 32920 20134 32972
rect 23201 32963 23259 32969
rect 23201 32929 23213 32963
rect 23247 32960 23259 32963
rect 23290 32960 23296 32972
rect 23247 32932 23296 32960
rect 23247 32929 23259 32932
rect 23201 32923 23259 32929
rect 23290 32920 23296 32932
rect 23348 32920 23354 32972
rect 25314 32920 25320 32972
rect 25372 32960 25378 32972
rect 25444 32963 25502 32969
rect 25444 32960 25456 32963
rect 25372 32932 25456 32960
rect 25372 32920 25378 32932
rect 25444 32929 25456 32932
rect 25490 32929 25502 32963
rect 30282 32960 30288 32972
rect 30243 32932 30288 32960
rect 25444 32923 25502 32929
rect 30282 32920 30288 32932
rect 30340 32920 30346 32972
rect 30558 32960 30564 32972
rect 30519 32932 30564 32960
rect 30558 32920 30564 32932
rect 30616 32920 30622 32972
rect 32306 32920 32312 32972
rect 32364 32920 32370 32972
rect 33873 32963 33931 32969
rect 33873 32929 33885 32963
rect 33919 32929 33931 32963
rect 34238 32960 34244 32972
rect 34199 32932 34244 32960
rect 33873 32923 33931 32929
rect 20993 32895 21051 32901
rect 20993 32892 21005 32895
rect 19812 32864 21005 32892
rect 20993 32861 21005 32864
rect 21039 32892 21051 32895
rect 22646 32892 22652 32904
rect 21039 32864 22652 32892
rect 21039 32861 21051 32864
rect 20993 32855 21051 32861
rect 22646 32852 22652 32864
rect 22704 32852 22710 32904
rect 26605 32895 26663 32901
rect 26605 32892 26617 32895
rect 26160 32864 26617 32892
rect 21545 32827 21603 32833
rect 21545 32793 21557 32827
rect 21591 32824 21603 32827
rect 21634 32824 21640 32836
rect 21591 32796 21640 32824
rect 21591 32793 21603 32796
rect 21545 32787 21603 32793
rect 21634 32784 21640 32796
rect 21692 32784 21698 32836
rect 26160 32768 26188 32864
rect 26605 32861 26617 32864
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 27249 32895 27307 32901
rect 27249 32861 27261 32895
rect 27295 32892 27307 32895
rect 27430 32892 27436 32904
rect 27295 32864 27436 32892
rect 27295 32861 27307 32864
rect 27249 32855 27307 32861
rect 27430 32852 27436 32864
rect 27488 32892 27494 32904
rect 27706 32892 27712 32904
rect 27488 32864 27712 32892
rect 27488 32852 27494 32864
rect 27706 32852 27712 32864
rect 27764 32852 27770 32904
rect 28534 32892 28540 32904
rect 28495 32864 28540 32892
rect 28534 32852 28540 32864
rect 28592 32852 28598 32904
rect 32324 32892 32352 32920
rect 32490 32892 32496 32904
rect 32324 32864 32496 32892
rect 32490 32852 32496 32864
rect 32548 32852 32554 32904
rect 32582 32852 32588 32904
rect 32640 32892 32646 32904
rect 32640 32864 32685 32892
rect 32640 32852 32646 32864
rect 29086 32824 29092 32836
rect 29047 32796 29092 32824
rect 29086 32784 29092 32796
rect 29144 32784 29150 32836
rect 31110 32784 31116 32836
rect 31168 32824 31174 32836
rect 31205 32827 31263 32833
rect 31205 32824 31217 32827
rect 31168 32796 31217 32824
rect 31168 32784 31174 32796
rect 31205 32793 31217 32796
rect 31251 32824 31263 32827
rect 31573 32827 31631 32833
rect 31573 32824 31585 32827
rect 31251 32796 31585 32824
rect 31251 32793 31263 32796
rect 31205 32787 31263 32793
rect 31573 32793 31585 32796
rect 31619 32824 31631 32827
rect 31846 32824 31852 32836
rect 31619 32796 31852 32824
rect 31619 32793 31631 32796
rect 31573 32787 31631 32793
rect 31846 32784 31852 32796
rect 31904 32824 31910 32836
rect 32263 32827 32321 32833
rect 32263 32824 32275 32827
rect 31904 32796 32275 32824
rect 31904 32784 31910 32796
rect 32263 32793 32275 32796
rect 32309 32793 32321 32827
rect 32263 32787 32321 32793
rect 33686 32784 33692 32836
rect 33744 32824 33750 32836
rect 33888 32824 33916 32923
rect 34238 32920 34244 32932
rect 34296 32960 34302 32972
rect 34977 32963 35035 32969
rect 34977 32960 34989 32963
rect 34296 32932 34989 32960
rect 34296 32920 34302 32932
rect 34977 32929 34989 32932
rect 35023 32929 35035 32963
rect 35250 32960 35256 32972
rect 35163 32932 35256 32960
rect 34977 32923 35035 32929
rect 34992 32892 35020 32923
rect 35250 32920 35256 32932
rect 35308 32960 35314 32972
rect 35434 32960 35440 32972
rect 35308 32932 35440 32960
rect 35308 32920 35314 32932
rect 35434 32920 35440 32932
rect 35492 32920 35498 32972
rect 36078 32920 36084 32972
rect 36136 32960 36142 32972
rect 37458 32960 37464 32972
rect 36136 32932 37464 32960
rect 36136 32920 36142 32932
rect 37458 32920 37464 32932
rect 37516 32960 37522 32972
rect 37737 32963 37795 32969
rect 37737 32960 37749 32963
rect 37516 32932 37749 32960
rect 37516 32920 37522 32932
rect 37737 32929 37749 32932
rect 37783 32929 37795 32963
rect 38194 32960 38200 32972
rect 38155 32932 38200 32960
rect 37737 32923 37795 32929
rect 38194 32920 38200 32932
rect 38252 32920 38258 32972
rect 39758 32920 39764 32972
rect 39816 32960 39822 32972
rect 39888 32963 39946 32969
rect 39888 32960 39900 32963
rect 39816 32932 39900 32960
rect 39816 32920 39822 32932
rect 39888 32929 39900 32932
rect 39934 32929 39946 32963
rect 39888 32923 39946 32929
rect 43692 32963 43750 32969
rect 43692 32929 43704 32963
rect 43738 32960 43750 32963
rect 43806 32960 43812 32972
rect 43738 32932 43812 32960
rect 43738 32929 43750 32932
rect 43692 32923 43750 32929
rect 43806 32920 43812 32932
rect 43864 32920 43870 32972
rect 45738 32920 45744 32972
rect 45796 32960 45802 32972
rect 46236 32963 46294 32969
rect 46236 32960 46248 32963
rect 45796 32932 46248 32960
rect 45796 32920 45802 32932
rect 46236 32929 46248 32932
rect 46282 32929 46294 32963
rect 46236 32923 46294 32929
rect 35621 32895 35679 32901
rect 35621 32892 35633 32895
rect 34992 32864 35633 32892
rect 35621 32861 35633 32864
rect 35667 32892 35679 32895
rect 35710 32892 35716 32904
rect 35667 32864 35716 32892
rect 35667 32861 35679 32864
rect 35621 32855 35679 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 38102 32852 38108 32904
rect 38160 32892 38166 32904
rect 38289 32895 38347 32901
rect 38289 32892 38301 32895
rect 38160 32864 38301 32892
rect 38160 32852 38166 32864
rect 38289 32861 38301 32864
rect 38335 32861 38347 32895
rect 38289 32855 38347 32861
rect 39991 32895 40049 32901
rect 39991 32861 40003 32895
rect 40037 32892 40049 32895
rect 40310 32892 40316 32904
rect 40037 32864 40316 32892
rect 40037 32861 40049 32864
rect 39991 32855 40049 32861
rect 40310 32852 40316 32864
rect 40368 32892 40374 32904
rect 40957 32895 41015 32901
rect 40957 32892 40969 32895
rect 40368 32864 40969 32892
rect 40368 32852 40374 32864
rect 40957 32861 40969 32864
rect 41003 32861 41015 32895
rect 40957 32855 41015 32861
rect 41601 32895 41659 32901
rect 41601 32861 41613 32895
rect 41647 32892 41659 32895
rect 41874 32892 41880 32904
rect 41647 32864 41880 32892
rect 41647 32861 41659 32864
rect 41601 32855 41659 32861
rect 41874 32852 41880 32864
rect 41932 32852 41938 32904
rect 44726 32892 44732 32904
rect 44687 32864 44732 32892
rect 44726 32852 44732 32864
rect 44784 32852 44790 32904
rect 45002 32892 45008 32904
rect 44963 32864 45008 32892
rect 45002 32852 45008 32864
rect 45060 32852 45066 32904
rect 33744 32796 33916 32824
rect 33744 32784 33750 32796
rect 18417 32759 18475 32765
rect 18417 32725 18429 32759
rect 18463 32756 18475 32759
rect 18598 32756 18604 32768
rect 18463 32728 18604 32756
rect 18463 32725 18475 32728
rect 18417 32719 18475 32725
rect 18598 32716 18604 32728
rect 18656 32756 18662 32768
rect 19242 32756 19248 32768
rect 18656 32728 19248 32756
rect 18656 32716 18662 32728
rect 19242 32716 19248 32728
rect 19300 32716 19306 32768
rect 20254 32756 20260 32768
rect 20215 32728 20260 32756
rect 20254 32716 20260 32728
rect 20312 32716 20318 32768
rect 20622 32716 20628 32768
rect 20680 32756 20686 32768
rect 25406 32756 25412 32768
rect 20680 32728 25412 32756
rect 20680 32716 20686 32728
rect 25406 32716 25412 32728
rect 25464 32716 25470 32768
rect 25547 32759 25605 32765
rect 25547 32725 25559 32759
rect 25593 32756 25605 32759
rect 26142 32756 26148 32768
rect 25593 32728 26148 32756
rect 25593 32725 25605 32728
rect 25547 32719 25605 32725
rect 26142 32716 26148 32728
rect 26200 32716 26206 32768
rect 27522 32756 27528 32768
rect 27483 32728 27528 32756
rect 27522 32716 27528 32728
rect 27580 32716 27586 32768
rect 31938 32756 31944 32768
rect 31899 32728 31944 32756
rect 31938 32716 31944 32728
rect 31996 32716 32002 32768
rect 32398 32756 32404 32768
rect 32359 32728 32404 32756
rect 32398 32716 32404 32728
rect 32456 32716 32462 32768
rect 33505 32759 33563 32765
rect 33505 32725 33517 32759
rect 33551 32756 33563 32759
rect 33594 32756 33600 32768
rect 33551 32728 33600 32756
rect 33551 32725 33563 32728
rect 33505 32719 33563 32725
rect 33594 32716 33600 32728
rect 33652 32716 33658 32768
rect 33778 32756 33784 32768
rect 33739 32728 33784 32756
rect 33778 32716 33784 32728
rect 33836 32716 33842 32768
rect 33888 32756 33916 32796
rect 33962 32784 33968 32836
rect 34020 32824 34026 32836
rect 35391 32827 35449 32833
rect 35391 32824 35403 32827
rect 34020 32796 35403 32824
rect 34020 32784 34026 32796
rect 35391 32793 35403 32796
rect 35437 32824 35449 32827
rect 35802 32824 35808 32836
rect 35437 32796 35808 32824
rect 35437 32793 35449 32796
rect 35391 32787 35449 32793
rect 35802 32784 35808 32796
rect 35860 32824 35866 32836
rect 36354 32824 36360 32836
rect 35860 32796 36360 32824
rect 35860 32784 35866 32796
rect 36354 32784 36360 32796
rect 36412 32824 36418 32836
rect 37185 32827 37243 32833
rect 37185 32824 37197 32827
rect 36412 32796 37197 32824
rect 36412 32784 36418 32796
rect 37185 32793 37197 32796
rect 37231 32793 37243 32827
rect 37185 32787 37243 32793
rect 34698 32756 34704 32768
rect 33888 32728 34704 32756
rect 34698 32716 34704 32728
rect 34756 32756 34762 32768
rect 35161 32759 35219 32765
rect 35161 32756 35173 32759
rect 34756 32728 35173 32756
rect 34756 32716 34762 32728
rect 35161 32725 35173 32728
rect 35207 32756 35219 32759
rect 35529 32759 35587 32765
rect 35529 32756 35541 32759
rect 35207 32728 35541 32756
rect 35207 32725 35219 32728
rect 35161 32719 35219 32725
rect 35529 32725 35541 32728
rect 35575 32725 35587 32759
rect 35894 32756 35900 32768
rect 35855 32728 35900 32756
rect 35529 32719 35587 32725
rect 35894 32716 35900 32728
rect 35952 32716 35958 32768
rect 38010 32716 38016 32768
rect 38068 32756 38074 32768
rect 38749 32759 38807 32765
rect 38749 32756 38761 32759
rect 38068 32728 38761 32756
rect 38068 32716 38074 32728
rect 38749 32725 38761 32728
rect 38795 32725 38807 32759
rect 38749 32719 38807 32725
rect 43763 32759 43821 32765
rect 43763 32725 43775 32759
rect 43809 32756 43821 32759
rect 44361 32759 44419 32765
rect 44361 32756 44373 32759
rect 43809 32728 44373 32756
rect 43809 32725 43821 32728
rect 43763 32719 43821 32725
rect 44361 32725 44373 32728
rect 44407 32756 44419 32759
rect 44450 32756 44456 32768
rect 44407 32728 44456 32756
rect 44407 32725 44419 32728
rect 44361 32719 44419 32725
rect 44450 32716 44456 32728
rect 44508 32716 44514 32768
rect 45830 32716 45836 32768
rect 45888 32756 45894 32768
rect 46339 32759 46397 32765
rect 46339 32756 46351 32759
rect 45888 32728 46351 32756
rect 45888 32716 45894 32728
rect 46339 32725 46351 32728
rect 46385 32725 46397 32759
rect 46339 32719 46397 32725
rect 1104 32666 48852 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 48852 32666
rect 1104 32592 48852 32614
rect 13495 32555 13553 32561
rect 13495 32521 13507 32555
rect 13541 32552 13553 32555
rect 13814 32552 13820 32564
rect 13541 32524 13820 32552
rect 13541 32521 13553 32524
rect 13495 32515 13553 32521
rect 13814 32512 13820 32524
rect 13872 32512 13878 32564
rect 13909 32555 13967 32561
rect 13909 32521 13921 32555
rect 13955 32552 13967 32555
rect 13998 32552 14004 32564
rect 13955 32524 14004 32552
rect 13955 32521 13967 32524
rect 13909 32515 13967 32521
rect 12897 32419 12955 32425
rect 12897 32385 12909 32419
rect 12943 32416 12955 32419
rect 13814 32416 13820 32428
rect 12943 32388 13820 32416
rect 12943 32385 12955 32388
rect 12897 32379 12955 32385
rect 13814 32376 13820 32388
rect 13872 32376 13878 32428
rect 13424 32351 13482 32357
rect 13424 32317 13436 32351
rect 13470 32348 13482 32351
rect 13538 32348 13544 32360
rect 13470 32320 13544 32348
rect 13470 32317 13482 32320
rect 13424 32311 13482 32317
rect 13538 32308 13544 32320
rect 13596 32348 13602 32360
rect 13924 32348 13952 32515
rect 13998 32512 14004 32524
rect 14056 32512 14062 32564
rect 14277 32555 14335 32561
rect 14277 32521 14289 32555
rect 14323 32552 14335 32555
rect 14550 32552 14556 32564
rect 14323 32524 14556 32552
rect 14323 32521 14335 32524
rect 14277 32515 14335 32521
rect 14550 32512 14556 32524
rect 14608 32512 14614 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 15933 32555 15991 32561
rect 15933 32552 15945 32555
rect 15436 32524 15945 32552
rect 15436 32512 15442 32524
rect 15933 32521 15945 32524
rect 15979 32521 15991 32555
rect 16850 32552 16856 32564
rect 16811 32524 16856 32552
rect 15933 32515 15991 32521
rect 16850 32512 16856 32524
rect 16908 32512 16914 32564
rect 17218 32512 17224 32564
rect 17276 32552 17282 32564
rect 17405 32555 17463 32561
rect 17405 32552 17417 32555
rect 17276 32524 17417 32552
rect 17276 32512 17282 32524
rect 17405 32521 17417 32524
rect 17451 32521 17463 32555
rect 17405 32515 17463 32521
rect 19058 32512 19064 32564
rect 19116 32552 19122 32564
rect 19613 32555 19671 32561
rect 19613 32552 19625 32555
rect 19116 32524 19625 32552
rect 19116 32512 19122 32524
rect 19613 32521 19625 32524
rect 19659 32521 19671 32555
rect 22646 32552 22652 32564
rect 22607 32524 22652 32552
rect 19613 32515 19671 32521
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 23290 32512 23296 32564
rect 23348 32552 23354 32564
rect 23845 32555 23903 32561
rect 23845 32552 23857 32555
rect 23348 32524 23857 32552
rect 23348 32512 23354 32524
rect 23845 32521 23857 32524
rect 23891 32521 23903 32555
rect 23845 32515 23903 32521
rect 24305 32555 24363 32561
rect 24305 32521 24317 32555
rect 24351 32552 24363 32555
rect 24578 32552 24584 32564
rect 24351 32524 24584 32552
rect 24351 32521 24363 32524
rect 24305 32515 24363 32521
rect 24578 32512 24584 32524
rect 24636 32512 24642 32564
rect 26142 32552 26148 32564
rect 26103 32524 26148 32552
rect 26142 32512 26148 32524
rect 26200 32512 26206 32564
rect 26467 32555 26525 32561
rect 26467 32521 26479 32555
rect 26513 32552 26525 32555
rect 26786 32552 26792 32564
rect 26513 32524 26792 32552
rect 26513 32521 26525 32524
rect 26467 32515 26525 32521
rect 26786 32512 26792 32524
rect 26844 32512 26850 32564
rect 27062 32512 27068 32564
rect 27120 32552 27126 32564
rect 27157 32555 27215 32561
rect 27157 32552 27169 32555
rect 27120 32524 27169 32552
rect 27120 32512 27126 32524
rect 27157 32521 27169 32524
rect 27203 32521 27215 32555
rect 27157 32515 27215 32521
rect 31757 32555 31815 32561
rect 31757 32521 31769 32555
rect 31803 32552 31815 32555
rect 32493 32555 32551 32561
rect 31803 32524 32306 32552
rect 31803 32521 31815 32524
rect 31757 32515 31815 32521
rect 15289 32487 15347 32493
rect 15289 32453 15301 32487
rect 15335 32484 15347 32487
rect 15562 32484 15568 32496
rect 15335 32456 15568 32484
rect 15335 32453 15347 32456
rect 15289 32447 15347 32453
rect 15562 32444 15568 32456
rect 15620 32444 15626 32496
rect 16390 32444 16396 32496
rect 16448 32484 16454 32496
rect 17773 32487 17831 32493
rect 17773 32484 17785 32487
rect 16448 32456 17785 32484
rect 16448 32444 16454 32456
rect 17773 32453 17785 32456
rect 17819 32453 17831 32487
rect 17773 32447 17831 32453
rect 14366 32416 14372 32428
rect 14327 32388 14372 32416
rect 14366 32376 14372 32388
rect 14424 32376 14430 32428
rect 13596 32320 13952 32348
rect 13596 32308 13602 32320
rect 16850 32308 16856 32360
rect 16908 32348 16914 32360
rect 16945 32351 17003 32357
rect 16945 32348 16957 32351
rect 16908 32320 16957 32348
rect 16908 32308 16914 32320
rect 16945 32317 16957 32320
rect 16991 32317 17003 32351
rect 16945 32311 17003 32317
rect 14550 32240 14556 32292
rect 14608 32280 14614 32292
rect 14690 32283 14748 32289
rect 14690 32280 14702 32283
rect 14608 32252 14702 32280
rect 14608 32240 14614 32252
rect 14690 32249 14702 32252
rect 14736 32249 14748 32283
rect 17788 32280 17816 32447
rect 20530 32444 20536 32496
rect 20588 32484 20594 32496
rect 20714 32484 20720 32496
rect 20588 32456 20720 32484
rect 20588 32444 20594 32456
rect 20714 32444 20720 32456
rect 20772 32484 20778 32496
rect 25314 32484 25320 32496
rect 20772 32456 25320 32484
rect 20772 32444 20778 32456
rect 25314 32444 25320 32456
rect 25372 32484 25378 32496
rect 25409 32487 25467 32493
rect 25409 32484 25421 32487
rect 25372 32456 25421 32484
rect 25372 32444 25378 32456
rect 25409 32453 25421 32456
rect 25455 32453 25467 32487
rect 25409 32447 25467 32453
rect 28626 32444 28632 32496
rect 28684 32484 28690 32496
rect 30193 32487 30251 32493
rect 30193 32484 30205 32487
rect 28684 32456 30205 32484
rect 28684 32444 28690 32456
rect 30193 32453 30205 32456
rect 30239 32453 30251 32487
rect 30193 32447 30251 32453
rect 18046 32416 18052 32428
rect 18007 32388 18052 32416
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 24486 32416 24492 32428
rect 24447 32388 24492 32416
rect 24486 32376 24492 32388
rect 24544 32376 24550 32428
rect 24762 32416 24768 32428
rect 24723 32388 24768 32416
rect 24762 32376 24768 32388
rect 24820 32376 24826 32428
rect 20140 32351 20198 32357
rect 20140 32317 20152 32351
rect 20186 32348 20198 32351
rect 20346 32348 20352 32360
rect 20186 32320 20352 32348
rect 20186 32317 20198 32320
rect 20140 32311 20198 32317
rect 20346 32308 20352 32320
rect 20404 32348 20410 32360
rect 20530 32348 20536 32360
rect 20404 32320 20536 32348
rect 20404 32308 20410 32320
rect 20530 32308 20536 32320
rect 20588 32308 20594 32360
rect 21085 32351 21143 32357
rect 21085 32317 21097 32351
rect 21131 32348 21143 32351
rect 21726 32348 21732 32360
rect 21131 32320 21732 32348
rect 21131 32317 21143 32320
rect 21085 32311 21143 32317
rect 21726 32308 21732 32320
rect 21784 32348 21790 32360
rect 21910 32348 21916 32360
rect 21784 32320 21916 32348
rect 21784 32308 21790 32320
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 25406 32308 25412 32360
rect 25464 32348 25470 32360
rect 26396 32351 26454 32357
rect 26396 32348 26408 32351
rect 25464 32320 26408 32348
rect 25464 32308 25470 32320
rect 26396 32317 26408 32320
rect 26442 32348 26454 32351
rect 29270 32348 29276 32360
rect 26442 32320 26924 32348
rect 29231 32320 29276 32348
rect 26442 32317 26454 32320
rect 26396 32311 26454 32317
rect 18370 32283 18428 32289
rect 18370 32280 18382 32283
rect 17788 32252 18382 32280
rect 14690 32243 14748 32249
rect 18370 32249 18382 32252
rect 18416 32280 18428 32283
rect 19245 32283 19303 32289
rect 19245 32280 19257 32283
rect 18416 32252 19257 32280
rect 18416 32249 18428 32252
rect 18370 32243 18428 32249
rect 19245 32249 19257 32252
rect 19291 32280 19303 32283
rect 19334 32280 19340 32292
rect 19291 32252 19340 32280
rect 19291 32249 19303 32252
rect 19245 32243 19303 32249
rect 19334 32240 19340 32252
rect 19392 32280 19398 32292
rect 20901 32283 20959 32289
rect 20901 32280 20913 32283
rect 19392 32252 20913 32280
rect 19392 32240 19398 32252
rect 20901 32249 20913 32252
rect 20947 32280 20959 32283
rect 21406 32283 21464 32289
rect 21406 32280 21418 32283
rect 20947 32252 21418 32280
rect 20947 32249 20959 32252
rect 20901 32243 20959 32249
rect 21406 32249 21418 32252
rect 21452 32280 21464 32283
rect 23106 32280 23112 32292
rect 21452 32252 23112 32280
rect 21452 32249 21464 32252
rect 21406 32243 21464 32249
rect 23106 32240 23112 32252
rect 23164 32280 23170 32292
rect 23201 32283 23259 32289
rect 23201 32280 23213 32283
rect 23164 32252 23213 32280
rect 23164 32240 23170 32252
rect 23201 32249 23213 32252
rect 23247 32249 23259 32283
rect 23201 32243 23259 32249
rect 24578 32240 24584 32292
rect 24636 32280 24642 32292
rect 24636 32252 24681 32280
rect 24636 32240 24642 32252
rect 13265 32215 13323 32221
rect 13265 32181 13277 32215
rect 13311 32212 13323 32215
rect 13630 32212 13636 32224
rect 13311 32184 13636 32212
rect 13311 32181 13323 32184
rect 13265 32175 13323 32181
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 16390 32212 16396 32224
rect 16351 32184 16396 32212
rect 16390 32172 16396 32184
rect 16448 32212 16454 32224
rect 17126 32212 17132 32224
rect 16448 32184 17132 32212
rect 16448 32172 16454 32184
rect 17126 32172 17132 32184
rect 17184 32172 17190 32224
rect 18966 32212 18972 32224
rect 18927 32184 18972 32212
rect 18966 32172 18972 32184
rect 19024 32172 19030 32224
rect 20211 32215 20269 32221
rect 20211 32181 20223 32215
rect 20257 32212 20269 32215
rect 20438 32212 20444 32224
rect 20257 32184 20444 32212
rect 20257 32181 20269 32184
rect 20211 32175 20269 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 21082 32172 21088 32224
rect 21140 32212 21146 32224
rect 26896 32221 26924 32320
rect 29270 32308 29276 32320
rect 29328 32308 29334 32360
rect 31662 32308 31668 32360
rect 31720 32348 31726 32360
rect 31772 32348 31800 32515
rect 31846 32444 31852 32496
rect 31904 32484 31910 32496
rect 31987 32487 32045 32493
rect 31987 32484 31999 32487
rect 31904 32456 31999 32484
rect 31904 32444 31910 32456
rect 31987 32453 31999 32456
rect 32033 32453 32045 32487
rect 32122 32484 32128 32496
rect 32083 32456 32128 32484
rect 31987 32447 32045 32453
rect 32122 32444 32128 32456
rect 32180 32444 32186 32496
rect 32278 32484 32306 32524
rect 32493 32521 32505 32555
rect 32539 32552 32551 32555
rect 33134 32552 33140 32564
rect 32539 32524 33140 32552
rect 32539 32521 32551 32524
rect 32493 32515 32551 32521
rect 33134 32512 33140 32524
rect 33192 32512 33198 32564
rect 33321 32555 33379 32561
rect 33321 32521 33333 32555
rect 33367 32552 33379 32555
rect 34238 32552 34244 32564
rect 33367 32524 34244 32552
rect 33367 32521 33379 32524
rect 33321 32515 33379 32521
rect 34238 32512 34244 32524
rect 34296 32512 34302 32564
rect 34698 32552 34704 32564
rect 34659 32524 34704 32552
rect 34698 32512 34704 32524
rect 34756 32512 34762 32564
rect 35161 32555 35219 32561
rect 35161 32521 35173 32555
rect 35207 32552 35219 32555
rect 35434 32552 35440 32564
rect 35207 32524 35440 32552
rect 35207 32521 35219 32524
rect 35161 32515 35219 32521
rect 35434 32512 35440 32524
rect 35492 32512 35498 32564
rect 35529 32555 35587 32561
rect 35529 32521 35541 32555
rect 35575 32552 35587 32555
rect 36262 32552 36268 32564
rect 35575 32524 36268 32552
rect 35575 32521 35587 32524
rect 35529 32515 35587 32521
rect 36262 32512 36268 32524
rect 36320 32512 36326 32564
rect 37458 32552 37464 32564
rect 37419 32524 37464 32552
rect 37458 32512 37464 32524
rect 37516 32512 37522 32564
rect 38194 32512 38200 32564
rect 38252 32552 38258 32564
rect 39209 32555 39267 32561
rect 39209 32552 39221 32555
rect 38252 32524 39221 32552
rect 38252 32512 38258 32524
rect 39209 32521 39221 32524
rect 39255 32521 39267 32555
rect 40310 32552 40316 32564
rect 40271 32524 40316 32552
rect 39209 32515 39267 32521
rect 40310 32512 40316 32524
rect 40368 32512 40374 32564
rect 40957 32555 41015 32561
rect 40957 32521 40969 32555
rect 41003 32552 41015 32555
rect 41046 32552 41052 32564
rect 41003 32524 41052 32552
rect 41003 32521 41015 32524
rect 40957 32515 41015 32521
rect 41046 32512 41052 32524
rect 41104 32512 41110 32564
rect 41877 32555 41935 32561
rect 41877 32521 41889 32555
rect 41923 32552 41935 32555
rect 43625 32555 43683 32561
rect 43625 32552 43637 32555
rect 41923 32524 43637 32552
rect 41923 32521 41935 32524
rect 41877 32515 41935 32521
rect 43625 32521 43637 32524
rect 43671 32552 43683 32555
rect 43671 32524 45140 32552
rect 43671 32521 43683 32524
rect 43625 32515 43683 32521
rect 32950 32484 32956 32496
rect 32278 32456 32956 32484
rect 32950 32444 32956 32456
rect 33008 32444 33014 32496
rect 34333 32487 34391 32493
rect 34333 32453 34345 32487
rect 34379 32484 34391 32487
rect 34606 32484 34612 32496
rect 34379 32456 34612 32484
rect 34379 32453 34391 32456
rect 34333 32447 34391 32453
rect 32217 32419 32275 32425
rect 32217 32385 32229 32419
rect 32263 32385 32275 32419
rect 33870 32416 33876 32428
rect 33831 32388 33876 32416
rect 32217 32379 32275 32385
rect 31849 32351 31907 32357
rect 31849 32348 31861 32351
rect 31720 32320 31861 32348
rect 31720 32308 31726 32320
rect 31849 32317 31861 32320
rect 31895 32317 31907 32351
rect 31849 32311 31907 32317
rect 31938 32308 31944 32360
rect 31996 32348 32002 32360
rect 32232 32348 32260 32379
rect 33870 32376 33876 32388
rect 33928 32376 33934 32428
rect 33594 32348 33600 32360
rect 31996 32320 32260 32348
rect 33555 32320 33600 32348
rect 31996 32308 32002 32320
rect 33594 32308 33600 32320
rect 33652 32308 33658 32360
rect 34348 32348 34376 32447
rect 34606 32444 34612 32456
rect 34664 32444 34670 32496
rect 35710 32444 35716 32496
rect 35768 32484 35774 32496
rect 35897 32487 35955 32493
rect 35897 32484 35909 32487
rect 35768 32456 35909 32484
rect 35768 32444 35774 32456
rect 35897 32453 35909 32456
rect 35943 32453 35955 32487
rect 35897 32447 35955 32453
rect 38933 32487 38991 32493
rect 38933 32453 38945 32487
rect 38979 32484 38991 32487
rect 44177 32487 44235 32493
rect 44177 32484 44189 32487
rect 38979 32456 44189 32484
rect 38979 32453 38991 32456
rect 38933 32447 38991 32453
rect 44177 32453 44189 32456
rect 44223 32453 44235 32487
rect 44177 32447 44235 32453
rect 35253 32419 35311 32425
rect 35253 32385 35265 32419
rect 35299 32416 35311 32419
rect 35342 32416 35348 32428
rect 35299 32388 35348 32416
rect 35299 32385 35311 32388
rect 35253 32379 35311 32385
rect 35342 32376 35348 32388
rect 35400 32376 35406 32428
rect 36538 32416 36544 32428
rect 36096 32388 36544 32416
rect 34072 32320 34376 32348
rect 27430 32280 27436 32292
rect 27391 32252 27436 32280
rect 27430 32240 27436 32252
rect 27488 32240 27494 32292
rect 27522 32240 27528 32292
rect 27580 32280 27586 32292
rect 27580 32252 27625 32280
rect 27580 32240 27586 32252
rect 27706 32240 27712 32292
rect 27764 32280 27770 32292
rect 28077 32283 28135 32289
rect 28077 32280 28089 32283
rect 27764 32252 28089 32280
rect 27764 32240 27770 32252
rect 28077 32249 28089 32252
rect 28123 32280 28135 32283
rect 28442 32280 28448 32292
rect 28123 32252 28448 32280
rect 28123 32249 28135 32252
rect 28077 32243 28135 32249
rect 28442 32240 28448 32252
rect 28500 32240 28506 32292
rect 29089 32283 29147 32289
rect 29089 32280 29101 32283
rect 28966 32252 29101 32280
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21140 32184 22017 32212
rect 21140 32172 21146 32184
rect 22005 32181 22017 32184
rect 22051 32212 22063 32215
rect 22281 32215 22339 32221
rect 22281 32212 22293 32215
rect 22051 32184 22293 32212
rect 22051 32181 22063 32184
rect 22005 32175 22063 32181
rect 22281 32181 22293 32184
rect 22327 32181 22339 32215
rect 22281 32175 22339 32181
rect 26881 32215 26939 32221
rect 26881 32181 26893 32215
rect 26927 32212 26939 32215
rect 27062 32212 27068 32224
rect 26927 32184 27068 32212
rect 26927 32181 26939 32184
rect 26881 32175 26939 32181
rect 27062 32172 27068 32184
rect 27120 32172 27126 32224
rect 27540 32212 27568 32240
rect 28537 32215 28595 32221
rect 28537 32212 28549 32215
rect 27540 32184 28549 32212
rect 28537 32181 28549 32184
rect 28583 32212 28595 32215
rect 28626 32212 28632 32224
rect 28583 32184 28632 32212
rect 28583 32181 28595 32184
rect 28537 32175 28595 32181
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 28718 32172 28724 32224
rect 28776 32212 28782 32224
rect 28966 32212 28994 32252
rect 29089 32249 29101 32252
rect 29135 32280 29147 32283
rect 29635 32283 29693 32289
rect 29635 32280 29647 32283
rect 29135 32252 29647 32280
rect 29135 32249 29147 32252
rect 29089 32243 29147 32249
rect 29635 32249 29647 32252
rect 29681 32280 29693 32283
rect 29822 32280 29828 32292
rect 29681 32252 29828 32280
rect 29681 32249 29693 32252
rect 29635 32243 29693 32249
rect 29822 32240 29828 32252
rect 29880 32240 29886 32292
rect 33413 32283 33471 32289
rect 33413 32249 33425 32283
rect 33459 32280 33471 32283
rect 34072 32280 34100 32320
rect 34790 32308 34796 32360
rect 34848 32348 34854 32360
rect 35032 32351 35090 32357
rect 35032 32348 35044 32351
rect 34848 32320 35044 32348
rect 34848 32308 34854 32320
rect 35032 32317 35044 32320
rect 35078 32348 35090 32351
rect 35986 32348 35992 32360
rect 35078 32320 35992 32348
rect 35078 32317 35090 32320
rect 35032 32311 35090 32317
rect 35986 32308 35992 32320
rect 36044 32308 36050 32360
rect 33459 32252 34100 32280
rect 33459 32249 33471 32252
rect 33413 32243 33471 32249
rect 34882 32240 34888 32292
rect 34940 32280 34946 32292
rect 36096 32280 36124 32388
rect 36538 32376 36544 32388
rect 36596 32376 36602 32428
rect 37185 32419 37243 32425
rect 37185 32385 37197 32419
rect 37231 32416 37243 32419
rect 38010 32416 38016 32428
rect 37231 32388 38016 32416
rect 37231 32385 37243 32388
rect 37185 32379 37243 32385
rect 38010 32376 38016 32388
rect 38068 32376 38074 32428
rect 40954 32376 40960 32428
rect 41012 32416 41018 32428
rect 41141 32419 41199 32425
rect 41141 32416 41153 32419
rect 41012 32388 41153 32416
rect 41012 32376 41018 32388
rect 41141 32385 41153 32388
rect 41187 32416 41199 32419
rect 42061 32419 42119 32425
rect 42061 32416 42073 32419
rect 41187 32388 42073 32416
rect 41187 32385 41199 32388
rect 41141 32379 41199 32385
rect 42061 32385 42073 32388
rect 42107 32385 42119 32419
rect 42061 32379 42119 32385
rect 42150 32376 42156 32428
rect 42208 32416 42214 32428
rect 42886 32416 42892 32428
rect 42208 32388 42892 32416
rect 42208 32376 42214 32388
rect 42886 32376 42892 32388
rect 42944 32376 42950 32428
rect 43533 32419 43591 32425
rect 43533 32385 43545 32419
rect 43579 32416 43591 32419
rect 43625 32419 43683 32425
rect 43625 32416 43637 32419
rect 43579 32388 43637 32416
rect 43579 32385 43591 32388
rect 43533 32379 43591 32385
rect 43625 32385 43637 32388
rect 43671 32385 43683 32419
rect 43625 32379 43683 32385
rect 36449 32351 36507 32357
rect 36449 32317 36461 32351
rect 36495 32348 36507 32351
rect 36630 32348 36636 32360
rect 36495 32320 36636 32348
rect 36495 32317 36507 32320
rect 36449 32311 36507 32317
rect 36262 32280 36268 32292
rect 34940 32252 36124 32280
rect 36223 32252 36268 32280
rect 34940 32240 34946 32252
rect 36262 32240 36268 32252
rect 36320 32280 36326 32292
rect 36464 32280 36492 32311
rect 36630 32308 36636 32320
rect 36688 32308 36694 32360
rect 36906 32308 36912 32360
rect 36964 32348 36970 32360
rect 37001 32351 37059 32357
rect 37001 32348 37013 32351
rect 36964 32320 37013 32348
rect 36964 32308 36970 32320
rect 37001 32317 37013 32320
rect 37047 32348 37059 32351
rect 38194 32348 38200 32360
rect 37047 32320 38200 32348
rect 37047 32317 37059 32320
rect 37001 32311 37059 32317
rect 38194 32308 38200 32320
rect 38252 32308 38258 32360
rect 41782 32308 41788 32360
rect 41840 32348 41846 32360
rect 41877 32351 41935 32357
rect 41877 32348 41889 32351
rect 41840 32320 41889 32348
rect 41840 32308 41846 32320
rect 41877 32317 41889 32320
rect 41923 32317 41935 32351
rect 41877 32311 41935 32317
rect 36320 32252 36492 32280
rect 37829 32283 37887 32289
rect 36320 32240 36326 32252
rect 37829 32249 37841 32283
rect 37875 32280 37887 32283
rect 38375 32283 38433 32289
rect 38375 32280 38387 32283
rect 37875 32252 38387 32280
rect 37875 32249 37887 32252
rect 37829 32243 37887 32249
rect 38375 32249 38387 32252
rect 38421 32280 38433 32283
rect 38654 32280 38660 32292
rect 38421 32252 38660 32280
rect 38421 32249 38433 32252
rect 38375 32243 38433 32249
rect 38654 32240 38660 32252
rect 38712 32240 38718 32292
rect 41138 32240 41144 32292
rect 41196 32280 41202 32292
rect 41233 32283 41291 32289
rect 41233 32280 41245 32283
rect 41196 32252 41245 32280
rect 41196 32240 41202 32252
rect 41233 32249 41245 32252
rect 41279 32249 41291 32283
rect 42886 32280 42892 32292
rect 42847 32252 42892 32280
rect 41233 32243 41291 32249
rect 42886 32240 42892 32252
rect 42944 32240 42950 32292
rect 42981 32283 43039 32289
rect 42981 32249 42993 32283
rect 43027 32249 43039 32283
rect 44192 32280 44220 32447
rect 44450 32416 44456 32428
rect 44411 32388 44456 32416
rect 44450 32376 44456 32388
rect 44508 32376 44514 32428
rect 45112 32357 45140 32524
rect 46201 32419 46259 32425
rect 46201 32385 46213 32419
rect 46247 32416 46259 32419
rect 46658 32416 46664 32428
rect 46247 32388 46664 32416
rect 46247 32385 46259 32388
rect 46201 32379 46259 32385
rect 46658 32376 46664 32388
rect 46716 32416 46722 32428
rect 47121 32419 47179 32425
rect 47121 32416 47133 32419
rect 46716 32388 47133 32416
rect 46716 32376 46722 32388
rect 47121 32385 47133 32388
rect 47167 32385 47179 32419
rect 47121 32379 47179 32385
rect 45097 32351 45155 32357
rect 45097 32317 45109 32351
rect 45143 32348 45155 32351
rect 45554 32348 45560 32360
rect 45143 32320 45560 32348
rect 45143 32317 45155 32320
rect 45097 32311 45155 32317
rect 45554 32308 45560 32320
rect 45612 32308 45618 32360
rect 44545 32283 44603 32289
rect 44545 32280 44557 32283
rect 44192 32252 44557 32280
rect 42981 32243 43039 32249
rect 44545 32249 44557 32252
rect 44591 32280 44603 32283
rect 44818 32280 44824 32292
rect 44591 32252 44824 32280
rect 44591 32249 44603 32252
rect 44545 32243 44603 32249
rect 30650 32212 30656 32224
rect 28776 32184 28994 32212
rect 30611 32184 30656 32212
rect 28776 32172 28782 32184
rect 30650 32172 30656 32184
rect 30708 32172 30714 32224
rect 31021 32215 31079 32221
rect 31021 32181 31033 32215
rect 31067 32212 31079 32215
rect 31389 32215 31447 32221
rect 31389 32212 31401 32215
rect 31067 32184 31401 32212
rect 31067 32181 31079 32184
rect 31021 32175 31079 32181
rect 31389 32181 31401 32184
rect 31435 32212 31447 32215
rect 32398 32212 32404 32224
rect 31435 32184 32404 32212
rect 31435 32181 31447 32184
rect 31389 32175 31447 32181
rect 32398 32172 32404 32184
rect 32456 32212 32462 32224
rect 35434 32212 35440 32224
rect 32456 32184 35440 32212
rect 32456 32172 32462 32184
rect 35434 32172 35440 32184
rect 35492 32172 35498 32224
rect 37918 32172 37924 32224
rect 37976 32212 37982 32224
rect 39758 32212 39764 32224
rect 37976 32184 39764 32212
rect 37976 32172 37982 32184
rect 39758 32172 39764 32184
rect 39816 32212 39822 32224
rect 39853 32215 39911 32221
rect 39853 32212 39865 32215
rect 39816 32184 39865 32212
rect 39816 32172 39822 32184
rect 39853 32181 39865 32184
rect 39899 32181 39911 32215
rect 42610 32212 42616 32224
rect 42571 32184 42616 32212
rect 39853 32175 39911 32181
rect 42610 32172 42616 32184
rect 42668 32212 42674 32224
rect 42996 32212 43024 32243
rect 44818 32240 44824 32252
rect 44876 32240 44882 32292
rect 46293 32283 46351 32289
rect 46293 32280 46305 32283
rect 45388 32252 46305 32280
rect 43806 32212 43812 32224
rect 42668 32184 43024 32212
rect 43767 32184 43812 32212
rect 42668 32172 42674 32184
rect 43806 32172 43812 32184
rect 43864 32172 43870 32224
rect 44836 32212 44864 32240
rect 45186 32212 45192 32224
rect 44836 32184 45192 32212
rect 45186 32172 45192 32184
rect 45244 32212 45250 32224
rect 45388 32221 45416 32252
rect 46293 32249 46305 32252
rect 46339 32249 46351 32283
rect 46842 32280 46848 32292
rect 46803 32252 46848 32280
rect 46293 32243 46351 32249
rect 46842 32240 46848 32252
rect 46900 32240 46906 32292
rect 45373 32215 45431 32221
rect 45373 32212 45385 32215
rect 45244 32184 45385 32212
rect 45244 32172 45250 32184
rect 45373 32181 45385 32184
rect 45419 32181 45431 32215
rect 45373 32175 45431 32181
rect 45738 32172 45744 32224
rect 45796 32212 45802 32224
rect 45833 32215 45891 32221
rect 45833 32212 45845 32215
rect 45796 32184 45845 32212
rect 45796 32172 45802 32184
rect 45833 32181 45845 32184
rect 45879 32181 45891 32215
rect 45833 32175 45891 32181
rect 1104 32122 48852 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 48852 32122
rect 1104 32048 48852 32070
rect 14366 31968 14372 32020
rect 14424 32008 14430 32020
rect 14645 32011 14703 32017
rect 14645 32008 14657 32011
rect 14424 31980 14657 32008
rect 14424 31968 14430 31980
rect 14645 31977 14657 31980
rect 14691 31977 14703 32011
rect 14645 31971 14703 31977
rect 14734 31968 14740 32020
rect 14792 32008 14798 32020
rect 19659 32011 19717 32017
rect 14792 31980 19196 32008
rect 14792 31968 14798 31980
rect 13817 31943 13875 31949
rect 13817 31909 13829 31943
rect 13863 31940 13875 31943
rect 15473 31943 15531 31949
rect 15473 31940 15485 31943
rect 13863 31912 15485 31940
rect 13863 31909 13875 31912
rect 13817 31903 13875 31909
rect 15473 31909 15485 31912
rect 15519 31940 15531 31943
rect 15562 31940 15568 31952
rect 15519 31912 15568 31940
rect 15519 31909 15531 31912
rect 15473 31903 15531 31909
rect 15562 31900 15568 31912
rect 15620 31900 15626 31952
rect 18046 31940 18052 31952
rect 17959 31912 18052 31940
rect 18046 31900 18052 31912
rect 18104 31940 18110 31952
rect 18966 31940 18972 31952
rect 18104 31912 18972 31940
rect 18104 31900 18110 31912
rect 18966 31900 18972 31912
rect 19024 31900 19030 31952
rect 16850 31872 16856 31884
rect 16811 31844 16856 31872
rect 16850 31832 16856 31844
rect 16908 31832 16914 31884
rect 13722 31804 13728 31816
rect 13683 31776 13728 31804
rect 13722 31764 13728 31776
rect 13780 31764 13786 31816
rect 14366 31804 14372 31816
rect 14327 31776 14372 31804
rect 14366 31764 14372 31776
rect 14424 31764 14430 31816
rect 15378 31804 15384 31816
rect 15339 31776 15384 31804
rect 15378 31764 15384 31776
rect 15436 31764 15442 31816
rect 16991 31807 17049 31813
rect 16991 31773 17003 31807
rect 17037 31804 17049 31807
rect 17678 31804 17684 31816
rect 17037 31776 17684 31804
rect 17037 31773 17049 31776
rect 16991 31767 17049 31773
rect 17678 31764 17684 31776
rect 17736 31804 17742 31816
rect 17957 31807 18015 31813
rect 17957 31804 17969 31807
rect 17736 31776 17969 31804
rect 17736 31764 17742 31776
rect 17957 31773 17969 31776
rect 18003 31773 18015 31807
rect 18230 31804 18236 31816
rect 18191 31776 18236 31804
rect 17957 31767 18015 31773
rect 18230 31764 18236 31776
rect 18288 31804 18294 31816
rect 18874 31804 18880 31816
rect 18288 31776 18880 31804
rect 18288 31764 18294 31776
rect 18874 31764 18880 31776
rect 18932 31764 18938 31816
rect 19168 31804 19196 31980
rect 19659 31977 19671 32011
rect 19705 32008 19717 32011
rect 20254 32008 20260 32020
rect 19705 31980 20260 32008
rect 19705 31977 19717 31980
rect 19659 31971 19717 31977
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 21910 32008 21916 32020
rect 21871 31980 21916 32008
rect 21910 31968 21916 31980
rect 21968 31968 21974 32020
rect 27430 31968 27436 32020
rect 27488 32008 27494 32020
rect 27709 32011 27767 32017
rect 27709 32008 27721 32011
rect 27488 31980 27721 32008
rect 27488 31968 27494 31980
rect 27709 31977 27721 31980
rect 27755 31977 27767 32011
rect 27709 31971 27767 31977
rect 28721 32011 28779 32017
rect 28721 31977 28733 32011
rect 28767 32008 28779 32011
rect 29270 32008 29276 32020
rect 28767 31980 29276 32008
rect 28767 31977 28779 31980
rect 28721 31971 28779 31977
rect 29270 31968 29276 31980
rect 29328 31968 29334 32020
rect 30558 32008 30564 32020
rect 30519 31980 30564 32008
rect 30558 31968 30564 31980
rect 30616 31968 30622 32020
rect 31754 31968 31760 32020
rect 31812 32008 31818 32020
rect 31849 32011 31907 32017
rect 31849 32008 31861 32011
rect 31812 31980 31861 32008
rect 31812 31968 31818 31980
rect 31849 31977 31861 31980
rect 31895 32008 31907 32011
rect 33229 32011 33287 32017
rect 33229 32008 33241 32011
rect 31895 31980 32168 32008
rect 31895 31977 31907 31980
rect 31849 31971 31907 31977
rect 32140 31952 32168 31980
rect 33106 31980 33241 32008
rect 19886 31900 19892 31952
rect 19944 31940 19950 31952
rect 21085 31943 21143 31949
rect 21085 31940 21097 31943
rect 19944 31912 21097 31940
rect 19944 31900 19950 31912
rect 21085 31909 21097 31912
rect 21131 31909 21143 31943
rect 21634 31940 21640 31952
rect 21595 31912 21640 31940
rect 21085 31903 21143 31909
rect 21634 31900 21640 31912
rect 21692 31900 21698 31952
rect 24578 31900 24584 31952
rect 24636 31940 24642 31952
rect 25041 31943 25099 31949
rect 25041 31940 25053 31943
rect 24636 31912 25053 31940
rect 24636 31900 24642 31912
rect 25041 31909 25053 31912
rect 25087 31940 25099 31943
rect 25406 31940 25412 31952
rect 25087 31912 25412 31940
rect 25087 31909 25099 31912
rect 25041 31903 25099 31909
rect 25406 31900 25412 31912
rect 25464 31940 25470 31952
rect 27249 31943 27307 31949
rect 25464 31912 27200 31940
rect 25464 31900 25470 31912
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19588 31875 19646 31881
rect 19588 31872 19600 31875
rect 19484 31844 19600 31872
rect 19484 31832 19490 31844
rect 19588 31841 19600 31844
rect 19634 31872 19646 31875
rect 19978 31872 19984 31884
rect 19634 31844 19984 31872
rect 19634 31841 19646 31844
rect 19588 31835 19646 31841
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 23014 31872 23020 31884
rect 22975 31844 23020 31872
rect 23014 31832 23020 31844
rect 23072 31832 23078 31884
rect 23198 31872 23204 31884
rect 23159 31844 23204 31872
rect 23198 31832 23204 31844
rect 23256 31832 23262 31884
rect 27172 31872 27200 31912
rect 27249 31909 27261 31943
rect 27295 31940 27307 31943
rect 28074 31940 28080 31952
rect 27295 31912 28080 31940
rect 27295 31909 27307 31912
rect 27249 31903 27307 31909
rect 28074 31900 28080 31912
rect 28132 31900 28138 31952
rect 28353 31943 28411 31949
rect 28353 31909 28365 31943
rect 28399 31940 28411 31943
rect 28534 31940 28540 31952
rect 28399 31912 28540 31940
rect 28399 31909 28411 31912
rect 28353 31903 28411 31909
rect 28534 31900 28540 31912
rect 28592 31940 28598 31952
rect 30883 31943 30941 31949
rect 30883 31940 30895 31943
rect 28592 31912 30895 31940
rect 28592 31900 28598 31912
rect 30883 31909 30895 31912
rect 30929 31909 30941 31943
rect 32122 31940 32128 31952
rect 32035 31912 32128 31940
rect 30883 31903 30941 31909
rect 32122 31900 32128 31912
rect 32180 31900 32186 31952
rect 32306 31900 32312 31952
rect 32364 31940 32370 31952
rect 33106 31940 33134 31980
rect 33229 31977 33241 31980
rect 33275 32008 33287 32011
rect 33778 32008 33784 32020
rect 33275 31980 33784 32008
rect 33275 31977 33287 31980
rect 33229 31971 33287 31977
rect 33778 31968 33784 31980
rect 33836 31968 33842 32020
rect 34425 32011 34483 32017
rect 34425 31977 34437 32011
rect 34471 32008 34483 32011
rect 34882 32008 34888 32020
rect 34471 31980 34888 32008
rect 34471 31977 34483 31980
rect 34425 31971 34483 31977
rect 33686 31940 33692 31952
rect 32364 31912 33134 31940
rect 33647 31912 33692 31940
rect 32364 31900 32370 31912
rect 33686 31900 33692 31912
rect 33744 31900 33750 31952
rect 27522 31872 27528 31884
rect 27172 31844 27528 31872
rect 27522 31832 27528 31844
rect 27580 31832 27586 31884
rect 28626 31832 28632 31884
rect 28684 31872 28690 31884
rect 29181 31875 29239 31881
rect 29181 31872 29193 31875
rect 28684 31844 29193 31872
rect 28684 31832 28690 31844
rect 29181 31841 29193 31844
rect 29227 31841 29239 31875
rect 29181 31835 29239 31841
rect 29733 31875 29791 31881
rect 29733 31841 29745 31875
rect 29779 31872 29791 31875
rect 30006 31872 30012 31884
rect 29779 31844 30012 31872
rect 29779 31841 29791 31844
rect 29733 31835 29791 31841
rect 30006 31832 30012 31844
rect 30064 31872 30070 31884
rect 30558 31872 30564 31884
rect 30064 31844 30564 31872
rect 30064 31832 30070 31844
rect 30558 31832 30564 31844
rect 30616 31832 30622 31884
rect 30742 31872 30748 31884
rect 30703 31844 30748 31872
rect 30742 31832 30748 31844
rect 30800 31872 30806 31884
rect 32030 31872 32036 31884
rect 30800 31844 32036 31872
rect 30800 31832 30806 31844
rect 32030 31832 32036 31844
rect 32088 31832 32094 31884
rect 32140 31872 32168 31900
rect 32140 31844 32628 31872
rect 20993 31807 21051 31813
rect 20993 31804 21005 31807
rect 19168 31776 21005 31804
rect 20993 31773 21005 31776
rect 21039 31804 21051 31807
rect 21726 31804 21732 31816
rect 21039 31776 21732 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21726 31764 21732 31776
rect 21784 31764 21790 31816
rect 23290 31804 23296 31816
rect 23251 31776 23296 31804
rect 23290 31764 23296 31776
rect 23348 31764 23354 31816
rect 24026 31764 24032 31816
rect 24084 31804 24090 31816
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 24084 31776 24961 31804
rect 24084 31764 24090 31776
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25593 31807 25651 31813
rect 25593 31773 25605 31807
rect 25639 31804 25651 31807
rect 26878 31804 26884 31816
rect 25639 31776 26884 31804
rect 25639 31773 25651 31776
rect 25593 31767 25651 31773
rect 26878 31764 26884 31776
rect 26936 31764 26942 31816
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 32306 31813 32312 31816
rect 32272 31807 32312 31813
rect 32272 31804 32284 31807
rect 31076 31776 32284 31804
rect 31076 31764 31082 31776
rect 32272 31773 32284 31776
rect 32272 31767 32312 31773
rect 32306 31764 32312 31767
rect 32364 31764 32370 31816
rect 32398 31764 32404 31816
rect 32456 31804 32462 31816
rect 32493 31807 32551 31813
rect 32493 31804 32505 31807
rect 32456 31776 32505 31804
rect 32456 31764 32462 31776
rect 32493 31773 32505 31776
rect 32539 31773 32551 31807
rect 32600 31804 32628 31844
rect 34440 31804 34468 31971
rect 34882 31968 34888 31980
rect 34940 31968 34946 32020
rect 35802 31968 35808 32020
rect 35860 32008 35866 32020
rect 35897 32011 35955 32017
rect 35897 32008 35909 32011
rect 35860 31980 35909 32008
rect 35860 31968 35866 31980
rect 35897 31977 35909 31980
rect 35943 31977 35955 32011
rect 35897 31971 35955 31977
rect 35986 31968 35992 32020
rect 36044 32008 36050 32020
rect 37277 32011 37335 32017
rect 37277 32008 37289 32011
rect 36044 31980 37289 32008
rect 36044 31968 36050 31980
rect 37277 31977 37289 31980
rect 37323 31977 37335 32011
rect 37277 31971 37335 31977
rect 40681 32011 40739 32017
rect 40681 31977 40693 32011
rect 40727 32008 40739 32011
rect 41046 32008 41052 32020
rect 40727 31980 41052 32008
rect 40727 31977 40739 31980
rect 40681 31971 40739 31977
rect 41046 31968 41052 31980
rect 41104 31968 41110 32020
rect 42886 32008 42892 32020
rect 42847 31980 42892 32008
rect 42886 31968 42892 31980
rect 42944 31968 42950 32020
rect 44726 32008 44732 32020
rect 44687 31980 44732 32008
rect 44726 31968 44732 31980
rect 44784 31968 44790 32020
rect 46658 32008 46664 32020
rect 46619 31980 46664 32008
rect 46658 31968 46664 31980
rect 46716 31968 46722 32020
rect 36906 31940 36912 31952
rect 36867 31912 36912 31940
rect 36906 31900 36912 31912
rect 36964 31900 36970 31952
rect 38375 31943 38433 31949
rect 38375 31909 38387 31943
rect 38421 31940 38433 31943
rect 38654 31940 38660 31952
rect 38421 31912 38660 31940
rect 38421 31909 38433 31912
rect 38375 31903 38433 31909
rect 38654 31900 38660 31912
rect 38712 31940 38718 31952
rect 40082 31943 40140 31949
rect 40082 31940 40094 31943
rect 38712 31912 40094 31940
rect 38712 31900 38718 31912
rect 40082 31909 40094 31912
rect 40128 31940 40140 31943
rect 40402 31940 40408 31952
rect 40128 31912 40408 31940
rect 40128 31909 40140 31912
rect 40082 31903 40140 31909
rect 40402 31900 40408 31912
rect 40460 31900 40466 31952
rect 40494 31900 40500 31952
rect 40552 31940 40558 31952
rect 41598 31940 41604 31952
rect 40552 31912 41604 31940
rect 40552 31900 40558 31912
rect 41598 31900 41604 31912
rect 41656 31900 41662 31952
rect 41690 31900 41696 31952
rect 41748 31940 41754 31952
rect 41748 31912 41793 31940
rect 41748 31900 41754 31912
rect 42610 31900 42616 31952
rect 42668 31940 42674 31952
rect 43533 31943 43591 31949
rect 43533 31940 43545 31943
rect 42668 31912 43545 31940
rect 42668 31900 42674 31912
rect 43533 31909 43545 31912
rect 43579 31909 43591 31943
rect 43533 31903 43591 31909
rect 44085 31943 44143 31949
rect 44085 31909 44097 31943
rect 44131 31940 44143 31943
rect 45002 31940 45008 31952
rect 44131 31912 45008 31940
rect 44131 31909 44143 31912
rect 44085 31903 44143 31909
rect 45002 31900 45008 31912
rect 45060 31900 45066 31952
rect 45097 31943 45155 31949
rect 45097 31909 45109 31943
rect 45143 31940 45155 31943
rect 45186 31940 45192 31952
rect 45143 31912 45192 31940
rect 45143 31909 45155 31912
rect 45097 31903 45155 31909
rect 45186 31900 45192 31912
rect 45244 31940 45250 31952
rect 46109 31943 46167 31949
rect 46109 31940 46121 31943
rect 45244 31912 46121 31940
rect 45244 31900 45250 31912
rect 46109 31909 46121 31912
rect 46155 31909 46167 31943
rect 46109 31903 46167 31909
rect 34977 31875 35035 31881
rect 34977 31841 34989 31875
rect 35023 31841 35035 31875
rect 34977 31835 35035 31841
rect 32600 31776 34468 31804
rect 32493 31767 32551 31773
rect 34698 31764 34704 31816
rect 34756 31804 34762 31816
rect 34992 31804 35020 31835
rect 35894 31832 35900 31884
rect 35952 31872 35958 31884
rect 36262 31872 36268 31884
rect 35952 31844 36268 31872
rect 35952 31832 35958 31844
rect 36262 31832 36268 31844
rect 36320 31872 36326 31884
rect 36449 31875 36507 31881
rect 36449 31872 36461 31875
rect 36320 31844 36461 31872
rect 36320 31832 36326 31844
rect 36449 31841 36461 31844
rect 36495 31841 36507 31875
rect 36449 31835 36507 31841
rect 38013 31875 38071 31881
rect 38013 31841 38025 31875
rect 38059 31872 38071 31875
rect 38102 31872 38108 31884
rect 38059 31844 38108 31872
rect 38059 31841 38071 31844
rect 38013 31835 38071 31841
rect 38102 31832 38108 31844
rect 38160 31832 38166 31884
rect 46382 31872 46388 31884
rect 46343 31844 46388 31872
rect 46382 31832 46388 31844
rect 46440 31832 46446 31884
rect 35066 31804 35072 31816
rect 34756 31776 35072 31804
rect 34756 31764 34762 31776
rect 35066 31764 35072 31776
rect 35124 31764 35130 31816
rect 35253 31807 35311 31813
rect 35253 31773 35265 31807
rect 35299 31804 35311 31807
rect 37274 31804 37280 31816
rect 35299 31776 37280 31804
rect 35299 31773 35311 31776
rect 35253 31767 35311 31773
rect 15105 31739 15163 31745
rect 15105 31705 15117 31739
rect 15151 31736 15163 31739
rect 15654 31736 15660 31748
rect 15151 31708 15660 31736
rect 15151 31705 15163 31708
rect 15105 31699 15163 31705
rect 15654 31696 15660 31708
rect 15712 31736 15718 31748
rect 15933 31739 15991 31745
rect 15933 31736 15945 31739
rect 15712 31708 15945 31736
rect 15712 31696 15718 31708
rect 15933 31705 15945 31708
rect 15979 31736 15991 31739
rect 31573 31739 31631 31745
rect 15979 31708 18092 31736
rect 15979 31705 15991 31708
rect 15933 31699 15991 31705
rect 14642 31628 14648 31680
rect 14700 31668 14706 31680
rect 15286 31668 15292 31680
rect 14700 31640 15292 31668
rect 14700 31628 14706 31640
rect 15286 31628 15292 31640
rect 15344 31628 15350 31680
rect 16298 31668 16304 31680
rect 16259 31640 16304 31668
rect 16298 31628 16304 31640
rect 16356 31628 16362 31680
rect 18064 31668 18092 31708
rect 31573 31705 31585 31739
rect 31619 31736 31631 31739
rect 31938 31736 31944 31748
rect 31619 31708 31944 31736
rect 31619 31705 31631 31708
rect 31573 31699 31631 31705
rect 31938 31696 31944 31708
rect 31996 31696 32002 31748
rect 32030 31696 32036 31748
rect 32088 31736 32094 31748
rect 32585 31739 32643 31745
rect 32585 31736 32597 31739
rect 32088 31708 32597 31736
rect 32088 31696 32094 31708
rect 32585 31705 32597 31708
rect 32631 31705 32643 31739
rect 32585 31699 32643 31705
rect 33594 31696 33600 31748
rect 33652 31736 33658 31748
rect 34054 31736 34060 31748
rect 33652 31708 34060 31736
rect 33652 31696 33658 31708
rect 34054 31696 34060 31708
rect 34112 31736 34118 31748
rect 35268 31736 35296 31767
rect 37274 31764 37280 31776
rect 37332 31764 37338 31816
rect 39758 31804 39764 31816
rect 39719 31776 39764 31804
rect 39758 31764 39764 31776
rect 39816 31764 39822 31816
rect 41874 31804 41880 31816
rect 41835 31776 41880 31804
rect 41874 31764 41880 31776
rect 41932 31804 41938 31816
rect 41932 31776 42794 31804
rect 41932 31764 41938 31776
rect 34112 31708 35296 31736
rect 34112 31696 34118 31708
rect 35434 31696 35440 31748
rect 35492 31736 35498 31748
rect 36633 31739 36691 31745
rect 35492 31708 36400 31736
rect 35492 31696 35498 31708
rect 18782 31668 18788 31680
rect 18064 31640 18788 31668
rect 18782 31628 18788 31640
rect 18840 31628 18846 31680
rect 24394 31668 24400 31680
rect 24355 31640 24400 31668
rect 24394 31628 24400 31640
rect 24452 31628 24458 31680
rect 28350 31628 28356 31680
rect 28408 31668 28414 31680
rect 29089 31671 29147 31677
rect 29089 31668 29101 31671
rect 28408 31640 29101 31668
rect 28408 31628 28414 31640
rect 29089 31637 29101 31640
rect 29135 31668 29147 31671
rect 29730 31668 29736 31680
rect 29135 31640 29736 31668
rect 29135 31637 29147 31640
rect 29089 31631 29147 31637
rect 29730 31628 29736 31640
rect 29788 31628 29794 31680
rect 30282 31668 30288 31680
rect 30243 31640 30288 31668
rect 30282 31628 30288 31640
rect 30340 31628 30346 31680
rect 32401 31671 32459 31677
rect 32401 31637 32413 31671
rect 32447 31668 32459 31671
rect 32490 31668 32496 31680
rect 32447 31640 32496 31668
rect 32447 31637 32459 31640
rect 32401 31631 32459 31637
rect 32490 31628 32496 31640
rect 32548 31628 32554 31680
rect 35526 31668 35532 31680
rect 35487 31640 35532 31668
rect 35526 31628 35532 31640
rect 35584 31628 35590 31680
rect 36372 31677 36400 31708
rect 36633 31705 36645 31739
rect 36679 31736 36691 31739
rect 36906 31736 36912 31748
rect 36679 31708 36912 31736
rect 36679 31705 36691 31708
rect 36633 31699 36691 31705
rect 36906 31696 36912 31708
rect 36964 31696 36970 31748
rect 38933 31739 38991 31745
rect 38933 31705 38945 31739
rect 38979 31736 38991 31739
rect 41690 31736 41696 31748
rect 38979 31708 41696 31736
rect 38979 31705 38991 31708
rect 38933 31699 38991 31705
rect 41690 31696 41696 31708
rect 41748 31696 41754 31748
rect 42766 31736 42794 31776
rect 43162 31764 43168 31816
rect 43220 31804 43226 31816
rect 43441 31807 43499 31813
rect 43441 31804 43453 31807
rect 43220 31776 43453 31804
rect 43220 31764 43226 31776
rect 43441 31773 43453 31776
rect 43487 31773 43499 31807
rect 43441 31767 43499 31773
rect 45005 31807 45063 31813
rect 45005 31773 45017 31807
rect 45051 31804 45063 31807
rect 45830 31804 45836 31816
rect 45051 31776 45836 31804
rect 45051 31773 45063 31776
rect 45005 31767 45063 31773
rect 45830 31764 45836 31776
rect 45888 31764 45894 31816
rect 44910 31736 44916 31748
rect 42766 31708 44916 31736
rect 44910 31696 44916 31708
rect 44968 31736 44974 31748
rect 45557 31739 45615 31745
rect 45557 31736 45569 31739
rect 44968 31708 45569 31736
rect 44968 31696 44974 31708
rect 45557 31705 45569 31708
rect 45603 31705 45615 31739
rect 45557 31699 45615 31705
rect 36357 31671 36415 31677
rect 36357 31637 36369 31671
rect 36403 31668 36415 31671
rect 37734 31668 37740 31680
rect 36403 31640 37740 31668
rect 36403 31637 36415 31640
rect 36357 31631 36415 31637
rect 37734 31628 37740 31640
rect 37792 31628 37798 31680
rect 1104 31578 48852 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 48852 31578
rect 1104 31504 48852 31526
rect 13722 31473 13728 31476
rect 13449 31467 13507 31473
rect 13449 31433 13461 31467
rect 13495 31464 13507 31467
rect 13679 31467 13728 31473
rect 13679 31464 13691 31467
rect 13495 31436 13691 31464
rect 13495 31433 13507 31436
rect 13449 31427 13507 31433
rect 13679 31433 13691 31436
rect 13725 31433 13728 31467
rect 13679 31427 13728 31433
rect 13722 31424 13728 31427
rect 13780 31424 13786 31476
rect 14691 31467 14749 31473
rect 14691 31433 14703 31467
rect 14737 31464 14749 31467
rect 15378 31464 15384 31476
rect 14737 31436 15384 31464
rect 14737 31433 14749 31436
rect 14691 31427 14749 31433
rect 15378 31424 15384 31436
rect 15436 31424 15442 31476
rect 15473 31467 15531 31473
rect 15473 31433 15485 31467
rect 15519 31464 15531 31467
rect 15562 31464 15568 31476
rect 15519 31436 15568 31464
rect 15519 31433 15531 31436
rect 15473 31427 15531 31433
rect 14461 31399 14519 31405
rect 14461 31365 14473 31399
rect 14507 31396 14519 31399
rect 15488 31396 15516 31427
rect 15562 31424 15568 31436
rect 15620 31424 15626 31476
rect 17497 31467 17555 31473
rect 17497 31433 17509 31467
rect 17543 31464 17555 31467
rect 17865 31467 17923 31473
rect 17865 31464 17877 31467
rect 17543 31436 17877 31464
rect 17543 31433 17555 31436
rect 17497 31427 17555 31433
rect 17865 31433 17877 31436
rect 17911 31464 17923 31467
rect 18046 31464 18052 31476
rect 17911 31436 18052 31464
rect 17911 31433 17923 31436
rect 17865 31427 17923 31433
rect 18046 31424 18052 31436
rect 18104 31424 18110 31476
rect 19886 31424 19892 31476
rect 19944 31464 19950 31476
rect 20073 31467 20131 31473
rect 20073 31464 20085 31467
rect 19944 31436 20085 31464
rect 19944 31424 19950 31436
rect 20073 31433 20085 31436
rect 20119 31464 20131 31467
rect 20165 31467 20223 31473
rect 20165 31464 20177 31467
rect 20119 31436 20177 31464
rect 20119 31433 20131 31436
rect 20073 31427 20131 31433
rect 20165 31433 20177 31436
rect 20211 31433 20223 31467
rect 21726 31464 21732 31476
rect 21687 31436 21732 31464
rect 20165 31427 20223 31433
rect 21726 31424 21732 31436
rect 21784 31424 21790 31476
rect 22695 31467 22753 31473
rect 22695 31433 22707 31467
rect 22741 31464 22753 31467
rect 24394 31464 24400 31476
rect 22741 31436 24400 31464
rect 22741 31433 22753 31436
rect 22695 31427 22753 31433
rect 24394 31424 24400 31436
rect 24452 31424 24458 31476
rect 25406 31424 25412 31476
rect 25464 31464 25470 31476
rect 25501 31467 25559 31473
rect 25501 31464 25513 31467
rect 25464 31436 25513 31464
rect 25464 31424 25470 31436
rect 25501 31433 25513 31436
rect 25547 31433 25559 31467
rect 25501 31427 25559 31433
rect 27430 31424 27436 31476
rect 27488 31464 27494 31476
rect 27847 31467 27905 31473
rect 27847 31464 27859 31467
rect 27488 31436 27859 31464
rect 27488 31424 27494 31436
rect 27847 31433 27859 31436
rect 27893 31433 27905 31467
rect 27847 31427 27905 31433
rect 31481 31467 31539 31473
rect 31481 31433 31493 31467
rect 31527 31464 31539 31467
rect 31527 31436 31892 31464
rect 31527 31433 31539 31436
rect 31481 31427 31539 31433
rect 14507 31368 15516 31396
rect 14507 31365 14519 31368
rect 14461 31359 14519 31365
rect 16850 31356 16856 31408
rect 16908 31396 16914 31408
rect 16945 31399 17003 31405
rect 16945 31396 16957 31399
rect 16908 31368 16957 31396
rect 16908 31356 16914 31368
rect 16945 31365 16957 31368
rect 16991 31396 17003 31399
rect 19426 31396 19432 31408
rect 16991 31368 19432 31396
rect 16991 31365 17003 31368
rect 16945 31359 17003 31365
rect 19426 31356 19432 31368
rect 19484 31356 19490 31408
rect 20438 31356 20444 31408
rect 20496 31396 20502 31408
rect 24026 31396 24032 31408
rect 20496 31368 24032 31396
rect 20496 31356 20502 31368
rect 24026 31356 24032 31368
rect 24084 31356 24090 31408
rect 27985 31399 28043 31405
rect 27985 31365 27997 31399
rect 28031 31396 28043 31399
rect 28258 31396 28264 31408
rect 28031 31368 28264 31396
rect 28031 31365 28043 31368
rect 27985 31359 28043 31365
rect 28258 31356 28264 31368
rect 28316 31396 28322 31408
rect 30190 31396 30196 31408
rect 28316 31368 30196 31396
rect 28316 31356 28322 31368
rect 30190 31356 30196 31368
rect 30248 31356 30254 31408
rect 31864 31405 31892 31436
rect 34330 31424 34336 31476
rect 34388 31464 34394 31476
rect 34609 31467 34667 31473
rect 34609 31464 34621 31467
rect 34388 31436 34621 31464
rect 34388 31424 34394 31436
rect 34609 31433 34621 31436
rect 34655 31464 34667 31467
rect 34698 31464 34704 31476
rect 34655 31436 34704 31464
rect 34655 31433 34667 31436
rect 34609 31427 34667 31433
rect 34698 31424 34704 31436
rect 34756 31424 34762 31476
rect 34790 31424 34796 31476
rect 34848 31464 34854 31476
rect 35069 31467 35127 31473
rect 35069 31464 35081 31467
rect 34848 31436 35081 31464
rect 34848 31424 34854 31436
rect 35069 31433 35081 31436
rect 35115 31433 35127 31467
rect 35069 31427 35127 31433
rect 35342 31424 35348 31476
rect 35400 31464 35406 31476
rect 35713 31467 35771 31473
rect 35713 31464 35725 31467
rect 35400 31436 35725 31464
rect 35400 31424 35406 31436
rect 35713 31433 35725 31436
rect 35759 31433 35771 31467
rect 36262 31464 36268 31476
rect 36223 31436 36268 31464
rect 35713 31427 35771 31433
rect 36262 31424 36268 31436
rect 36320 31424 36326 31476
rect 38102 31424 38108 31476
rect 38160 31464 38166 31476
rect 39393 31467 39451 31473
rect 39393 31464 39405 31467
rect 38160 31436 39405 31464
rect 38160 31424 38166 31436
rect 39393 31433 39405 31436
rect 39439 31433 39451 31467
rect 39393 31427 39451 31433
rect 40957 31467 41015 31473
rect 40957 31433 40969 31467
rect 41003 31464 41015 31467
rect 41046 31464 41052 31476
rect 41003 31436 41052 31464
rect 41003 31433 41015 31436
rect 40957 31427 41015 31433
rect 41046 31424 41052 31436
rect 41104 31424 41110 31476
rect 41690 31424 41696 31476
rect 41748 31464 41754 31476
rect 42061 31467 42119 31473
rect 42061 31464 42073 31467
rect 41748 31436 42073 31464
rect 41748 31424 41754 31436
rect 42061 31433 42073 31436
rect 42107 31433 42119 31467
rect 42061 31427 42119 31433
rect 42521 31467 42579 31473
rect 42521 31433 42533 31467
rect 42567 31464 42579 31467
rect 43162 31464 43168 31476
rect 42567 31436 43168 31464
rect 42567 31433 42579 31436
rect 42521 31427 42579 31433
rect 31849 31399 31907 31405
rect 31849 31365 31861 31399
rect 31895 31396 31907 31399
rect 32582 31396 32588 31408
rect 31895 31368 32588 31396
rect 31895 31365 31907 31368
rect 31849 31359 31907 31365
rect 32582 31356 32588 31368
rect 32640 31356 32646 31408
rect 42076 31396 42104 31427
rect 43162 31424 43168 31436
rect 43220 31424 43226 31476
rect 45186 31424 45192 31476
rect 45244 31464 45250 31476
rect 45373 31467 45431 31473
rect 45373 31464 45385 31467
rect 45244 31436 45385 31464
rect 45244 31424 45250 31436
rect 45373 31433 45385 31436
rect 45419 31433 45431 31467
rect 45830 31464 45836 31476
rect 45791 31436 45836 31464
rect 45373 31427 45431 31433
rect 45830 31424 45836 31436
rect 45888 31424 45894 31476
rect 42610 31396 42616 31408
rect 42076 31368 42616 31396
rect 42610 31356 42616 31368
rect 42668 31396 42674 31408
rect 42797 31399 42855 31405
rect 42797 31396 42809 31399
rect 42668 31368 42809 31396
rect 42668 31356 42674 31368
rect 42797 31365 42809 31368
rect 42843 31365 42855 31399
rect 42797 31359 42855 31365
rect 15010 31328 15016 31340
rect 14635 31300 15016 31328
rect 14635 31269 14663 31300
rect 15010 31288 15016 31300
rect 15068 31328 15074 31340
rect 15105 31331 15163 31337
rect 15105 31328 15117 31331
rect 15068 31300 15117 31328
rect 15068 31288 15074 31300
rect 15105 31297 15117 31300
rect 15151 31328 15163 31331
rect 15194 31328 15200 31340
rect 15151 31300 15200 31328
rect 15151 31297 15163 31300
rect 15105 31291 15163 31297
rect 15194 31288 15200 31300
rect 15252 31288 15258 31340
rect 15654 31328 15660 31340
rect 15615 31300 15660 31328
rect 15654 31288 15660 31300
rect 15712 31288 15718 31340
rect 17310 31288 17316 31340
rect 17368 31328 17374 31340
rect 18141 31331 18199 31337
rect 18141 31328 18153 31331
rect 17368 31300 18153 31328
rect 17368 31288 17374 31300
rect 18141 31297 18153 31300
rect 18187 31328 18199 31331
rect 19061 31331 19119 31337
rect 19061 31328 19073 31331
rect 18187 31300 19073 31328
rect 18187 31297 18199 31300
rect 18141 31291 18199 31297
rect 19061 31297 19073 31300
rect 19107 31297 19119 31331
rect 21634 31328 21640 31340
rect 19061 31291 19119 31297
rect 20174 31300 21640 31328
rect 13608 31263 13666 31269
rect 13608 31229 13620 31263
rect 13654 31260 13666 31263
rect 14620 31263 14678 31269
rect 13654 31232 13814 31260
rect 13654 31229 13666 31232
rect 13608 31223 13666 31229
rect 13786 31124 13814 31232
rect 14620 31229 14632 31263
rect 14666 31229 14678 31263
rect 14620 31223 14678 31229
rect 18782 31220 18788 31272
rect 18840 31260 18846 31272
rect 20174 31260 20202 31300
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 22465 31331 22523 31337
rect 22465 31297 22477 31331
rect 22511 31328 22523 31331
rect 23198 31328 23204 31340
rect 22511 31300 23204 31328
rect 22511 31297 22523 31300
rect 22465 31291 22523 31297
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 24762 31288 24768 31340
rect 24820 31328 24826 31340
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 24820 31300 24869 31328
rect 24820 31288 24826 31300
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 28997 31331 29055 31337
rect 28997 31328 29009 31331
rect 25004 31300 29009 31328
rect 25004 31288 25010 31300
rect 28997 31297 29009 31300
rect 29043 31328 29055 31331
rect 31938 31328 31944 31340
rect 29043 31300 29316 31328
rect 31899 31300 31944 31328
rect 29043 31297 29055 31300
rect 28997 31291 29055 31297
rect 18840 31232 20202 31260
rect 18840 31220 18846 31232
rect 22278 31220 22284 31272
rect 22336 31260 22342 31272
rect 22592 31263 22650 31269
rect 22592 31260 22604 31263
rect 22336 31232 22604 31260
rect 22336 31220 22342 31232
rect 22592 31229 22604 31232
rect 22638 31229 22650 31263
rect 22592 31223 22650 31229
rect 15749 31195 15807 31201
rect 15749 31161 15761 31195
rect 15795 31192 15807 31195
rect 16114 31192 16120 31204
rect 15795 31164 16120 31192
rect 15795 31161 15807 31164
rect 15749 31155 15807 31161
rect 16114 31152 16120 31164
rect 16172 31152 16178 31204
rect 16301 31195 16359 31201
rect 16301 31161 16313 31195
rect 16347 31192 16359 31195
rect 16482 31192 16488 31204
rect 16347 31164 16488 31192
rect 16347 31161 16359 31164
rect 16301 31155 16359 31161
rect 16482 31152 16488 31164
rect 16540 31152 16546 31204
rect 18233 31195 18291 31201
rect 18233 31161 18245 31195
rect 18279 31161 18291 31195
rect 18233 31155 18291 31161
rect 14093 31127 14151 31133
rect 14093 31124 14105 31127
rect 13786 31096 14105 31124
rect 14093 31093 14105 31096
rect 14139 31124 14151 31127
rect 14734 31124 14740 31136
rect 14139 31096 14740 31124
rect 14139 31093 14151 31096
rect 14093 31087 14151 31093
rect 14734 31084 14740 31096
rect 14792 31084 14798 31136
rect 18046 31084 18052 31136
rect 18104 31124 18110 31136
rect 18248 31124 18276 31155
rect 20254 31152 20260 31204
rect 20312 31192 20318 31204
rect 20441 31195 20499 31201
rect 20441 31192 20453 31195
rect 20312 31164 20453 31192
rect 20312 31152 20318 31164
rect 20441 31161 20453 31164
rect 20487 31161 20499 31195
rect 20441 31155 20499 31161
rect 20533 31195 20591 31201
rect 20533 31161 20545 31195
rect 20579 31161 20591 31195
rect 20533 31155 20591 31161
rect 21085 31195 21143 31201
rect 21085 31161 21097 31195
rect 21131 31192 21143 31195
rect 21266 31192 21272 31204
rect 21131 31164 21272 31192
rect 21131 31161 21143 31164
rect 21085 31155 21143 31161
rect 18104 31096 18276 31124
rect 19613 31127 19671 31133
rect 18104 31084 18110 31096
rect 19613 31093 19625 31127
rect 19659 31124 19671 31127
rect 19978 31124 19984 31136
rect 19659 31096 19984 31124
rect 19659 31093 19671 31096
rect 19613 31087 19671 31093
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 20073 31127 20131 31133
rect 20073 31093 20085 31127
rect 20119 31124 20131 31127
rect 20548 31124 20576 31155
rect 21266 31152 21272 31164
rect 21324 31152 21330 31204
rect 22607 31192 22635 31223
rect 23014 31220 23020 31272
rect 23072 31260 23078 31272
rect 23477 31263 23535 31269
rect 23477 31260 23489 31263
rect 23072 31232 23489 31260
rect 23072 31220 23078 31232
rect 23477 31229 23489 31232
rect 23523 31260 23535 31263
rect 23934 31260 23940 31272
rect 23523 31232 23940 31260
rect 23523 31229 23535 31232
rect 23477 31223 23535 31229
rect 23934 31220 23940 31232
rect 23992 31220 23998 31272
rect 29288 31269 29316 31300
rect 31938 31288 31944 31300
rect 31996 31288 32002 31340
rect 37826 31328 37832 31340
rect 37200 31300 37832 31328
rect 37200 31272 37228 31300
rect 37826 31288 37832 31300
rect 37884 31288 37890 31340
rect 39117 31331 39175 31337
rect 39117 31297 39129 31331
rect 39163 31328 39175 31331
rect 39758 31328 39764 31340
rect 39163 31300 39764 31328
rect 39163 31297 39175 31300
rect 39117 31291 39175 31297
rect 39758 31288 39764 31300
rect 39816 31328 39822 31340
rect 40129 31331 40187 31337
rect 40129 31328 40141 31331
rect 39816 31300 40141 31328
rect 39816 31288 39822 31300
rect 40129 31297 40141 31300
rect 40175 31297 40187 31331
rect 40129 31291 40187 31297
rect 40586 31288 40592 31340
rect 40644 31328 40650 31340
rect 41138 31328 41144 31340
rect 40644 31300 41144 31328
rect 40644 31288 40650 31300
rect 41138 31288 41144 31300
rect 41196 31288 41202 31340
rect 27776 31263 27834 31269
rect 27776 31229 27788 31263
rect 27822 31260 27834 31263
rect 27985 31263 28043 31269
rect 27985 31260 27997 31263
rect 27822 31232 27997 31260
rect 27822 31229 27834 31232
rect 27776 31223 27834 31229
rect 27985 31229 27997 31232
rect 28031 31229 28043 31263
rect 27985 31223 28043 31229
rect 29273 31263 29331 31269
rect 29273 31229 29285 31263
rect 29319 31229 29331 31263
rect 29730 31260 29736 31272
rect 29691 31232 29736 31260
rect 29273 31223 29331 31229
rect 29730 31220 29736 31232
rect 29788 31220 29794 31272
rect 31720 31263 31778 31269
rect 31720 31260 31732 31263
rect 30484 31232 31732 31260
rect 23109 31195 23167 31201
rect 23109 31192 23121 31195
rect 22607 31164 23121 31192
rect 23109 31161 23121 31164
rect 23155 31161 23167 31195
rect 24578 31192 24584 31204
rect 24539 31164 24584 31192
rect 23109 31155 23167 31161
rect 24578 31152 24584 31164
rect 24636 31152 24642 31204
rect 24682 31195 24740 31201
rect 24682 31161 24694 31195
rect 24728 31192 24740 31195
rect 25682 31192 25688 31204
rect 24728 31164 25688 31192
rect 24728 31161 24740 31164
rect 24682 31155 24740 31161
rect 25682 31152 25688 31164
rect 25740 31192 25746 31204
rect 25961 31195 26019 31201
rect 25961 31192 25973 31195
rect 25740 31164 25973 31192
rect 25740 31152 25746 31164
rect 25961 31161 25973 31164
rect 26007 31161 26019 31195
rect 26234 31192 26240 31204
rect 26195 31164 26240 31192
rect 25961 31155 26019 31161
rect 21174 31124 21180 31136
rect 20119 31096 21180 31124
rect 20119 31093 20131 31096
rect 20073 31087 20131 31093
rect 21174 31084 21180 31096
rect 21232 31124 21238 31136
rect 21361 31127 21419 31133
rect 21361 31124 21373 31127
rect 21232 31096 21373 31124
rect 21232 31084 21238 31096
rect 21361 31093 21373 31096
rect 21407 31093 21419 31127
rect 24394 31124 24400 31136
rect 24355 31096 24400 31124
rect 21361 31087 21419 31093
rect 24394 31084 24400 31096
rect 24452 31084 24458 31136
rect 25976 31124 26004 31155
rect 26234 31152 26240 31164
rect 26292 31152 26298 31204
rect 26329 31195 26387 31201
rect 26329 31161 26341 31195
rect 26375 31161 26387 31195
rect 26329 31155 26387 31161
rect 26881 31195 26939 31201
rect 26881 31161 26893 31195
rect 26927 31192 26939 31195
rect 28442 31192 28448 31204
rect 26927 31164 28448 31192
rect 26927 31161 26939 31164
rect 26881 31155 26939 31161
rect 26344 31124 26372 31155
rect 28442 31152 28448 31164
rect 28500 31152 28506 31204
rect 30484 31136 30512 31232
rect 31720 31229 31732 31232
rect 31766 31260 31778 31263
rect 31846 31260 31852 31272
rect 31766 31232 31852 31260
rect 31766 31229 31778 31232
rect 31720 31223 31778 31229
rect 31846 31220 31852 31232
rect 31904 31220 31910 31272
rect 33137 31263 33195 31269
rect 33137 31229 33149 31263
rect 33183 31260 33195 31263
rect 33873 31263 33931 31269
rect 33873 31260 33885 31263
rect 33183 31232 33885 31260
rect 33183 31229 33195 31232
rect 33137 31223 33195 31229
rect 33873 31229 33885 31232
rect 33919 31260 33931 31263
rect 34146 31260 34152 31272
rect 33919 31232 34152 31260
rect 33919 31229 33931 31232
rect 33873 31223 33931 31229
rect 31570 31192 31576 31204
rect 31531 31164 31576 31192
rect 31570 31152 31576 31164
rect 31628 31152 31634 31204
rect 26694 31124 26700 31136
rect 25976 31096 26700 31124
rect 26694 31084 26700 31096
rect 26752 31084 26758 31136
rect 28626 31124 28632 31136
rect 28587 31096 28632 31124
rect 28626 31084 28632 31096
rect 28684 31084 28690 31136
rect 29362 31124 29368 31136
rect 29323 31096 29368 31124
rect 29362 31084 29368 31096
rect 29420 31084 29426 31136
rect 30466 31124 30472 31136
rect 30427 31096 30472 31124
rect 30466 31084 30472 31096
rect 30524 31084 30530 31136
rect 30834 31124 30840 31136
rect 30795 31096 30840 31124
rect 30834 31084 30840 31096
rect 30892 31084 30898 31136
rect 32214 31124 32220 31136
rect 32175 31096 32220 31124
rect 32214 31084 32220 31096
rect 32272 31084 32278 31136
rect 32582 31124 32588 31136
rect 32543 31096 32588 31124
rect 32582 31084 32588 31096
rect 32640 31124 32646 31136
rect 33152 31124 33180 31223
rect 34146 31220 34152 31232
rect 34204 31220 34210 31272
rect 34698 31220 34704 31272
rect 34756 31260 34762 31272
rect 34885 31263 34943 31269
rect 34885 31260 34897 31263
rect 34756 31232 34897 31260
rect 34756 31220 34762 31232
rect 34885 31229 34897 31232
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 36725 31263 36783 31269
rect 36725 31229 36737 31263
rect 36771 31260 36783 31263
rect 37093 31263 37151 31269
rect 37093 31260 37105 31263
rect 36771 31232 37105 31260
rect 36771 31229 36783 31232
rect 36725 31223 36783 31229
rect 37093 31229 37105 31232
rect 37139 31260 37151 31263
rect 37182 31260 37188 31272
rect 37139 31232 37188 31260
rect 37139 31229 37151 31232
rect 37093 31223 37151 31229
rect 37182 31220 37188 31232
rect 37240 31220 37246 31272
rect 37369 31263 37427 31269
rect 37369 31229 37381 31263
rect 37415 31260 37427 31263
rect 37458 31260 37464 31272
rect 37415 31232 37464 31260
rect 37415 31229 37427 31232
rect 37369 31223 37427 31229
rect 37458 31220 37464 31232
rect 37516 31220 37522 31272
rect 38286 31220 38292 31272
rect 38344 31260 38350 31272
rect 38381 31263 38439 31269
rect 38381 31260 38393 31263
rect 38344 31232 38393 31260
rect 38344 31220 38350 31232
rect 38381 31229 38393 31232
rect 38427 31229 38439 31263
rect 38838 31260 38844 31272
rect 38799 31232 38844 31260
rect 38381 31223 38439 31229
rect 38838 31220 38844 31232
rect 38896 31220 38902 31272
rect 33965 31195 34023 31201
rect 33965 31161 33977 31195
rect 34011 31192 34023 31195
rect 35894 31192 35900 31204
rect 34011 31164 35900 31192
rect 34011 31161 34023 31164
rect 33965 31155 34023 31161
rect 35894 31152 35900 31164
rect 35952 31152 35958 31204
rect 37550 31192 37556 31204
rect 37511 31164 37556 31192
rect 37550 31152 37556 31164
rect 37608 31152 37614 31204
rect 41233 31195 41291 31201
rect 41233 31161 41245 31195
rect 41279 31161 41291 31195
rect 41233 31155 41291 31161
rect 41785 31195 41843 31201
rect 41785 31161 41797 31195
rect 41831 31192 41843 31195
rect 42058 31192 42064 31204
rect 41831 31164 42064 31192
rect 41831 31161 41843 31164
rect 41785 31155 41843 31161
rect 32640 31096 33180 31124
rect 32640 31084 32646 31096
rect 34698 31084 34704 31136
rect 34756 31124 34762 31136
rect 35345 31127 35403 31133
rect 35345 31124 35357 31127
rect 34756 31096 35357 31124
rect 34756 31084 34762 31096
rect 35345 31093 35357 31096
rect 35391 31093 35403 31127
rect 35345 31087 35403 31093
rect 38105 31127 38163 31133
rect 38105 31093 38117 31127
rect 38151 31124 38163 31127
rect 38654 31124 38660 31136
rect 38151 31096 38660 31124
rect 38151 31093 38163 31096
rect 38105 31087 38163 31093
rect 38654 31084 38660 31096
rect 38712 31124 38718 31136
rect 39761 31127 39819 31133
rect 39761 31124 39773 31127
rect 38712 31096 39773 31124
rect 38712 31084 38718 31096
rect 39761 31093 39773 31096
rect 39807 31093 39819 31127
rect 39761 31087 39819 31093
rect 41046 31084 41052 31136
rect 41104 31124 41110 31136
rect 41248 31124 41276 31155
rect 42058 31152 42064 31164
rect 42116 31152 42122 31204
rect 41104 31096 41276 31124
rect 42812 31124 42840 31359
rect 43898 31288 43904 31340
rect 43956 31328 43962 31340
rect 45278 31328 45284 31340
rect 43956 31300 45284 31328
rect 43956 31288 43962 31300
rect 45278 31288 45284 31300
rect 45336 31288 45342 31340
rect 44612 31263 44670 31269
rect 44612 31229 44624 31263
rect 44658 31260 44670 31263
rect 45005 31263 45063 31269
rect 45005 31260 45017 31263
rect 44658 31232 45017 31260
rect 44658 31229 44670 31232
rect 44612 31223 44670 31229
rect 45005 31229 45017 31232
rect 45051 31260 45063 31263
rect 45646 31260 45652 31272
rect 45051 31232 45652 31260
rect 45051 31229 45063 31232
rect 45005 31223 45063 31229
rect 45646 31220 45652 31232
rect 45704 31220 45710 31272
rect 46106 31260 46112 31272
rect 46067 31232 46112 31260
rect 46106 31220 46112 31232
rect 46164 31260 46170 31272
rect 46569 31263 46627 31269
rect 46569 31260 46581 31263
rect 46164 31232 46581 31260
rect 46164 31220 46170 31232
rect 46569 31229 46581 31232
rect 46615 31229 46627 31263
rect 46569 31223 46627 31229
rect 43070 31192 43076 31204
rect 43031 31164 43076 31192
rect 43070 31152 43076 31164
rect 43128 31152 43134 31204
rect 43165 31195 43223 31201
rect 43165 31161 43177 31195
rect 43211 31161 43223 31195
rect 43714 31192 43720 31204
rect 43627 31164 43720 31192
rect 43165 31155 43223 31161
rect 43180 31124 43208 31155
rect 43714 31152 43720 31164
rect 43772 31192 43778 31204
rect 45094 31192 45100 31204
rect 43772 31164 45100 31192
rect 43772 31152 43778 31164
rect 45094 31152 45100 31164
rect 45152 31152 45158 31204
rect 45278 31152 45284 31204
rect 45336 31192 45342 31204
rect 46382 31192 46388 31204
rect 45336 31164 46388 31192
rect 45336 31152 45342 31164
rect 46382 31152 46388 31164
rect 46440 31192 46446 31204
rect 46937 31195 46995 31201
rect 46937 31192 46949 31195
rect 46440 31164 46949 31192
rect 46440 31152 46446 31164
rect 46937 31161 46949 31164
rect 46983 31161 46995 31195
rect 46937 31155 46995 31161
rect 43993 31127 44051 31133
rect 43993 31124 44005 31127
rect 42812 31096 44005 31124
rect 41104 31084 41110 31096
rect 43993 31093 44005 31096
rect 44039 31093 44051 31127
rect 43993 31087 44051 31093
rect 44683 31127 44741 31133
rect 44683 31093 44695 31127
rect 44729 31124 44741 31127
rect 44818 31124 44824 31136
rect 44729 31096 44824 31124
rect 44729 31093 44741 31096
rect 44683 31087 44741 31093
rect 44818 31084 44824 31096
rect 44876 31084 44882 31136
rect 46290 31124 46296 31136
rect 46251 31096 46296 31124
rect 46290 31084 46296 31096
rect 46348 31084 46354 31136
rect 1104 31034 48852 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 48852 31034
rect 1104 30960 48852 30982
rect 15105 30923 15163 30929
rect 15105 30889 15117 30923
rect 15151 30920 15163 30923
rect 15378 30920 15384 30932
rect 15151 30892 15384 30920
rect 15151 30889 15163 30892
rect 15105 30883 15163 30889
rect 15378 30880 15384 30892
rect 15436 30880 15442 30932
rect 16209 30923 16267 30929
rect 16209 30889 16221 30923
rect 16255 30920 16267 30923
rect 16298 30920 16304 30932
rect 16255 30892 16304 30920
rect 16255 30889 16267 30892
rect 16209 30883 16267 30889
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 17678 30920 17684 30932
rect 17639 30892 17684 30920
rect 17678 30880 17684 30892
rect 17736 30880 17742 30932
rect 20162 30880 20168 30932
rect 20220 30920 20226 30932
rect 22278 30920 22284 30932
rect 20220 30892 22284 30920
rect 20220 30880 20226 30892
rect 22278 30880 22284 30892
rect 22336 30880 22342 30932
rect 23109 30923 23167 30929
rect 23109 30889 23121 30923
rect 23155 30920 23167 30923
rect 23290 30920 23296 30932
rect 23155 30892 23296 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 14550 30812 14556 30864
rect 14608 30852 14614 30864
rect 15286 30852 15292 30864
rect 14608 30824 15292 30852
rect 14608 30812 14614 30824
rect 15286 30812 15292 30824
rect 15344 30852 15350 30864
rect 15610 30855 15668 30861
rect 15610 30852 15622 30855
rect 15344 30824 15622 30852
rect 15344 30812 15350 30824
rect 15610 30821 15622 30824
rect 15656 30821 15668 30855
rect 18046 30852 18052 30864
rect 18007 30824 18052 30852
rect 15610 30815 15668 30821
rect 18046 30812 18052 30824
rect 18104 30812 18110 30864
rect 21085 30855 21143 30861
rect 21085 30821 21097 30855
rect 21131 30852 21143 30855
rect 21174 30852 21180 30864
rect 21131 30824 21180 30852
rect 21131 30821 21143 30824
rect 21085 30815 21143 30821
rect 21174 30812 21180 30824
rect 21232 30812 21238 30864
rect 12621 30787 12679 30793
rect 12621 30753 12633 30787
rect 12667 30784 12679 30787
rect 12710 30784 12716 30796
rect 12667 30756 12716 30784
rect 12667 30753 12679 30756
rect 12621 30747 12679 30753
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 13262 30744 13268 30796
rect 13320 30784 13326 30796
rect 13633 30787 13691 30793
rect 13633 30784 13645 30787
rect 13320 30756 13645 30784
rect 13320 30744 13326 30756
rect 13633 30753 13645 30756
rect 13679 30753 13691 30787
rect 13633 30747 13691 30753
rect 13906 30744 13912 30796
rect 13964 30784 13970 30796
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 13964 30756 14105 30784
rect 13964 30744 13970 30756
rect 14093 30753 14105 30756
rect 14139 30753 14151 30787
rect 14093 30747 14151 30753
rect 19848 30787 19906 30793
rect 19848 30753 19860 30787
rect 19894 30784 19906 30787
rect 20438 30784 20444 30796
rect 19894 30756 20444 30784
rect 19894 30753 19906 30756
rect 19848 30747 19906 30753
rect 20438 30744 20444 30756
rect 20496 30784 20502 30796
rect 20714 30784 20720 30796
rect 20496 30756 20720 30784
rect 20496 30744 20502 30756
rect 20714 30744 20720 30756
rect 20772 30744 20778 30796
rect 23216 30793 23244 30892
rect 23290 30880 23296 30892
rect 23348 30880 23354 30932
rect 23569 30923 23627 30929
rect 23569 30920 23581 30923
rect 23446 30892 23581 30920
rect 23201 30787 23259 30793
rect 23201 30753 23213 30787
rect 23247 30753 23259 30787
rect 23201 30747 23259 30753
rect 14369 30719 14427 30725
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 15289 30719 15347 30725
rect 15289 30716 15301 30719
rect 14415 30688 15301 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15289 30685 15301 30688
rect 15335 30716 15347 30719
rect 16574 30716 16580 30728
rect 15335 30688 16580 30716
rect 15335 30685 15347 30688
rect 15289 30679 15347 30685
rect 16574 30676 16580 30688
rect 16632 30676 16638 30728
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 19935 30719 19993 30725
rect 19935 30685 19947 30719
rect 19981 30716 19993 30719
rect 20346 30716 20352 30728
rect 19981 30688 20352 30716
rect 19981 30685 19993 30688
rect 19935 30679 19993 30685
rect 12759 30651 12817 30657
rect 12759 30617 12771 30651
rect 12805 30648 12817 30651
rect 17972 30648 18000 30679
rect 20346 30676 20352 30688
rect 20404 30716 20410 30728
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 20404 30688 21005 30716
rect 20404 30676 20410 30688
rect 20993 30685 21005 30688
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 21269 30719 21327 30725
rect 21269 30685 21281 30719
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 18414 30648 18420 30660
rect 12805 30620 18420 30648
rect 12805 30617 12817 30620
rect 12759 30611 12817 30617
rect 18414 30608 18420 30620
rect 18472 30608 18478 30660
rect 18509 30651 18567 30657
rect 18509 30617 18521 30651
rect 18555 30648 18567 30651
rect 21284 30648 21312 30679
rect 23106 30676 23112 30728
rect 23164 30716 23170 30728
rect 23446 30716 23474 30892
rect 23569 30889 23581 30892
rect 23615 30889 23627 30923
rect 24578 30920 24584 30932
rect 24539 30892 24584 30920
rect 23569 30883 23627 30889
rect 24578 30880 24584 30892
rect 24636 30920 24642 30932
rect 25087 30923 25145 30929
rect 25087 30920 25099 30923
rect 24636 30892 25099 30920
rect 24636 30880 24642 30892
rect 25087 30889 25099 30892
rect 25133 30889 25145 30923
rect 30006 30920 30012 30932
rect 29967 30892 30012 30920
rect 25087 30883 25145 30889
rect 30006 30880 30012 30892
rect 30064 30880 30070 30932
rect 31205 30923 31263 30929
rect 31205 30889 31217 30923
rect 31251 30920 31263 30923
rect 31386 30920 31392 30932
rect 31251 30892 31392 30920
rect 31251 30889 31263 30892
rect 31205 30883 31263 30889
rect 31386 30880 31392 30892
rect 31444 30880 31450 30932
rect 31662 30920 31668 30932
rect 31623 30892 31668 30920
rect 31662 30880 31668 30892
rect 31720 30880 31726 30932
rect 31754 30880 31760 30932
rect 31812 30920 31818 30932
rect 32398 30920 32404 30932
rect 31812 30892 32404 30920
rect 31812 30880 31818 30892
rect 32398 30880 32404 30892
rect 32456 30880 32462 30932
rect 34054 30920 34060 30932
rect 34015 30892 34060 30920
rect 34054 30880 34060 30892
rect 34112 30880 34118 30932
rect 34698 30920 34704 30932
rect 34624 30892 34704 30920
rect 26694 30852 26700 30864
rect 26655 30824 26700 30852
rect 26694 30812 26700 30824
rect 26752 30812 26758 30864
rect 26878 30812 26884 30864
rect 26936 30852 26942 30864
rect 27249 30855 27307 30861
rect 27249 30852 27261 30855
rect 26936 30824 27261 30852
rect 26936 30812 26942 30824
rect 27249 30821 27261 30824
rect 27295 30821 27307 30855
rect 29178 30852 29184 30864
rect 29139 30824 29184 30852
rect 27249 30815 27307 30821
rect 29178 30812 29184 30824
rect 29236 30812 29242 30864
rect 32122 30852 32128 30864
rect 32083 30824 32128 30852
rect 32122 30812 32128 30824
rect 32180 30812 32186 30864
rect 33689 30855 33747 30861
rect 33689 30821 33701 30855
rect 33735 30852 33747 30855
rect 34624 30852 34652 30892
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 35894 30920 35900 30932
rect 35855 30892 35900 30920
rect 35894 30880 35900 30892
rect 35952 30880 35958 30932
rect 39390 30880 39396 30932
rect 39448 30920 39454 30932
rect 40586 30920 40592 30932
rect 39448 30892 40592 30920
rect 39448 30880 39454 30892
rect 40586 30880 40592 30892
rect 40644 30880 40650 30932
rect 41138 30920 41144 30932
rect 41099 30892 41144 30920
rect 41138 30880 41144 30892
rect 41196 30880 41202 30932
rect 41598 30880 41604 30932
rect 41656 30920 41662 30932
rect 42337 30923 42395 30929
rect 42337 30920 42349 30923
rect 41656 30892 42349 30920
rect 41656 30880 41662 30892
rect 42337 30889 42349 30892
rect 42383 30889 42395 30923
rect 43070 30920 43076 30932
rect 43031 30892 43076 30920
rect 42337 30883 42395 30889
rect 43070 30880 43076 30892
rect 43128 30920 43134 30932
rect 43487 30923 43545 30929
rect 43487 30920 43499 30923
rect 43128 30892 43499 30920
rect 43128 30880 43134 30892
rect 43487 30889 43499 30892
rect 43533 30889 43545 30923
rect 43487 30883 43545 30889
rect 41506 30852 41512 30864
rect 33735 30824 34652 30852
rect 41467 30824 41512 30852
rect 33735 30821 33747 30824
rect 33689 30815 33747 30821
rect 41506 30812 41512 30824
rect 41564 30812 41570 30864
rect 44545 30855 44603 30861
rect 44545 30821 44557 30855
rect 44591 30852 44603 30855
rect 44634 30852 44640 30864
rect 44591 30824 44640 30852
rect 44591 30821 44603 30824
rect 44545 30815 44603 30821
rect 44634 30812 44640 30824
rect 44692 30812 44698 30864
rect 45094 30852 45100 30864
rect 45007 30824 45100 30852
rect 45094 30812 45100 30824
rect 45152 30852 45158 30864
rect 46842 30852 46848 30864
rect 45152 30824 46848 30852
rect 45152 30812 45158 30824
rect 46842 30812 46848 30824
rect 46900 30812 46906 30864
rect 24946 30784 24952 30796
rect 24907 30756 24952 30784
rect 24946 30744 24952 30756
rect 25004 30744 25010 30796
rect 31021 30787 31079 30793
rect 31021 30753 31033 30787
rect 31067 30784 31079 30787
rect 31110 30784 31116 30796
rect 31067 30756 31116 30784
rect 31067 30753 31079 30756
rect 31021 30747 31079 30753
rect 31110 30744 31116 30756
rect 31168 30744 31174 30796
rect 31846 30744 31852 30796
rect 31904 30784 31910 30796
rect 32272 30787 32330 30793
rect 32272 30784 32284 30787
rect 31904 30756 32284 30784
rect 31904 30744 31910 30756
rect 32272 30753 32284 30756
rect 32318 30753 32330 30787
rect 34514 30784 34520 30796
rect 34475 30756 34520 30784
rect 32272 30747 32330 30753
rect 34514 30744 34520 30756
rect 34572 30744 34578 30796
rect 34664 30787 34722 30793
rect 34664 30753 34676 30787
rect 34710 30784 34722 30787
rect 36081 30787 36139 30793
rect 36081 30784 36093 30787
rect 34710 30756 36093 30784
rect 34710 30753 34722 30756
rect 34664 30747 34722 30753
rect 36081 30753 36093 30756
rect 36127 30784 36139 30787
rect 36170 30784 36176 30796
rect 36127 30756 36176 30784
rect 36127 30753 36139 30756
rect 36081 30747 36139 30753
rect 36170 30744 36176 30756
rect 36228 30744 36234 30796
rect 36906 30744 36912 30796
rect 36964 30784 36970 30796
rect 37737 30787 37795 30793
rect 37737 30784 37749 30787
rect 36964 30756 37749 30784
rect 36964 30744 36970 30756
rect 37737 30753 37749 30756
rect 37783 30784 37795 30787
rect 38010 30784 38016 30796
rect 37783 30756 38016 30784
rect 37783 30753 37795 30756
rect 37737 30747 37795 30753
rect 38010 30744 38016 30756
rect 38068 30744 38074 30796
rect 38930 30744 38936 30796
rect 38988 30784 38994 30796
rect 39209 30787 39267 30793
rect 39209 30784 39221 30787
rect 38988 30756 39221 30784
rect 38988 30744 38994 30756
rect 39209 30753 39221 30756
rect 39255 30784 39267 30787
rect 39390 30784 39396 30796
rect 39255 30756 39396 30784
rect 39255 30753 39267 30756
rect 39209 30747 39267 30753
rect 39390 30744 39396 30756
rect 39448 30744 39454 30796
rect 39485 30787 39543 30793
rect 39485 30753 39497 30787
rect 39531 30784 39543 30787
rect 39574 30784 39580 30796
rect 39531 30756 39580 30784
rect 39531 30753 39543 30756
rect 39485 30747 39543 30753
rect 23164 30688 23474 30716
rect 26605 30719 26663 30725
rect 23164 30676 23170 30688
rect 26605 30685 26617 30719
rect 26651 30716 26663 30719
rect 27430 30716 27436 30728
rect 26651 30688 27436 30716
rect 26651 30685 26663 30688
rect 26605 30679 26663 30685
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 28905 30719 28963 30725
rect 28905 30685 28917 30719
rect 28951 30716 28963 30719
rect 29086 30716 29092 30728
rect 28951 30688 29092 30716
rect 28951 30685 28963 30688
rect 28905 30679 28963 30685
rect 29086 30676 29092 30688
rect 29144 30676 29150 30728
rect 30650 30676 30656 30728
rect 30708 30716 30714 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30708 30688 30941 30716
rect 30708 30676 30714 30688
rect 30929 30685 30941 30688
rect 30975 30716 30987 30719
rect 31754 30716 31760 30728
rect 30975 30688 31760 30716
rect 30975 30685 30987 30688
rect 30929 30679 30987 30685
rect 31754 30676 31760 30688
rect 31812 30676 31818 30728
rect 31938 30676 31944 30728
rect 31996 30716 32002 30728
rect 32493 30719 32551 30725
rect 32493 30716 32505 30719
rect 31996 30688 32505 30716
rect 31996 30676 32002 30688
rect 32493 30685 32505 30688
rect 32539 30716 32551 30719
rect 33226 30716 33232 30728
rect 32539 30688 33232 30716
rect 32539 30685 32551 30688
rect 32493 30679 32551 30685
rect 33226 30676 33232 30688
rect 33284 30676 33290 30728
rect 34882 30716 34888 30728
rect 34843 30688 34888 30716
rect 34882 30676 34888 30688
rect 34940 30676 34946 30728
rect 38838 30716 38844 30728
rect 37936 30688 38844 30716
rect 21358 30648 21364 30660
rect 18555 30620 21364 30648
rect 18555 30617 18567 30620
rect 18509 30611 18567 30617
rect 15470 30540 15476 30592
rect 15528 30580 15534 30592
rect 18524 30580 18552 30611
rect 21358 30608 21364 30620
rect 21416 30608 21422 30660
rect 29638 30648 29644 30660
rect 29599 30620 29644 30648
rect 29638 30608 29644 30620
rect 29696 30608 29702 30660
rect 29730 30608 29736 30660
rect 29788 30648 29794 30660
rect 32585 30651 32643 30657
rect 32585 30648 32597 30651
rect 29788 30620 32597 30648
rect 29788 30608 29794 30620
rect 32585 30617 32597 30620
rect 32631 30617 32643 30651
rect 32585 30611 32643 30617
rect 33134 30608 33140 30660
rect 33192 30648 33198 30660
rect 33192 30620 34376 30648
rect 33192 30608 33198 30620
rect 15528 30552 18552 30580
rect 15528 30540 15534 30552
rect 20254 30540 20260 30592
rect 20312 30580 20318 30592
rect 20349 30583 20407 30589
rect 20349 30580 20361 30583
rect 20312 30552 20361 30580
rect 20312 30540 20318 30552
rect 20349 30549 20361 30552
rect 20395 30549 20407 30583
rect 24118 30580 24124 30592
rect 24079 30552 24124 30580
rect 20349 30543 20407 30549
rect 24118 30540 24124 30552
rect 24176 30540 24182 30592
rect 26234 30580 26240 30592
rect 26195 30552 26240 30580
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 32401 30583 32459 30589
rect 32401 30549 32413 30583
rect 32447 30580 32459 30583
rect 32490 30580 32496 30592
rect 32447 30552 32496 30580
rect 32447 30549 32459 30552
rect 32401 30543 32459 30549
rect 32490 30540 32496 30552
rect 32548 30540 32554 30592
rect 33321 30583 33379 30589
rect 33321 30549 33333 30583
rect 33367 30580 33379 30583
rect 33410 30580 33416 30592
rect 33367 30552 33416 30580
rect 33367 30549 33379 30552
rect 33321 30543 33379 30549
rect 33410 30540 33416 30552
rect 33468 30540 33474 30592
rect 34348 30580 34376 30620
rect 34606 30608 34612 30660
rect 34664 30648 34670 30660
rect 34793 30651 34851 30657
rect 34793 30648 34805 30651
rect 34664 30620 34805 30648
rect 34664 30608 34670 30620
rect 34793 30617 34805 30620
rect 34839 30617 34851 30651
rect 34793 30611 34851 30617
rect 36909 30651 36967 30657
rect 36909 30617 36921 30651
rect 36955 30648 36967 30651
rect 37458 30648 37464 30660
rect 36955 30620 37464 30648
rect 36955 30617 36967 30620
rect 36909 30611 36967 30617
rect 37458 30608 37464 30620
rect 37516 30648 37522 30660
rect 37936 30657 37964 30688
rect 38838 30676 38844 30688
rect 38896 30716 38902 30728
rect 39500 30716 39528 30747
rect 39574 30744 39580 30756
rect 39632 30744 39638 30796
rect 43254 30744 43260 30796
rect 43312 30784 43318 30796
rect 43384 30787 43442 30793
rect 43384 30784 43396 30787
rect 43312 30756 43396 30784
rect 43312 30744 43318 30756
rect 43384 30753 43396 30756
rect 43430 30753 43442 30787
rect 45922 30784 45928 30796
rect 45883 30756 45928 30784
rect 43384 30747 43442 30753
rect 45922 30744 45928 30756
rect 45980 30744 45986 30796
rect 39666 30716 39672 30728
rect 38896 30688 39528 30716
rect 39627 30688 39672 30716
rect 38896 30676 38902 30688
rect 39666 30676 39672 30688
rect 39724 30676 39730 30728
rect 41417 30719 41475 30725
rect 41417 30685 41429 30719
rect 41463 30716 41475 30719
rect 41874 30716 41880 30728
rect 41463 30688 41880 30716
rect 41463 30685 41475 30688
rect 41417 30679 41475 30685
rect 41874 30676 41880 30688
rect 41932 30676 41938 30728
rect 42061 30719 42119 30725
rect 42061 30685 42073 30719
rect 42107 30716 42119 30719
rect 43070 30716 43076 30728
rect 42107 30688 43076 30716
rect 42107 30685 42119 30688
rect 42061 30679 42119 30685
rect 43070 30676 43076 30688
rect 43128 30676 43134 30728
rect 44453 30719 44511 30725
rect 44453 30685 44465 30719
rect 44499 30716 44511 30719
rect 45462 30716 45468 30728
rect 44499 30688 45468 30716
rect 44499 30685 44511 30688
rect 44453 30679 44511 30685
rect 45462 30676 45468 30688
rect 45520 30716 45526 30728
rect 46063 30719 46121 30725
rect 46063 30716 46075 30719
rect 45520 30688 46075 30716
rect 45520 30676 45526 30688
rect 46063 30685 46075 30688
rect 46109 30685 46121 30719
rect 46063 30679 46121 30685
rect 37921 30651 37979 30657
rect 37921 30648 37933 30651
rect 37516 30620 37933 30648
rect 37516 30608 37522 30620
rect 37921 30617 37933 30620
rect 37967 30617 37979 30651
rect 37921 30611 37979 30617
rect 34977 30583 35035 30589
rect 34977 30580 34989 30583
rect 34348 30552 34989 30580
rect 34977 30549 34989 30552
rect 35023 30549 35035 30583
rect 35618 30580 35624 30592
rect 35579 30552 35624 30580
rect 34977 30543 35035 30549
rect 35618 30540 35624 30552
rect 35676 30540 35682 30592
rect 36262 30580 36268 30592
rect 36223 30552 36268 30580
rect 36262 30540 36268 30552
rect 36320 30540 36326 30592
rect 38286 30540 38292 30592
rect 38344 30580 38350 30592
rect 38381 30583 38439 30589
rect 38381 30580 38393 30583
rect 38344 30552 38393 30580
rect 38344 30540 38350 30552
rect 38381 30549 38393 30552
rect 38427 30549 38439 30583
rect 40494 30580 40500 30592
rect 40455 30552 40500 30580
rect 38381 30543 38439 30549
rect 40494 30540 40500 30552
rect 40552 30540 40558 30592
rect 46753 30583 46811 30589
rect 46753 30549 46765 30583
rect 46799 30580 46811 30583
rect 47026 30580 47032 30592
rect 46799 30552 47032 30580
rect 46799 30549 46811 30552
rect 46753 30543 46811 30549
rect 47026 30540 47032 30552
rect 47084 30540 47090 30592
rect 1104 30490 48852 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 48852 30490
rect 1104 30416 48852 30438
rect 13262 30336 13268 30388
rect 13320 30376 13326 30388
rect 13357 30379 13415 30385
rect 13357 30376 13369 30379
rect 13320 30348 13369 30376
rect 13320 30336 13326 30348
rect 13357 30345 13369 30348
rect 13403 30376 13415 30379
rect 15102 30376 15108 30388
rect 13403 30348 15108 30376
rect 13403 30345 13415 30348
rect 13357 30339 13415 30345
rect 15102 30336 15108 30348
rect 15160 30336 15166 30388
rect 15286 30376 15292 30388
rect 15247 30348 15292 30376
rect 15286 30336 15292 30348
rect 15344 30336 15350 30388
rect 16574 30376 16580 30388
rect 16535 30348 16580 30376
rect 16574 30336 16580 30348
rect 16632 30336 16638 30388
rect 17497 30379 17555 30385
rect 17497 30345 17509 30379
rect 17543 30376 17555 30379
rect 18046 30376 18052 30388
rect 17543 30348 18052 30376
rect 17543 30345 17555 30348
rect 17497 30339 17555 30345
rect 18046 30336 18052 30348
rect 18104 30336 18110 30388
rect 18414 30336 18420 30388
rect 18472 30376 18478 30388
rect 19061 30379 19119 30385
rect 19061 30376 19073 30379
rect 18472 30348 19073 30376
rect 18472 30336 18478 30348
rect 19061 30345 19073 30348
rect 19107 30345 19119 30379
rect 20162 30376 20168 30388
rect 20123 30348 20168 30376
rect 19061 30339 19119 30345
rect 20162 30336 20168 30348
rect 20220 30336 20226 30388
rect 21174 30336 21180 30388
rect 21232 30376 21238 30388
rect 21637 30379 21695 30385
rect 21637 30376 21649 30379
rect 21232 30348 21649 30376
rect 21232 30336 21238 30348
rect 21637 30345 21649 30348
rect 21683 30345 21695 30379
rect 22370 30376 22376 30388
rect 22331 30348 22376 30376
rect 21637 30339 21695 30345
rect 22370 30336 22376 30348
rect 22428 30336 22434 30388
rect 23106 30336 23112 30388
rect 23164 30376 23170 30388
rect 23201 30379 23259 30385
rect 23201 30376 23213 30379
rect 23164 30348 23213 30376
rect 23164 30336 23170 30348
rect 23201 30345 23213 30348
rect 23247 30376 23259 30379
rect 23750 30376 23756 30388
rect 23247 30348 23756 30376
rect 23247 30345 23259 30348
rect 23201 30339 23259 30345
rect 23750 30336 23756 30348
rect 23808 30336 23814 30388
rect 24394 30336 24400 30388
rect 24452 30376 24458 30388
rect 24581 30379 24639 30385
rect 24581 30376 24593 30379
rect 24452 30348 24593 30376
rect 24452 30336 24458 30348
rect 24581 30345 24593 30348
rect 24627 30376 24639 30379
rect 25682 30376 25688 30388
rect 24627 30348 25688 30376
rect 24627 30345 24639 30348
rect 24581 30339 24639 30345
rect 25682 30336 25688 30348
rect 25740 30336 25746 30388
rect 27430 30376 27436 30388
rect 27391 30348 27436 30376
rect 27430 30336 27436 30348
rect 27488 30376 27494 30388
rect 28123 30379 28181 30385
rect 28123 30376 28135 30379
rect 27488 30348 28135 30376
rect 27488 30336 27494 30348
rect 28123 30345 28135 30348
rect 28169 30345 28181 30379
rect 28123 30339 28181 30345
rect 30653 30379 30711 30385
rect 30653 30345 30665 30379
rect 30699 30376 30711 30379
rect 31018 30376 31024 30388
rect 30699 30348 31024 30376
rect 30699 30345 30711 30348
rect 30653 30339 30711 30345
rect 31018 30336 31024 30348
rect 31076 30336 31082 30388
rect 31389 30379 31447 30385
rect 31389 30345 31401 30379
rect 31435 30376 31447 30379
rect 31757 30379 31815 30385
rect 31757 30376 31769 30379
rect 31435 30348 31769 30376
rect 31435 30345 31447 30348
rect 31389 30339 31447 30345
rect 31757 30345 31769 30348
rect 31803 30376 31815 30379
rect 32582 30376 32588 30388
rect 31803 30348 32588 30376
rect 31803 30345 31815 30348
rect 31757 30339 31815 30345
rect 32582 30336 32588 30348
rect 32640 30336 32646 30388
rect 33689 30379 33747 30385
rect 33689 30376 33701 30379
rect 32692 30348 33701 30376
rect 13679 30311 13737 30317
rect 13679 30277 13691 30311
rect 13725 30308 13737 30311
rect 20254 30308 20260 30320
rect 13725 30280 20260 30308
rect 13725 30277 13737 30280
rect 13679 30271 13737 30277
rect 20254 30268 20260 30280
rect 20312 30268 20318 30320
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 21266 30308 21272 30320
rect 20395 30280 21272 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 21266 30268 21272 30280
rect 21324 30268 21330 30320
rect 22830 30268 22836 30320
rect 22888 30308 22894 30320
rect 28626 30308 28632 30320
rect 22888 30280 28632 30308
rect 22888 30268 22894 30280
rect 28626 30268 28632 30280
rect 28684 30268 28690 30320
rect 31036 30308 31064 30336
rect 31619 30311 31677 30317
rect 31619 30308 31631 30311
rect 31036 30280 31631 30308
rect 31619 30277 31631 30280
rect 31665 30277 31677 30311
rect 31619 30271 31677 30277
rect 31938 30268 31944 30320
rect 31996 30308 32002 30320
rect 32692 30308 32720 30348
rect 33689 30345 33701 30348
rect 33735 30345 33747 30379
rect 33689 30339 33747 30345
rect 33778 30336 33784 30388
rect 33836 30376 33842 30388
rect 34517 30379 34575 30385
rect 34517 30376 34529 30379
rect 33836 30348 34529 30376
rect 33836 30336 33842 30348
rect 34517 30345 34529 30348
rect 34563 30376 34575 30379
rect 34790 30376 34796 30388
rect 34563 30348 34796 30376
rect 34563 30345 34575 30348
rect 34517 30339 34575 30345
rect 34790 30336 34796 30348
rect 34848 30336 34854 30388
rect 35069 30379 35127 30385
rect 35069 30345 35081 30379
rect 35115 30376 35127 30379
rect 35526 30376 35532 30388
rect 35115 30348 35532 30376
rect 35115 30345 35127 30348
rect 35069 30339 35127 30345
rect 35526 30336 35532 30348
rect 35584 30336 35590 30388
rect 35894 30336 35900 30388
rect 35952 30376 35958 30388
rect 36265 30379 36323 30385
rect 36265 30376 36277 30379
rect 35952 30348 36277 30376
rect 35952 30336 35958 30348
rect 36265 30345 36277 30348
rect 36311 30345 36323 30379
rect 37458 30376 37464 30388
rect 37419 30348 37464 30376
rect 36265 30339 36323 30345
rect 37458 30336 37464 30348
rect 37516 30336 37522 30388
rect 37734 30376 37740 30388
rect 37695 30348 37740 30376
rect 37734 30336 37740 30348
rect 37792 30336 37798 30388
rect 38010 30376 38016 30388
rect 37971 30348 38016 30376
rect 38010 30336 38016 30348
rect 38068 30336 38074 30388
rect 38470 30376 38476 30388
rect 38431 30348 38476 30376
rect 38470 30336 38476 30348
rect 38528 30336 38534 30388
rect 41874 30336 41880 30388
rect 41932 30376 41938 30388
rect 42061 30379 42119 30385
rect 42061 30376 42073 30379
rect 41932 30348 42073 30376
rect 41932 30336 41938 30348
rect 42061 30345 42073 30348
rect 42107 30345 42119 30379
rect 42061 30339 42119 30345
rect 43254 30336 43260 30388
rect 43312 30376 43318 30388
rect 43717 30379 43775 30385
rect 43717 30376 43729 30379
rect 43312 30348 43729 30376
rect 43312 30336 43318 30348
rect 43717 30345 43729 30348
rect 43763 30345 43775 30379
rect 43717 30339 43775 30345
rect 44358 30336 44364 30388
rect 44416 30376 44422 30388
rect 45094 30376 45100 30388
rect 44416 30348 45100 30376
rect 44416 30336 44422 30348
rect 45094 30336 45100 30348
rect 45152 30376 45158 30388
rect 45462 30376 45468 30388
rect 45152 30348 45324 30376
rect 45423 30348 45468 30376
rect 45152 30336 45158 30348
rect 31996 30280 32720 30308
rect 33137 30311 33195 30317
rect 31996 30268 32002 30280
rect 33137 30277 33149 30311
rect 33183 30308 33195 30311
rect 33505 30311 33563 30317
rect 33505 30308 33517 30311
rect 33183 30280 33517 30308
rect 33183 30277 33195 30280
rect 33137 30271 33195 30277
rect 33505 30277 33517 30280
rect 33551 30308 33563 30311
rect 34606 30308 34612 30320
rect 33551 30280 34612 30308
rect 33551 30277 33563 30280
rect 33505 30271 33563 30277
rect 34606 30268 34612 30280
rect 34664 30308 34670 30320
rect 35345 30311 35403 30317
rect 35345 30308 35357 30311
rect 34664 30280 35357 30308
rect 34664 30268 34670 30280
rect 35345 30277 35357 30280
rect 35391 30277 35403 30311
rect 35345 30271 35403 30277
rect 35713 30311 35771 30317
rect 35713 30277 35725 30311
rect 35759 30308 35771 30311
rect 36170 30308 36176 30320
rect 35759 30280 36176 30308
rect 35759 30277 35771 30280
rect 35713 30271 35771 30277
rect 14691 30243 14749 30249
rect 14691 30209 14703 30243
rect 14737 30240 14749 30243
rect 20717 30243 20775 30249
rect 20717 30240 20729 30243
rect 14737 30212 20729 30240
rect 14737 30209 14749 30212
rect 14691 30203 14749 30209
rect 20717 30209 20729 30212
rect 20763 30240 20775 30243
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 20763 30212 22017 30240
rect 20763 30209 20775 30212
rect 20717 30203 20775 30209
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 29273 30243 29331 30249
rect 29273 30209 29285 30243
rect 29319 30240 29331 30243
rect 29362 30240 29368 30252
rect 29319 30212 29368 30240
rect 29319 30209 29331 30212
rect 29273 30203 29331 30209
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 31846 30240 31852 30252
rect 31807 30212 31852 30240
rect 31846 30200 31852 30212
rect 31904 30200 31910 30252
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30240 33655 30243
rect 34054 30240 34060 30252
rect 33643 30212 34060 30240
rect 33643 30209 33655 30212
rect 33597 30203 33655 30209
rect 34054 30200 34060 30212
rect 34112 30200 34118 30252
rect 34514 30200 34520 30252
rect 34572 30240 34578 30252
rect 34701 30243 34759 30249
rect 34701 30240 34713 30243
rect 34572 30212 34713 30240
rect 34572 30200 34578 30212
rect 34701 30209 34713 30212
rect 34747 30209 34759 30243
rect 35728 30240 35756 30271
rect 36170 30268 36176 30280
rect 36228 30268 36234 30320
rect 45296 30308 45324 30348
rect 45462 30336 45468 30348
rect 45520 30336 45526 30388
rect 47578 30376 47584 30388
rect 47539 30348 47584 30376
rect 47578 30336 47584 30348
rect 47636 30336 47642 30388
rect 45922 30308 45928 30320
rect 42812 30280 45048 30308
rect 45296 30280 45928 30308
rect 42812 30252 42840 30280
rect 45020 30252 45048 30280
rect 45922 30268 45928 30280
rect 45980 30308 45986 30320
rect 46293 30311 46351 30317
rect 46293 30308 46305 30311
rect 45980 30280 46305 30308
rect 45980 30268 45986 30280
rect 46293 30277 46305 30280
rect 46339 30277 46351 30311
rect 46293 30271 46351 30277
rect 34701 30203 34759 30209
rect 34808 30212 35756 30240
rect 13608 30175 13666 30181
rect 13608 30141 13620 30175
rect 13654 30172 13666 30175
rect 14588 30175 14646 30181
rect 13654 30144 13814 30172
rect 13654 30141 13666 30144
rect 13608 30135 13666 30141
rect 12710 30036 12716 30048
rect 12671 30008 12716 30036
rect 12710 29996 12716 30008
rect 12768 29996 12774 30048
rect 13078 30036 13084 30048
rect 13039 30008 13084 30036
rect 13078 29996 13084 30008
rect 13136 29996 13142 30048
rect 13786 30036 13814 30144
rect 14588 30141 14600 30175
rect 14634 30141 14646 30175
rect 14588 30135 14646 30141
rect 19680 30175 19738 30181
rect 19680 30141 19692 30175
rect 19726 30172 19738 30175
rect 20162 30172 20168 30184
rect 19726 30144 20168 30172
rect 19726 30141 19738 30144
rect 19680 30135 19738 30141
rect 14090 30036 14096 30048
rect 13786 30008 14096 30036
rect 14090 29996 14096 30008
rect 14148 29996 14154 30048
rect 14461 30039 14519 30045
rect 14461 30005 14473 30039
rect 14507 30036 14519 30039
rect 14603 30036 14631 30135
rect 20162 30132 20168 30144
rect 20220 30172 20226 30184
rect 22189 30175 22247 30181
rect 20220 30144 20576 30172
rect 20220 30132 20226 30144
rect 15470 30064 15476 30116
rect 15528 30104 15534 30116
rect 15657 30107 15715 30113
rect 15657 30104 15669 30107
rect 15528 30076 15669 30104
rect 15528 30064 15534 30076
rect 15657 30073 15669 30076
rect 15703 30073 15715 30107
rect 15657 30067 15715 30073
rect 15746 30064 15752 30116
rect 15804 30104 15810 30116
rect 16301 30107 16359 30113
rect 15804 30076 15849 30104
rect 15804 30064 15810 30076
rect 16301 30073 16313 30107
rect 16347 30104 16359 30107
rect 16482 30104 16488 30116
rect 16347 30076 16488 30104
rect 16347 30073 16359 30076
rect 16301 30067 16359 30073
rect 16482 30064 16488 30076
rect 16540 30064 16546 30116
rect 18141 30107 18199 30113
rect 18141 30073 18153 30107
rect 18187 30073 18199 30107
rect 18141 30067 18199 30073
rect 16574 30036 16580 30048
rect 14507 30008 16580 30036
rect 14507 30005 14519 30008
rect 14461 29999 14519 30005
rect 16574 29996 16580 30008
rect 16632 29996 16638 30048
rect 16942 30036 16948 30048
rect 16903 30008 16948 30036
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 17770 30036 17776 30048
rect 17731 30008 17776 30036
rect 17770 29996 17776 30008
rect 17828 30036 17834 30048
rect 18156 30036 18184 30067
rect 18230 30064 18236 30116
rect 18288 30104 18294 30116
rect 18782 30104 18788 30116
rect 18288 30076 18333 30104
rect 18695 30076 18788 30104
rect 18288 30064 18294 30076
rect 18782 30064 18788 30076
rect 18840 30104 18846 30116
rect 20349 30107 20407 30113
rect 20349 30104 20361 30107
rect 18840 30076 20361 30104
rect 18840 30064 18846 30076
rect 20349 30073 20361 30076
rect 20395 30073 20407 30107
rect 20548 30104 20576 30144
rect 22189 30141 22201 30175
rect 22235 30172 22247 30175
rect 22738 30172 22744 30184
rect 22235 30144 22744 30172
rect 22235 30141 22247 30144
rect 22189 30135 22247 30141
rect 22738 30132 22744 30144
rect 22796 30132 22802 30184
rect 23658 30172 23664 30184
rect 23619 30144 23664 30172
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 26237 30175 26295 30181
rect 26237 30141 26249 30175
rect 26283 30172 26295 30175
rect 26326 30172 26332 30184
rect 26283 30144 26332 30172
rect 26283 30141 26295 30144
rect 26237 30135 26295 30141
rect 26326 30132 26332 30144
rect 26384 30132 26390 30184
rect 28052 30175 28110 30181
rect 28052 30141 28064 30175
rect 28098 30141 28110 30175
rect 28052 30135 28110 30141
rect 20714 30104 20720 30116
rect 20548 30076 20720 30104
rect 20349 30067 20407 30073
rect 20714 30064 20720 30076
rect 20772 30064 20778 30116
rect 20809 30107 20867 30113
rect 20809 30073 20821 30107
rect 20855 30104 20867 30107
rect 21082 30104 21088 30116
rect 20855 30076 21088 30104
rect 20855 30073 20867 30076
rect 20809 30067 20867 30073
rect 21082 30064 21088 30076
rect 21140 30064 21146 30116
rect 23750 30064 23756 30116
rect 23808 30104 23814 30116
rect 24023 30107 24081 30113
rect 24023 30104 24035 30107
rect 23808 30076 24035 30104
rect 23808 30064 23814 30076
rect 24023 30073 24035 30076
rect 24069 30104 24081 30107
rect 26142 30104 26148 30116
rect 24069 30076 26148 30104
rect 24069 30073 24081 30076
rect 24023 30067 24081 30073
rect 26142 30064 26148 30076
rect 26200 30104 26206 30116
rect 26599 30107 26657 30113
rect 26599 30104 26611 30107
rect 26200 30076 26611 30104
rect 26200 30064 26206 30076
rect 26599 30073 26611 30076
rect 26645 30104 26657 30107
rect 28067 30104 28095 30135
rect 29178 30132 29184 30184
rect 29236 30172 29242 30184
rect 30193 30175 30251 30181
rect 30193 30172 30205 30175
rect 29236 30144 30205 30172
rect 29236 30132 29242 30144
rect 30193 30141 30205 30144
rect 30239 30141 30251 30175
rect 30193 30135 30251 30141
rect 31021 30175 31079 30181
rect 31021 30141 31033 30175
rect 31067 30172 31079 30175
rect 31110 30172 31116 30184
rect 31067 30144 31116 30172
rect 31067 30141 31079 30144
rect 31021 30135 31079 30141
rect 31110 30132 31116 30144
rect 31168 30172 31174 30184
rect 32490 30172 32496 30184
rect 31168 30144 32496 30172
rect 31168 30132 31174 30144
rect 32490 30132 32496 30144
rect 32548 30132 32554 30184
rect 33410 30181 33416 30184
rect 33376 30175 33416 30181
rect 33376 30172 33388 30175
rect 33323 30144 33388 30172
rect 33376 30141 33388 30144
rect 33468 30172 33474 30184
rect 34808 30172 34836 30212
rect 36354 30200 36360 30252
rect 36412 30240 36418 30252
rect 36412 30212 36457 30240
rect 36412 30200 36418 30212
rect 39298 30200 39304 30252
rect 39356 30240 39362 30252
rect 41506 30240 41512 30252
rect 39356 30212 41512 30240
rect 39356 30200 39362 30212
rect 41506 30200 41512 30212
rect 41564 30240 41570 30252
rect 41693 30243 41751 30249
rect 41693 30240 41705 30243
rect 41564 30212 41705 30240
rect 41564 30200 41570 30212
rect 41693 30209 41705 30212
rect 41739 30209 41751 30243
rect 41693 30203 41751 30209
rect 42794 30200 42800 30252
rect 42852 30240 42858 30252
rect 43070 30240 43076 30252
rect 42852 30212 42945 30240
rect 43031 30212 43076 30240
rect 42852 30200 42858 30212
rect 43070 30200 43076 30212
rect 43128 30200 43134 30252
rect 45002 30240 45008 30252
rect 44963 30212 45008 30240
rect 45002 30200 45008 30212
rect 45060 30200 45066 30252
rect 46934 30240 46940 30252
rect 46676 30212 46940 30240
rect 33468 30144 34836 30172
rect 36136 30175 36194 30181
rect 33376 30135 33416 30141
rect 33410 30132 33416 30135
rect 33468 30132 33474 30144
rect 36136 30141 36148 30175
rect 36182 30172 36194 30175
rect 36262 30172 36268 30184
rect 36182 30144 36268 30172
rect 36182 30141 36194 30144
rect 36136 30135 36194 30141
rect 36262 30132 36268 30144
rect 36320 30132 36326 30184
rect 37550 30172 37556 30184
rect 37511 30144 37556 30172
rect 37550 30132 37556 30144
rect 37608 30132 37614 30184
rect 38470 30132 38476 30184
rect 38528 30172 38534 30184
rect 38565 30175 38623 30181
rect 38565 30172 38577 30175
rect 38528 30144 38577 30172
rect 38528 30132 38534 30144
rect 38565 30141 38577 30144
rect 38611 30141 38623 30175
rect 38565 30135 38623 30141
rect 39117 30175 39175 30181
rect 39117 30141 39129 30175
rect 39163 30172 39175 30175
rect 39574 30172 39580 30184
rect 39163 30144 39580 30172
rect 39163 30141 39175 30144
rect 39117 30135 39175 30141
rect 39574 30132 39580 30144
rect 39632 30132 39638 30184
rect 39758 30132 39764 30184
rect 39816 30172 39822 30184
rect 40494 30172 40500 30184
rect 39816 30144 40500 30172
rect 39816 30132 39822 30144
rect 40494 30132 40500 30144
rect 40552 30132 40558 30184
rect 46676 30181 46704 30212
rect 46934 30200 46940 30212
rect 46992 30240 46998 30252
rect 47596 30240 47624 30336
rect 46992 30212 47624 30240
rect 46992 30200 46998 30212
rect 46661 30175 46719 30181
rect 46661 30141 46673 30175
rect 46707 30141 46719 30175
rect 46661 30135 46719 30141
rect 46845 30175 46903 30181
rect 46845 30141 46857 30175
rect 46891 30172 46903 30175
rect 47026 30172 47032 30184
rect 46891 30144 47032 30172
rect 46891 30141 46903 30144
rect 46845 30135 46903 30141
rect 47026 30132 47032 30144
rect 47084 30132 47090 30184
rect 28537 30107 28595 30113
rect 28537 30104 28549 30107
rect 26645 30076 27936 30104
rect 28067 30076 28549 30104
rect 26645 30073 26657 30076
rect 26599 30067 26657 30073
rect 17828 30008 18184 30036
rect 19751 30039 19809 30045
rect 17828 29996 17834 30008
rect 19751 30005 19763 30039
rect 19797 30036 19809 30039
rect 19978 30036 19984 30048
rect 19797 30008 19984 30036
rect 19797 30005 19809 30008
rect 19751 29999 19809 30005
rect 19978 29996 19984 30008
rect 20036 29996 20042 30048
rect 20438 30036 20444 30048
rect 20399 30008 20444 30036
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 24946 30036 24952 30048
rect 24907 30008 24952 30036
rect 24946 29996 24952 30008
rect 25004 29996 25010 30048
rect 27154 30036 27160 30048
rect 27115 30008 27160 30036
rect 27154 29996 27160 30008
rect 27212 29996 27218 30048
rect 27908 30036 27936 30076
rect 28537 30073 28549 30076
rect 28583 30104 28595 30107
rect 29086 30104 29092 30116
rect 28583 30076 29092 30104
rect 28583 30073 28595 30076
rect 28537 30067 28595 30073
rect 29086 30064 29092 30076
rect 29144 30064 29150 30116
rect 29594 30107 29652 30113
rect 29594 30073 29606 30107
rect 29640 30073 29652 30107
rect 29594 30067 29652 30073
rect 31481 30107 31539 30113
rect 31481 30073 31493 30107
rect 31527 30104 31539 30107
rect 31662 30104 31668 30116
rect 31527 30076 31668 30104
rect 31527 30073 31539 30076
rect 31481 30067 31539 30073
rect 28718 30036 28724 30048
rect 27908 30008 28724 30036
rect 28718 29996 28724 30008
rect 28776 30036 28782 30048
rect 28997 30039 29055 30045
rect 28997 30036 29009 30039
rect 28776 30008 29009 30036
rect 28776 29996 28782 30008
rect 28997 30005 29009 30008
rect 29043 30036 29055 30039
rect 29609 30036 29637 30067
rect 31662 30064 31668 30076
rect 31720 30064 31726 30116
rect 32950 30064 32956 30116
rect 33008 30104 33014 30116
rect 33229 30107 33287 30113
rect 33229 30104 33241 30107
rect 33008 30076 33241 30104
rect 33008 30064 33014 30076
rect 33229 30073 33241 30076
rect 33275 30104 33287 30107
rect 34698 30104 34704 30116
rect 33275 30076 34704 30104
rect 33275 30073 33287 30076
rect 33229 30067 33287 30073
rect 34698 30064 34704 30076
rect 34756 30064 34762 30116
rect 35618 30064 35624 30116
rect 35676 30104 35682 30116
rect 35989 30107 36047 30113
rect 35989 30104 36001 30107
rect 35676 30076 36001 30104
rect 35676 30064 35682 30076
rect 35989 30073 36001 30076
rect 36035 30104 36047 30107
rect 36035 30076 37136 30104
rect 36035 30073 36047 30076
rect 35989 30067 36047 30073
rect 37108 30048 37136 30076
rect 37274 30064 37280 30116
rect 37332 30104 37338 30116
rect 38488 30104 38516 30132
rect 37332 30076 38516 30104
rect 39301 30107 39359 30113
rect 37332 30064 37338 30076
rect 39301 30073 39313 30107
rect 39347 30104 39359 30107
rect 40678 30104 40684 30116
rect 39347 30076 40684 30104
rect 39347 30073 39359 30076
rect 39301 30067 39359 30073
rect 40678 30064 40684 30076
rect 40736 30064 40742 30116
rect 40818 30107 40876 30113
rect 40818 30073 40830 30107
rect 40864 30073 40876 30107
rect 40818 30067 40876 30073
rect 42889 30107 42947 30113
rect 42889 30073 42901 30107
rect 42935 30073 42947 30107
rect 42889 30067 42947 30073
rect 44361 30107 44419 30113
rect 44361 30073 44373 30107
rect 44407 30104 44419 30107
rect 44542 30104 44548 30116
rect 44407 30076 44548 30104
rect 44407 30073 44419 30076
rect 44361 30067 44419 30073
rect 29043 30008 29637 30036
rect 29043 30005 29055 30008
rect 28997 29999 29055 30005
rect 31386 29996 31392 30048
rect 31444 30036 31450 30048
rect 32125 30039 32183 30045
rect 32125 30036 32137 30039
rect 31444 30008 32137 30036
rect 31444 29996 31450 30008
rect 32125 30005 32137 30008
rect 32171 30005 32183 30039
rect 32582 30036 32588 30048
rect 32543 30008 32588 30036
rect 32125 29999 32183 30005
rect 32582 29996 32588 30008
rect 32640 29996 32646 30048
rect 35802 29996 35808 30048
rect 35860 30036 35866 30048
rect 36633 30039 36691 30045
rect 36633 30036 36645 30039
rect 35860 30008 36645 30036
rect 35860 29996 35866 30008
rect 36633 30005 36645 30008
rect 36679 30005 36691 30039
rect 37090 30036 37096 30048
rect 37051 30008 37096 30036
rect 36633 29999 36691 30005
rect 37090 29996 37096 30008
rect 37148 29996 37154 30048
rect 39482 29996 39488 30048
rect 39540 30036 39546 30048
rect 39577 30039 39635 30045
rect 39577 30036 39589 30039
rect 39540 30008 39589 30036
rect 39540 29996 39546 30008
rect 39577 30005 39589 30008
rect 39623 30005 39635 30039
rect 40218 30036 40224 30048
rect 40179 30008 40224 30036
rect 39577 29999 39635 30005
rect 40218 29996 40224 30008
rect 40276 30036 40282 30048
rect 40833 30036 40861 30067
rect 41414 30036 41420 30048
rect 40276 30008 40861 30036
rect 41375 30008 41420 30036
rect 40276 29996 40282 30008
rect 41414 29996 41420 30008
rect 41472 29996 41478 30048
rect 42426 29996 42432 30048
rect 42484 30036 42490 30048
rect 42613 30039 42671 30045
rect 42613 30036 42625 30039
rect 42484 30008 42625 30036
rect 42484 29996 42490 30008
rect 42613 30005 42625 30008
rect 42659 30036 42671 30039
rect 42904 30036 42932 30067
rect 44542 30064 44548 30076
rect 44600 30064 44606 30116
rect 44634 30064 44640 30116
rect 44692 30104 44698 30116
rect 44692 30076 44737 30104
rect 44692 30064 44698 30076
rect 42659 30008 42932 30036
rect 42659 30005 42671 30008
rect 42613 29999 42671 30005
rect 46382 29996 46388 30048
rect 46440 30036 46446 30048
rect 46937 30039 46995 30045
rect 46937 30036 46949 30039
rect 46440 30008 46949 30036
rect 46440 29996 46446 30008
rect 46937 30005 46949 30008
rect 46983 30005 46995 30039
rect 46937 29999 46995 30005
rect 1104 29946 48852 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 48852 29946
rect 1104 29872 48852 29894
rect 14366 29792 14372 29844
rect 14424 29832 14430 29844
rect 15013 29835 15071 29841
rect 15013 29832 15025 29835
rect 14424 29804 15025 29832
rect 14424 29792 14430 29804
rect 15013 29801 15025 29804
rect 15059 29832 15071 29835
rect 15470 29832 15476 29844
rect 15059 29804 15476 29832
rect 15059 29801 15071 29804
rect 15013 29795 15071 29801
rect 15470 29792 15476 29804
rect 15528 29792 15534 29844
rect 15746 29792 15752 29844
rect 15804 29832 15810 29844
rect 16209 29835 16267 29841
rect 16209 29832 16221 29835
rect 15804 29804 16221 29832
rect 15804 29792 15810 29804
rect 16209 29801 16221 29804
rect 16255 29832 16267 29835
rect 16942 29832 16948 29844
rect 16255 29804 16948 29832
rect 16255 29801 16267 29804
rect 16209 29795 16267 29801
rect 16942 29792 16948 29804
rect 17000 29792 17006 29844
rect 17221 29835 17279 29841
rect 17221 29801 17233 29835
rect 17267 29832 17279 29835
rect 17770 29832 17776 29844
rect 17267 29804 17776 29832
rect 17267 29801 17279 29804
rect 17221 29795 17279 29801
rect 17770 29792 17776 29804
rect 17828 29792 17834 29844
rect 18046 29832 18052 29844
rect 18007 29804 18052 29832
rect 18046 29792 18052 29804
rect 18104 29792 18110 29844
rect 20346 29832 20352 29844
rect 20307 29804 20352 29832
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 23750 29832 23756 29844
rect 23711 29804 23756 29832
rect 23750 29792 23756 29804
rect 23808 29792 23814 29844
rect 28718 29792 28724 29844
rect 28776 29832 28782 29844
rect 28813 29835 28871 29841
rect 28813 29832 28825 29835
rect 28776 29804 28825 29832
rect 28776 29792 28782 29804
rect 28813 29801 28825 29804
rect 28859 29801 28871 29835
rect 28813 29795 28871 29801
rect 29362 29792 29368 29844
rect 29420 29832 29426 29844
rect 30009 29835 30067 29841
rect 30009 29832 30021 29835
rect 29420 29804 30021 29832
rect 29420 29792 29426 29804
rect 30009 29801 30021 29804
rect 30055 29801 30067 29835
rect 30009 29795 30067 29801
rect 30466 29792 30472 29844
rect 30524 29832 30530 29844
rect 30837 29835 30895 29841
rect 30837 29832 30849 29835
rect 30524 29804 30849 29832
rect 30524 29792 30530 29804
rect 30837 29801 30849 29804
rect 30883 29801 30895 29835
rect 30837 29795 30895 29801
rect 31205 29835 31263 29841
rect 31205 29801 31217 29835
rect 31251 29832 31263 29835
rect 31478 29832 31484 29844
rect 31251 29804 31484 29832
rect 31251 29801 31263 29804
rect 31205 29795 31263 29801
rect 31478 29792 31484 29804
rect 31536 29792 31542 29844
rect 31573 29835 31631 29841
rect 31573 29801 31585 29835
rect 31619 29832 31631 29835
rect 31662 29832 31668 29844
rect 31619 29804 31668 29832
rect 31619 29801 31631 29804
rect 31573 29795 31631 29801
rect 31662 29792 31668 29804
rect 31720 29792 31726 29844
rect 32122 29792 32128 29844
rect 32180 29832 32186 29844
rect 32309 29835 32367 29841
rect 32309 29832 32321 29835
rect 32180 29804 32321 29832
rect 32180 29792 32186 29804
rect 32309 29801 32321 29804
rect 32355 29801 32367 29835
rect 32309 29795 32367 29801
rect 33226 29792 33232 29844
rect 33284 29832 33290 29844
rect 34514 29832 34520 29844
rect 33284 29804 34520 29832
rect 33284 29792 33290 29804
rect 34514 29792 34520 29804
rect 34572 29832 34578 29844
rect 35618 29832 35624 29844
rect 34572 29804 35624 29832
rect 34572 29792 34578 29804
rect 35618 29792 35624 29804
rect 35676 29792 35682 29844
rect 35805 29835 35863 29841
rect 35805 29801 35817 29835
rect 35851 29832 35863 29835
rect 35894 29832 35900 29844
rect 35851 29804 35900 29832
rect 35851 29801 35863 29804
rect 35805 29795 35863 29801
rect 35894 29792 35900 29804
rect 35952 29792 35958 29844
rect 36170 29832 36176 29844
rect 36131 29804 36176 29832
rect 36170 29792 36176 29804
rect 36228 29792 36234 29844
rect 36262 29792 36268 29844
rect 36320 29832 36326 29844
rect 36449 29835 36507 29841
rect 36449 29832 36461 29835
rect 36320 29804 36461 29832
rect 36320 29792 36326 29804
rect 36449 29801 36461 29804
rect 36495 29801 36507 29835
rect 36449 29795 36507 29801
rect 36817 29835 36875 29841
rect 36817 29801 36829 29835
rect 36863 29832 36875 29835
rect 36998 29832 37004 29844
rect 36863 29804 37004 29832
rect 36863 29801 36875 29804
rect 36817 29795 36875 29801
rect 36998 29792 37004 29804
rect 37056 29792 37062 29844
rect 38654 29792 38660 29844
rect 38712 29832 38718 29844
rect 38749 29835 38807 29841
rect 38749 29832 38761 29835
rect 38712 29804 38761 29832
rect 38712 29792 38718 29804
rect 38749 29801 38761 29804
rect 38795 29801 38807 29835
rect 39298 29832 39304 29844
rect 39259 29804 39304 29832
rect 38749 29795 38807 29801
rect 39298 29792 39304 29804
rect 39356 29792 39362 29844
rect 39666 29792 39672 29844
rect 39724 29832 39730 29844
rect 40494 29832 40500 29844
rect 39724 29804 40500 29832
rect 39724 29792 39730 29804
rect 40494 29792 40500 29804
rect 40552 29832 40558 29844
rect 40589 29835 40647 29841
rect 40589 29832 40601 29835
rect 40552 29804 40601 29832
rect 40552 29792 40558 29804
rect 40589 29801 40601 29804
rect 40635 29801 40647 29835
rect 42426 29832 42432 29844
rect 42387 29804 42432 29832
rect 40589 29795 40647 29801
rect 42426 29792 42432 29804
rect 42484 29792 42490 29844
rect 43717 29835 43775 29841
rect 43717 29832 43729 29835
rect 42766 29804 43729 29832
rect 14550 29764 14556 29776
rect 13832 29736 14556 29764
rect 13832 29705 13860 29736
rect 14550 29724 14556 29736
rect 14608 29724 14614 29776
rect 15286 29724 15292 29776
rect 15344 29764 15350 29776
rect 15610 29767 15668 29773
rect 15610 29764 15622 29767
rect 15344 29736 15622 29764
rect 15344 29724 15350 29736
rect 15610 29733 15622 29736
rect 15656 29733 15668 29767
rect 18414 29764 18420 29776
rect 18375 29736 18420 29764
rect 15610 29727 15668 29733
rect 18414 29724 18420 29736
rect 18472 29724 18478 29776
rect 20717 29767 20775 29773
rect 20717 29733 20729 29767
rect 20763 29764 20775 29767
rect 21082 29764 21088 29776
rect 20763 29736 21088 29764
rect 20763 29733 20775 29736
rect 20717 29727 20775 29733
rect 21082 29724 21088 29736
rect 21140 29724 21146 29776
rect 23385 29767 23443 29773
rect 23385 29733 23397 29767
rect 23431 29764 23443 29767
rect 23658 29764 23664 29776
rect 23431 29736 23664 29764
rect 23431 29733 23443 29736
rect 23385 29727 23443 29733
rect 23658 29724 23664 29736
rect 23716 29764 23722 29776
rect 24029 29767 24087 29773
rect 24029 29764 24041 29767
rect 23716 29736 24041 29764
rect 23716 29724 23722 29736
rect 24029 29733 24041 29736
rect 24075 29733 24087 29767
rect 24029 29727 24087 29733
rect 24118 29724 24124 29776
rect 24176 29764 24182 29776
rect 24397 29767 24455 29773
rect 24397 29764 24409 29767
rect 24176 29736 24409 29764
rect 24176 29724 24182 29736
rect 24397 29733 24409 29736
rect 24443 29733 24455 29767
rect 24397 29727 24455 29733
rect 26881 29767 26939 29773
rect 26881 29733 26893 29767
rect 26927 29764 26939 29767
rect 27154 29764 27160 29776
rect 26927 29736 27160 29764
rect 26927 29733 26939 29736
rect 26881 29727 26939 29733
rect 27154 29724 27160 29736
rect 27212 29724 27218 29776
rect 29178 29724 29184 29776
rect 29236 29764 29242 29776
rect 29641 29767 29699 29773
rect 29641 29764 29653 29767
rect 29236 29736 29653 29764
rect 29236 29724 29242 29736
rect 29641 29733 29653 29736
rect 29687 29733 29699 29767
rect 29641 29727 29699 29733
rect 30561 29767 30619 29773
rect 30561 29733 30573 29767
rect 30607 29764 30619 29767
rect 31846 29764 31852 29776
rect 30607 29736 31852 29764
rect 30607 29733 30619 29736
rect 30561 29727 30619 29733
rect 31846 29724 31852 29736
rect 31904 29724 31910 29776
rect 34149 29767 34207 29773
rect 34149 29733 34161 29767
rect 34195 29764 34207 29767
rect 34330 29764 34336 29776
rect 34195 29736 34336 29764
rect 34195 29733 34207 29736
rect 34149 29727 34207 29733
rect 34330 29724 34336 29736
rect 34388 29764 34394 29776
rect 35912 29764 35940 29792
rect 37461 29767 37519 29773
rect 37461 29764 37473 29767
rect 34388 29736 35480 29764
rect 35912 29736 37473 29764
rect 34388 29724 34394 29736
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29665 13875 29699
rect 13817 29659 13875 29665
rect 13906 29656 13912 29708
rect 13964 29696 13970 29708
rect 14093 29699 14151 29705
rect 14093 29696 14105 29699
rect 13964 29668 14105 29696
rect 13964 29656 13970 29668
rect 14093 29665 14105 29668
rect 14139 29665 14151 29699
rect 14093 29659 14151 29665
rect 19797 29699 19855 29705
rect 19797 29665 19809 29699
rect 19843 29696 19855 29699
rect 19886 29696 19892 29708
rect 19843 29668 19892 29696
rect 19843 29665 19855 29668
rect 19797 29659 19855 29665
rect 19886 29656 19892 29668
rect 19944 29696 19950 29708
rect 20806 29696 20812 29708
rect 19944 29668 20812 29696
rect 19944 29656 19950 29668
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 22922 29696 22928 29708
rect 22883 29668 22928 29696
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23198 29696 23204 29708
rect 23159 29668 23204 29696
rect 23198 29656 23204 29668
rect 23256 29656 23262 29708
rect 31018 29696 31024 29708
rect 30979 29668 31024 29696
rect 31018 29656 31024 29668
rect 31076 29656 31082 29708
rect 31941 29699 31999 29705
rect 31941 29665 31953 29699
rect 31987 29696 31999 29699
rect 33192 29699 33250 29705
rect 31987 29668 33134 29696
rect 31987 29665 31999 29668
rect 31941 29659 31999 29665
rect 13722 29588 13728 29640
rect 13780 29628 13786 29640
rect 14366 29628 14372 29640
rect 13780 29600 14372 29628
rect 13780 29588 13786 29600
rect 14366 29588 14372 29600
rect 14424 29588 14430 29640
rect 15286 29628 15292 29640
rect 15247 29600 15292 29628
rect 15286 29588 15292 29600
rect 15344 29588 15350 29640
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29628 18383 29631
rect 18782 29628 18788 29640
rect 18371 29600 18788 29628
rect 18371 29597 18383 29600
rect 18325 29591 18383 29597
rect 18782 29588 18788 29600
rect 18840 29588 18846 29640
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20036 29600 21005 29628
rect 20036 29588 20042 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21269 29631 21327 29637
rect 21269 29597 21281 29631
rect 21315 29597 21327 29631
rect 21269 29591 21327 29597
rect 24305 29631 24363 29637
rect 24305 29597 24317 29631
rect 24351 29628 24363 29631
rect 24762 29628 24768 29640
rect 24351 29600 24768 29628
rect 24351 29597 24363 29600
rect 24305 29591 24363 29597
rect 16482 29520 16488 29572
rect 16540 29560 16546 29572
rect 18877 29563 18935 29569
rect 18877 29560 18889 29563
rect 16540 29532 18889 29560
rect 16540 29520 16546 29532
rect 18877 29529 18889 29532
rect 18923 29529 18935 29563
rect 18877 29523 18935 29529
rect 18966 29520 18972 29572
rect 19024 29560 19030 29572
rect 21284 29560 21312 29591
rect 24762 29588 24768 29600
rect 24820 29588 24826 29640
rect 26789 29631 26847 29637
rect 26789 29597 26801 29631
rect 26835 29628 26847 29631
rect 26878 29628 26884 29640
rect 26835 29600 26884 29628
rect 26835 29597 26847 29600
rect 26789 29591 26847 29597
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 28258 29588 28264 29640
rect 28316 29628 28322 29640
rect 28445 29631 28503 29637
rect 28445 29628 28457 29631
rect 28316 29600 28457 29628
rect 28316 29588 28322 29600
rect 28445 29597 28457 29600
rect 28491 29597 28503 29631
rect 33106 29628 33134 29668
rect 33192 29665 33204 29699
rect 33238 29696 33250 29699
rect 33686 29696 33692 29708
rect 33238 29668 33692 29696
rect 33238 29665 33250 29668
rect 33192 29659 33250 29665
rect 33686 29656 33692 29668
rect 33744 29656 33750 29708
rect 34609 29699 34667 29705
rect 34609 29665 34621 29699
rect 34655 29696 34667 29699
rect 34698 29696 34704 29708
rect 34655 29668 34704 29696
rect 34655 29665 34667 29668
rect 34609 29659 34667 29665
rect 34698 29656 34704 29668
rect 34756 29656 34762 29708
rect 33318 29628 33324 29640
rect 33106 29600 33324 29628
rect 28445 29591 28503 29597
rect 33318 29588 33324 29600
rect 33376 29628 33382 29640
rect 33413 29631 33471 29637
rect 33413 29628 33425 29631
rect 33376 29600 33425 29628
rect 33376 29588 33382 29600
rect 33413 29597 33425 29600
rect 33459 29628 33471 29631
rect 34977 29631 35035 29637
rect 34977 29628 34989 29631
rect 33459 29600 34989 29628
rect 33459 29597 33471 29600
rect 33413 29591 33471 29597
rect 34977 29597 34989 29600
rect 35023 29628 35035 29631
rect 35342 29628 35348 29640
rect 35023 29600 35348 29628
rect 35023 29597 35035 29600
rect 34977 29591 35035 29597
rect 35342 29588 35348 29600
rect 35400 29588 35406 29640
rect 19024 29532 21312 29560
rect 19024 29520 19030 29532
rect 24670 29520 24676 29572
rect 24728 29560 24734 29572
rect 24857 29563 24915 29569
rect 24857 29560 24869 29563
rect 24728 29532 24869 29560
rect 24728 29520 24734 29532
rect 24857 29529 24869 29532
rect 24903 29560 24915 29563
rect 27341 29563 27399 29569
rect 27341 29560 27353 29563
rect 24903 29532 27353 29560
rect 24903 29529 24915 29532
rect 24857 29523 24915 29529
rect 27341 29529 27353 29532
rect 27387 29560 27399 29563
rect 29638 29560 29644 29572
rect 27387 29532 29644 29560
rect 27387 29529 27399 29532
rect 27341 29523 27399 29529
rect 29638 29520 29644 29532
rect 29696 29520 29702 29572
rect 33042 29520 33048 29572
rect 33100 29560 33106 29572
rect 33505 29563 33563 29569
rect 33505 29560 33517 29563
rect 33100 29532 33517 29560
rect 33100 29520 33106 29532
rect 33505 29529 33517 29532
rect 33551 29529 33563 29563
rect 33505 29523 33563 29529
rect 33962 29520 33968 29572
rect 34020 29560 34026 29572
rect 35069 29563 35127 29569
rect 35069 29560 35081 29563
rect 34020 29532 35081 29560
rect 34020 29520 34026 29532
rect 35069 29529 35081 29532
rect 35115 29529 35127 29563
rect 35452 29560 35480 29736
rect 37461 29733 37473 29736
rect 37507 29764 37519 29767
rect 37550 29764 37556 29776
rect 37507 29736 37556 29764
rect 37507 29733 37519 29736
rect 37461 29727 37519 29733
rect 37550 29724 37556 29736
rect 37608 29724 37614 29776
rect 41871 29767 41929 29773
rect 41871 29733 41883 29767
rect 41917 29764 41929 29767
rect 42518 29764 42524 29776
rect 41917 29736 42524 29764
rect 41917 29733 41929 29736
rect 41871 29727 41929 29733
rect 42518 29724 42524 29736
rect 42576 29764 42582 29776
rect 42766 29764 42794 29804
rect 43717 29801 43729 29804
rect 43763 29801 43775 29835
rect 43717 29795 43775 29801
rect 44269 29835 44327 29841
rect 44269 29801 44281 29835
rect 44315 29832 44327 29835
rect 44634 29832 44640 29844
rect 44315 29804 44640 29832
rect 44315 29801 44327 29804
rect 44269 29795 44327 29801
rect 44634 29792 44640 29804
rect 44692 29832 44698 29844
rect 44913 29835 44971 29841
rect 44913 29832 44925 29835
rect 44692 29804 44925 29832
rect 44692 29792 44698 29804
rect 44913 29801 44925 29804
rect 44959 29832 44971 29835
rect 44959 29804 45324 29832
rect 44959 29801 44971 29804
rect 44913 29795 44971 29801
rect 45296 29773 45324 29804
rect 42576 29736 42794 29764
rect 45281 29767 45339 29773
rect 42576 29724 42582 29736
rect 45281 29733 45293 29767
rect 45327 29733 45339 29767
rect 45281 29727 45339 29733
rect 36630 29696 36636 29708
rect 36591 29668 36636 29696
rect 36630 29656 36636 29668
rect 36688 29656 36694 29708
rect 40126 29696 40132 29708
rect 40087 29668 40132 29696
rect 40126 29656 40132 29668
rect 40184 29656 40190 29708
rect 40678 29656 40684 29708
rect 40736 29696 40742 29708
rect 41506 29696 41512 29708
rect 40736 29668 41512 29696
rect 40736 29656 40742 29668
rect 41506 29656 41512 29668
rect 41564 29656 41570 29708
rect 42794 29656 42800 29708
rect 42852 29696 42858 29708
rect 43346 29696 43352 29708
rect 42852 29668 42897 29696
rect 43307 29668 43352 29696
rect 42852 29656 42858 29668
rect 43346 29656 43352 29668
rect 43404 29656 43410 29708
rect 46934 29696 46940 29708
rect 46895 29668 46940 29696
rect 46934 29656 46940 29668
rect 46992 29656 46998 29708
rect 47210 29656 47216 29708
rect 47268 29696 47274 29708
rect 47305 29699 47363 29705
rect 47305 29696 47317 29699
rect 47268 29668 47317 29696
rect 47268 29656 47274 29668
rect 47305 29665 47317 29668
rect 47351 29665 47363 29699
rect 47305 29659 47363 29665
rect 38378 29628 38384 29640
rect 38339 29600 38384 29628
rect 38378 29588 38384 29600
rect 38436 29588 38442 29640
rect 45189 29631 45247 29637
rect 45189 29597 45201 29631
rect 45235 29628 45247 29631
rect 45370 29628 45376 29640
rect 45235 29600 45376 29628
rect 45235 29597 45247 29600
rect 45189 29591 45247 29597
rect 45370 29588 45376 29600
rect 45428 29588 45434 29640
rect 45554 29628 45560 29640
rect 45515 29600 45560 29628
rect 45554 29588 45560 29600
rect 45612 29588 45618 29640
rect 37734 29560 37740 29572
rect 35069 29523 35127 29529
rect 35268 29532 37740 29560
rect 19935 29495 19993 29501
rect 19935 29461 19947 29495
rect 19981 29492 19993 29495
rect 20162 29492 20168 29504
rect 19981 29464 20168 29492
rect 19981 29461 19993 29464
rect 19935 29455 19993 29461
rect 20162 29452 20168 29464
rect 20220 29452 20226 29504
rect 26326 29492 26332 29504
rect 26287 29464 26332 29492
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 29365 29495 29423 29501
rect 29365 29461 29377 29495
rect 29411 29492 29423 29495
rect 29454 29492 29460 29504
rect 29411 29464 29460 29492
rect 29411 29461 29423 29464
rect 29365 29455 29423 29461
rect 29454 29452 29460 29464
rect 29512 29452 29518 29504
rect 32953 29495 33011 29501
rect 32953 29461 32965 29495
rect 32999 29492 33011 29495
rect 33226 29492 33232 29504
rect 32999 29464 33232 29492
rect 32999 29461 33011 29464
rect 32953 29455 33011 29461
rect 33226 29452 33232 29464
rect 33284 29452 33290 29504
rect 33321 29495 33379 29501
rect 33321 29461 33333 29495
rect 33367 29492 33379 29495
rect 34330 29492 34336 29504
rect 33367 29464 34336 29492
rect 33367 29461 33379 29464
rect 33321 29455 33379 29461
rect 34330 29452 34336 29464
rect 34388 29452 34394 29504
rect 34514 29452 34520 29504
rect 34572 29492 34578 29504
rect 34747 29495 34805 29501
rect 34747 29492 34759 29495
rect 34572 29464 34759 29492
rect 34572 29452 34578 29464
rect 34747 29461 34759 29464
rect 34793 29461 34805 29495
rect 34747 29455 34805 29461
rect 34885 29495 34943 29501
rect 34885 29461 34897 29495
rect 34931 29492 34943 29495
rect 35268 29492 35296 29532
rect 37734 29520 37740 29532
rect 37792 29520 37798 29572
rect 40310 29560 40316 29572
rect 40271 29532 40316 29560
rect 40310 29520 40316 29532
rect 40368 29520 40374 29572
rect 34931 29464 35296 29492
rect 34931 29461 34943 29464
rect 34885 29455 34943 29461
rect 36354 29452 36360 29504
rect 36412 29492 36418 29504
rect 37185 29495 37243 29501
rect 37185 29492 37197 29495
rect 36412 29464 37197 29492
rect 36412 29452 36418 29464
rect 37185 29461 37197 29464
rect 37231 29492 37243 29495
rect 37458 29492 37464 29504
rect 37231 29464 37464 29492
rect 37231 29461 37243 29464
rect 37185 29455 37243 29461
rect 37458 29452 37464 29464
rect 37516 29452 37522 29504
rect 38010 29492 38016 29504
rect 37971 29464 38016 29492
rect 38010 29452 38016 29464
rect 38068 29452 38074 29504
rect 39574 29492 39580 29504
rect 39535 29464 39580 29492
rect 39574 29452 39580 29464
rect 39632 29452 39638 29504
rect 46842 29492 46848 29504
rect 46803 29464 46848 29492
rect 46842 29452 46848 29464
rect 46900 29452 46906 29504
rect 1104 29402 48852 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 48852 29402
rect 1104 29328 48852 29350
rect 13173 29291 13231 29297
rect 13173 29257 13185 29291
rect 13219 29288 13231 29291
rect 13354 29288 13360 29300
rect 13219 29260 13360 29288
rect 13219 29257 13231 29260
rect 13173 29251 13231 29257
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 14737 29291 14795 29297
rect 14737 29257 14749 29291
rect 14783 29288 14795 29291
rect 15194 29288 15200 29300
rect 14783 29260 15200 29288
rect 14783 29257 14795 29260
rect 14737 29251 14795 29257
rect 15194 29248 15200 29260
rect 15252 29288 15258 29300
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15252 29260 16037 29288
rect 15252 29248 15258 29260
rect 16025 29257 16037 29260
rect 16071 29288 16083 29291
rect 17773 29291 17831 29297
rect 17773 29288 17785 29291
rect 16071 29260 17785 29288
rect 16071 29257 16083 29260
rect 16025 29251 16083 29257
rect 17773 29257 17785 29260
rect 17819 29257 17831 29291
rect 17773 29251 17831 29257
rect 16666 29180 16672 29232
rect 16724 29220 16730 29232
rect 17129 29223 17187 29229
rect 17129 29220 17141 29223
rect 16724 29192 17141 29220
rect 16724 29180 16730 29192
rect 17129 29189 17141 29192
rect 17175 29220 17187 29223
rect 17218 29220 17224 29232
rect 17175 29192 17224 29220
rect 17175 29189 17187 29192
rect 17129 29183 17187 29189
rect 17218 29180 17224 29192
rect 17276 29180 17282 29232
rect 14366 29112 14372 29164
rect 14424 29152 14430 29164
rect 14829 29155 14887 29161
rect 14829 29152 14841 29155
rect 14424 29124 14841 29152
rect 14424 29112 14430 29124
rect 14829 29121 14841 29124
rect 14875 29121 14887 29155
rect 14829 29115 14887 29121
rect 13354 29084 13360 29096
rect 13315 29056 13360 29084
rect 13354 29044 13360 29056
rect 13412 29044 13418 29096
rect 13814 29044 13820 29096
rect 13872 29084 13878 29096
rect 14001 29087 14059 29093
rect 13872 29056 13917 29084
rect 13872 29044 13878 29056
rect 14001 29053 14013 29087
rect 14047 29084 14059 29087
rect 15286 29084 15292 29096
rect 14047 29056 15292 29084
rect 14047 29053 14059 29056
rect 14001 29047 14059 29053
rect 15286 29044 15292 29056
rect 15344 29044 15350 29096
rect 16945 29087 17003 29093
rect 16945 29053 16957 29087
rect 16991 29084 17003 29087
rect 16991 29056 17540 29084
rect 16991 29053 17003 29056
rect 16945 29047 17003 29053
rect 14369 28951 14427 28957
rect 14369 28917 14381 28951
rect 14415 28948 14427 28951
rect 14550 28948 14556 28960
rect 14415 28920 14556 28948
rect 14415 28917 14427 28920
rect 14369 28911 14427 28917
rect 14550 28908 14556 28920
rect 14608 28908 14614 28960
rect 15194 28948 15200 28960
rect 15155 28920 15200 28948
rect 15194 28908 15200 28920
rect 15252 28908 15258 28960
rect 15749 28951 15807 28957
rect 15749 28917 15761 28951
rect 15795 28948 15807 28951
rect 15930 28948 15936 28960
rect 15795 28920 15936 28948
rect 15795 28917 15807 28920
rect 15749 28911 15807 28917
rect 15930 28908 15936 28920
rect 15988 28908 15994 28960
rect 17512 28957 17540 29056
rect 17788 29016 17816 29251
rect 18414 29248 18420 29300
rect 18472 29288 18478 29300
rect 18969 29291 19027 29297
rect 18969 29288 18981 29291
rect 18472 29260 18981 29288
rect 18472 29248 18478 29260
rect 18969 29257 18981 29260
rect 19015 29257 19027 29291
rect 18969 29251 19027 29257
rect 19978 29248 19984 29300
rect 20036 29288 20042 29300
rect 20165 29291 20223 29297
rect 20165 29288 20177 29291
rect 20036 29260 20177 29288
rect 20036 29248 20042 29260
rect 20165 29257 20177 29260
rect 20211 29257 20223 29291
rect 20165 29251 20223 29257
rect 20625 29291 20683 29297
rect 20625 29257 20637 29291
rect 20671 29288 20683 29291
rect 21082 29288 21088 29300
rect 20671 29260 21088 29288
rect 20671 29257 20683 29260
rect 20625 29251 20683 29257
rect 21082 29248 21088 29260
rect 21140 29288 21146 29300
rect 21729 29291 21787 29297
rect 21729 29288 21741 29291
rect 21140 29260 21741 29288
rect 21140 29248 21146 29260
rect 21729 29257 21741 29260
rect 21775 29257 21787 29291
rect 21729 29251 21787 29257
rect 22465 29291 22523 29297
rect 22465 29257 22477 29291
rect 22511 29288 22523 29291
rect 23198 29288 23204 29300
rect 22511 29260 23204 29288
rect 22511 29257 22523 29260
rect 22465 29251 22523 29257
rect 23198 29248 23204 29260
rect 23256 29248 23262 29300
rect 24118 29248 24124 29300
rect 24176 29288 24182 29300
rect 24305 29291 24363 29297
rect 24305 29288 24317 29291
rect 24176 29260 24317 29288
rect 24176 29248 24182 29260
rect 24305 29257 24317 29260
rect 24351 29257 24363 29291
rect 24670 29288 24676 29300
rect 24631 29260 24676 29288
rect 24305 29251 24363 29257
rect 24670 29248 24676 29260
rect 24728 29248 24734 29300
rect 24762 29248 24768 29300
rect 24820 29288 24826 29300
rect 25041 29291 25099 29297
rect 25041 29288 25053 29291
rect 24820 29260 25053 29288
rect 24820 29248 24826 29260
rect 25041 29257 25053 29260
rect 25087 29257 25099 29291
rect 25041 29251 25099 29257
rect 26881 29291 26939 29297
rect 26881 29257 26893 29291
rect 26927 29288 26939 29291
rect 27154 29288 27160 29300
rect 26927 29260 27160 29288
rect 26927 29257 26939 29260
rect 26881 29251 26939 29257
rect 27154 29248 27160 29260
rect 27212 29248 27218 29300
rect 28350 29288 28356 29300
rect 28311 29260 28356 29288
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 29089 29291 29147 29297
rect 29089 29257 29101 29291
rect 29135 29288 29147 29291
rect 30006 29288 30012 29300
rect 29135 29260 30012 29288
rect 29135 29257 29147 29260
rect 29089 29251 29147 29257
rect 18782 29180 18788 29232
rect 18840 29220 18846 29232
rect 19245 29223 19303 29229
rect 19245 29220 19257 29223
rect 18840 29192 19257 29220
rect 18840 29180 18846 29192
rect 19245 29189 19257 29192
rect 19291 29189 19303 29223
rect 21358 29220 21364 29232
rect 21319 29192 21364 29220
rect 19245 29183 19303 29189
rect 21358 29180 21364 29192
rect 21416 29180 21422 29232
rect 20162 29112 20168 29164
rect 20220 29152 20226 29164
rect 20809 29155 20867 29161
rect 20809 29152 20821 29155
rect 20220 29124 20821 29152
rect 20220 29112 20226 29124
rect 20809 29121 20821 29124
rect 20855 29152 20867 29155
rect 21266 29152 21272 29164
rect 20855 29124 21272 29152
rect 20855 29121 20867 29124
rect 20809 29115 20867 29121
rect 21266 29112 21272 29124
rect 21324 29112 21330 29164
rect 26326 29152 26332 29164
rect 26287 29124 26332 29152
rect 26326 29112 26332 29124
rect 26384 29112 26390 29164
rect 26878 29112 26884 29164
rect 26936 29152 26942 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 26936 29124 27169 29152
rect 26936 29112 26942 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 18046 29084 18052 29096
rect 18007 29056 18052 29084
rect 18046 29044 18052 29056
rect 18104 29044 18110 29096
rect 22557 29087 22615 29093
rect 22557 29053 22569 29087
rect 22603 29084 22615 29087
rect 23912 29087 23970 29093
rect 22603 29056 23474 29084
rect 22603 29053 22615 29056
rect 22557 29047 22615 29053
rect 18370 29019 18428 29025
rect 18370 29016 18382 29019
rect 17788 28988 18382 29016
rect 18370 28985 18382 28988
rect 18416 28985 18428 29019
rect 19886 29016 19892 29028
rect 19847 28988 19892 29016
rect 18370 28979 18428 28985
rect 19886 28976 19892 28988
rect 19944 28976 19950 29028
rect 20901 29019 20959 29025
rect 20901 28985 20913 29019
rect 20947 29016 20959 29019
rect 21082 29016 21088 29028
rect 20947 28988 21088 29016
rect 20947 28985 20959 28988
rect 20901 28979 20959 28985
rect 21082 28976 21088 28988
rect 21140 28976 21146 29028
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22922 29016 22928 29028
rect 21876 28988 22928 29016
rect 21876 28976 21882 28988
rect 22922 28976 22928 28988
rect 22980 29016 22986 29028
rect 23017 29019 23075 29025
rect 23017 29016 23029 29019
rect 22980 28988 23029 29016
rect 22980 28976 22986 28988
rect 23017 28985 23029 28988
rect 23063 28985 23075 29019
rect 23017 28979 23075 28985
rect 23446 28960 23474 29056
rect 23912 29053 23924 29087
rect 23958 29084 23970 29087
rect 24670 29084 24676 29096
rect 23958 29056 24676 29084
rect 23958 29053 23970 29056
rect 23912 29047 23970 29053
rect 24670 29044 24676 29056
rect 24728 29044 24734 29096
rect 25777 29087 25835 29093
rect 25777 29053 25789 29087
rect 25823 29053 25835 29087
rect 25777 29047 25835 29053
rect 26237 29087 26295 29093
rect 26237 29053 26249 29087
rect 26283 29053 26295 29087
rect 26237 29047 26295 29053
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29084 28227 29087
rect 29104 29084 29132 29251
rect 30006 29248 30012 29260
rect 30064 29248 30070 29300
rect 32582 29248 32588 29300
rect 32640 29288 32646 29300
rect 32640 29260 33548 29288
rect 32640 29248 32646 29260
rect 33520 29232 33548 29260
rect 35894 29248 35900 29300
rect 35952 29288 35958 29300
rect 36265 29291 36323 29297
rect 36265 29288 36277 29291
rect 35952 29260 36277 29288
rect 35952 29248 35958 29260
rect 36265 29257 36277 29260
rect 36311 29257 36323 29291
rect 36265 29251 36323 29257
rect 36998 29248 37004 29300
rect 37056 29288 37062 29300
rect 37461 29291 37519 29297
rect 37461 29288 37473 29291
rect 37056 29260 37473 29288
rect 37056 29248 37062 29260
rect 37461 29257 37473 29260
rect 37507 29257 37519 29291
rect 37461 29251 37519 29257
rect 33502 29220 33508 29232
rect 33463 29192 33508 29220
rect 33502 29180 33508 29192
rect 33560 29180 33566 29232
rect 35161 29223 35219 29229
rect 35161 29189 35173 29223
rect 35207 29220 35219 29223
rect 37274 29220 37280 29232
rect 35207 29192 37280 29220
rect 35207 29189 35219 29192
rect 35161 29183 35219 29189
rect 37274 29180 37280 29192
rect 37332 29180 37338 29232
rect 29638 29152 29644 29164
rect 29599 29124 29644 29152
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 33137 29155 33195 29161
rect 33137 29121 33149 29155
rect 33183 29152 33195 29155
rect 33597 29155 33655 29161
rect 33597 29152 33609 29155
rect 33183 29124 33609 29152
rect 33183 29121 33195 29124
rect 33137 29115 33195 29121
rect 33597 29121 33609 29124
rect 33643 29152 33655 29155
rect 33778 29152 33784 29164
rect 33643 29124 33784 29152
rect 33643 29121 33655 29124
rect 33597 29115 33655 29121
rect 33778 29112 33784 29124
rect 33836 29112 33842 29164
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 34701 29155 34759 29161
rect 34701 29152 34713 29155
rect 34572 29124 34713 29152
rect 34572 29112 34578 29124
rect 34701 29121 34713 29124
rect 34747 29152 34759 29155
rect 35250 29152 35256 29164
rect 34747 29124 35256 29152
rect 34747 29121 34759 29124
rect 34701 29115 34759 29121
rect 35250 29112 35256 29124
rect 35308 29152 35314 29164
rect 35897 29155 35955 29161
rect 35897 29152 35909 29155
rect 35308 29124 35909 29152
rect 35308 29112 35314 29124
rect 35897 29121 35909 29124
rect 35943 29152 35955 29155
rect 36136 29155 36194 29161
rect 36136 29152 36148 29155
rect 35943 29124 36148 29152
rect 35943 29121 35955 29124
rect 35897 29115 35955 29121
rect 36136 29121 36148 29124
rect 36182 29152 36194 29155
rect 36262 29152 36268 29164
rect 36182 29124 36268 29152
rect 36182 29121 36194 29124
rect 36136 29115 36194 29121
rect 36262 29112 36268 29124
rect 36320 29112 36326 29164
rect 36354 29112 36360 29164
rect 36412 29152 36418 29164
rect 36412 29124 36457 29152
rect 36412 29112 36418 29124
rect 36630 29112 36636 29164
rect 36688 29152 36694 29164
rect 36998 29152 37004 29164
rect 36688 29124 37004 29152
rect 36688 29112 36694 29124
rect 36998 29112 37004 29124
rect 37056 29112 37062 29164
rect 28215 29056 29132 29084
rect 31481 29087 31539 29093
rect 28215 29053 28227 29056
rect 28169 29047 28227 29053
rect 31481 29053 31493 29087
rect 31527 29053 31539 29087
rect 31662 29084 31668 29096
rect 31623 29056 31668 29084
rect 31481 29047 31539 29053
rect 17497 28951 17555 28957
rect 17497 28917 17509 28951
rect 17543 28948 17555 28951
rect 17586 28948 17592 28960
rect 17543 28920 17592 28948
rect 17543 28917 17555 28920
rect 17497 28911 17555 28917
rect 17586 28908 17592 28920
rect 17644 28908 17650 28960
rect 22646 28908 22652 28960
rect 22704 28948 22710 28960
rect 22741 28951 22799 28957
rect 22741 28948 22753 28951
rect 22704 28920 22753 28948
rect 22704 28908 22710 28920
rect 22741 28917 22753 28920
rect 22787 28917 22799 28951
rect 23446 28920 23480 28960
rect 22741 28911 22799 28917
rect 23474 28908 23480 28920
rect 23532 28948 23538 28960
rect 23983 28951 24041 28957
rect 23532 28920 23577 28948
rect 23532 28908 23538 28920
rect 23983 28917 23995 28951
rect 24029 28948 24041 28951
rect 24118 28948 24124 28960
rect 24029 28920 24124 28948
rect 24029 28917 24041 28920
rect 23983 28911 24041 28917
rect 24118 28908 24124 28920
rect 24176 28908 24182 28960
rect 25685 28951 25743 28957
rect 25685 28917 25697 28951
rect 25731 28948 25743 28951
rect 25792 28948 25820 29047
rect 25866 28976 25872 29028
rect 25924 29016 25930 29028
rect 26252 29016 26280 29047
rect 28350 29016 28356 29028
rect 25924 28988 28356 29016
rect 25924 28976 25930 28988
rect 28350 28976 28356 28988
rect 28408 28976 28414 29028
rect 28442 28976 28448 29028
rect 28500 29016 28506 29028
rect 29362 29016 29368 29028
rect 28500 28988 29368 29016
rect 28500 28976 28506 28988
rect 29362 28976 29368 28988
rect 29420 28976 29426 29028
rect 29454 28976 29460 29028
rect 29512 29016 29518 29028
rect 30745 29019 30803 29025
rect 29512 28988 29557 29016
rect 29512 28976 29518 28988
rect 30745 28985 30757 29019
rect 30791 29016 30803 29019
rect 31018 29016 31024 29028
rect 30791 28988 31024 29016
rect 30791 28985 30803 28988
rect 30745 28979 30803 28985
rect 31018 28976 31024 28988
rect 31076 29016 31082 29028
rect 31113 29019 31171 29025
rect 31113 29016 31125 29019
rect 31076 28988 31125 29016
rect 31076 28976 31082 28988
rect 31113 28985 31125 28988
rect 31159 29016 31171 29019
rect 31496 29016 31524 29047
rect 31662 29044 31668 29056
rect 31720 29044 31726 29096
rect 32769 29087 32827 29093
rect 32769 29053 32781 29087
rect 32815 29084 32827 29087
rect 33376 29087 33434 29093
rect 33376 29084 33388 29087
rect 32815 29056 33388 29084
rect 32815 29053 32827 29056
rect 32769 29047 32827 29053
rect 33376 29053 33388 29056
rect 33422 29084 33434 29087
rect 33686 29084 33692 29096
rect 33422 29056 33692 29084
rect 33422 29053 33434 29056
rect 33376 29047 33434 29053
rect 33686 29044 33692 29056
rect 33744 29044 33750 29096
rect 34977 29087 35035 29093
rect 34977 29084 34989 29087
rect 34256 29056 34989 29084
rect 31570 29016 31576 29028
rect 31159 28988 31576 29016
rect 31159 28985 31171 28988
rect 31113 28979 31171 28985
rect 31570 28976 31576 28988
rect 31628 28976 31634 29028
rect 32401 29019 32459 29025
rect 32401 28985 32413 29019
rect 32447 29016 32459 29019
rect 32950 29016 32956 29028
rect 32447 28988 32956 29016
rect 32447 28985 32459 28988
rect 32401 28979 32459 28985
rect 32950 28976 32956 28988
rect 33008 29016 33014 29028
rect 33229 29019 33287 29025
rect 33229 29016 33241 29019
rect 33008 28988 33241 29016
rect 33008 28976 33014 28988
rect 33229 28985 33241 28988
rect 33275 28985 33287 29019
rect 33229 28979 33287 28985
rect 34256 28960 34284 29056
rect 34977 29053 34989 29056
rect 35023 29053 35035 29087
rect 37476 29084 37504 29251
rect 43346 29248 43352 29300
rect 43404 29288 43410 29300
rect 43717 29291 43775 29297
rect 43717 29288 43729 29291
rect 43404 29260 43729 29288
rect 43404 29248 43410 29260
rect 43717 29257 43729 29260
rect 43763 29257 43775 29291
rect 43717 29251 43775 29257
rect 44361 29291 44419 29297
rect 44361 29257 44373 29291
rect 44407 29288 44419 29291
rect 44634 29288 44640 29300
rect 44407 29260 44640 29288
rect 44407 29257 44419 29260
rect 44361 29251 44419 29257
rect 44634 29248 44640 29260
rect 44692 29288 44698 29300
rect 45465 29291 45523 29297
rect 45465 29288 45477 29291
rect 44692 29260 45477 29288
rect 44692 29248 44698 29260
rect 45465 29257 45477 29260
rect 45511 29257 45523 29291
rect 47026 29288 47032 29300
rect 46987 29260 47032 29288
rect 45465 29251 45523 29257
rect 47026 29248 47032 29260
rect 47084 29248 47090 29300
rect 39022 29180 39028 29232
rect 39080 29220 39086 29232
rect 39853 29223 39911 29229
rect 39853 29220 39865 29223
rect 39080 29192 39865 29220
rect 39080 29180 39086 29192
rect 39853 29189 39865 29192
rect 39899 29220 39911 29223
rect 40126 29220 40132 29232
rect 39899 29192 40132 29220
rect 39899 29189 39911 29192
rect 39853 29183 39911 29189
rect 40126 29180 40132 29192
rect 40184 29180 40190 29232
rect 41877 29223 41935 29229
rect 41877 29189 41889 29223
rect 41923 29220 41935 29223
rect 42518 29220 42524 29232
rect 41923 29192 42524 29220
rect 41923 29189 41935 29192
rect 41877 29183 41935 29189
rect 42518 29180 42524 29192
rect 42576 29180 42582 29232
rect 46661 29223 46719 29229
rect 46661 29189 46673 29223
rect 46707 29220 46719 29223
rect 46934 29220 46940 29232
rect 46707 29192 46940 29220
rect 46707 29189 46719 29192
rect 46661 29183 46719 29189
rect 46934 29180 46940 29192
rect 46992 29180 46998 29232
rect 38010 29112 38016 29164
rect 38068 29152 38074 29164
rect 39574 29152 39580 29164
rect 38068 29124 39580 29152
rect 38068 29112 38074 29124
rect 38212 29093 38240 29124
rect 39574 29112 39580 29124
rect 39632 29112 39638 29164
rect 40494 29152 40500 29164
rect 40455 29124 40500 29152
rect 40494 29112 40500 29124
rect 40552 29112 40558 29164
rect 42150 29112 42156 29164
rect 42208 29152 42214 29164
rect 42334 29152 42340 29164
rect 42208 29124 42340 29152
rect 42208 29112 42214 29124
rect 42334 29112 42340 29124
rect 42392 29112 42398 29164
rect 42981 29155 43039 29161
rect 42981 29121 42993 29155
rect 43027 29152 43039 29155
rect 43070 29152 43076 29164
rect 43027 29124 43076 29152
rect 43027 29121 43039 29124
rect 42981 29115 43039 29121
rect 43070 29112 43076 29124
rect 43128 29112 43134 29164
rect 44545 29155 44603 29161
rect 44545 29121 44557 29155
rect 44591 29152 44603 29155
rect 44818 29152 44824 29164
rect 44591 29124 44824 29152
rect 44591 29121 44603 29124
rect 44545 29115 44603 29121
rect 44818 29112 44824 29124
rect 44876 29112 44882 29164
rect 44910 29112 44916 29164
rect 44968 29152 44974 29164
rect 44968 29124 45013 29152
rect 44968 29112 44974 29124
rect 37645 29087 37703 29093
rect 37645 29084 37657 29087
rect 37476 29056 37657 29084
rect 34977 29047 35035 29053
rect 37645 29053 37657 29056
rect 37691 29053 37703 29087
rect 37645 29047 37703 29053
rect 38197 29087 38255 29093
rect 38197 29053 38209 29087
rect 38243 29053 38255 29087
rect 38378 29084 38384 29096
rect 38339 29056 38384 29084
rect 38197 29047 38255 29053
rect 38378 29044 38384 29056
rect 38436 29044 38442 29096
rect 39209 29087 39267 29093
rect 39209 29053 39221 29087
rect 39255 29053 39267 29087
rect 39209 29047 39267 29053
rect 41417 29087 41475 29093
rect 41417 29053 41429 29087
rect 41463 29084 41475 29087
rect 42061 29087 42119 29093
rect 42061 29084 42073 29087
rect 41463 29056 42073 29084
rect 41463 29053 41475 29056
rect 41417 29047 41475 29053
rect 42061 29053 42073 29056
rect 42107 29053 42119 29087
rect 42061 29047 42119 29053
rect 45925 29087 45983 29093
rect 45925 29053 45937 29087
rect 45971 29084 45983 29087
rect 47210 29084 47216 29096
rect 45971 29056 47216 29084
rect 45971 29053 45983 29056
rect 45925 29047 45983 29053
rect 34330 28976 34336 29028
rect 34388 29016 34394 29028
rect 34514 29016 34520 29028
rect 34388 28988 34520 29016
rect 34388 28976 34394 28988
rect 34514 28976 34520 28988
rect 34572 28976 34578 29028
rect 34698 28976 34704 29028
rect 34756 29016 34762 29028
rect 35529 29019 35587 29025
rect 35529 29016 35541 29019
rect 34756 28988 35541 29016
rect 34756 28976 34762 28988
rect 35529 28985 35541 28988
rect 35575 29016 35587 29019
rect 35989 29019 36047 29025
rect 35989 29016 36001 29019
rect 35575 28988 36001 29016
rect 35575 28985 35587 28988
rect 35529 28979 35587 28985
rect 35989 28985 36001 28988
rect 36035 29016 36047 29019
rect 36078 29016 36084 29028
rect 36035 28988 36084 29016
rect 36035 28985 36047 28988
rect 35989 28979 36047 28985
rect 36078 28976 36084 28988
rect 36136 28976 36142 29028
rect 36725 29019 36783 29025
rect 36725 28985 36737 29019
rect 36771 29016 36783 29019
rect 39025 29019 39083 29025
rect 39025 29016 39037 29019
rect 36771 28988 39037 29016
rect 36771 28985 36783 28988
rect 36725 28979 36783 28985
rect 39025 28985 39037 28988
rect 39071 29016 39083 29019
rect 39224 29016 39252 29047
rect 39071 28988 39252 29016
rect 40859 29019 40917 29025
rect 39071 28985 39083 28988
rect 39025 28979 39083 28985
rect 40859 28985 40871 29019
rect 40905 28985 40917 29019
rect 40859 28979 40917 28985
rect 26418 28948 26424 28960
rect 25731 28920 26424 28948
rect 25731 28917 25743 28920
rect 25685 28911 25743 28917
rect 26418 28908 26424 28920
rect 26476 28908 26482 28960
rect 28077 28951 28135 28957
rect 28077 28917 28089 28951
rect 28123 28948 28135 28951
rect 28258 28948 28264 28960
rect 28123 28920 28264 28948
rect 28123 28917 28135 28920
rect 28077 28911 28135 28917
rect 28258 28908 28264 28920
rect 28316 28908 28322 28960
rect 28718 28948 28724 28960
rect 28679 28920 28724 28948
rect 28718 28908 28724 28920
rect 28776 28908 28782 28960
rect 31478 28948 31484 28960
rect 31439 28920 31484 28948
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 31754 28908 31760 28960
rect 31812 28948 31818 28960
rect 33873 28951 33931 28957
rect 33873 28948 33885 28951
rect 31812 28920 33885 28948
rect 31812 28908 31818 28920
rect 33873 28917 33885 28920
rect 33919 28917 33931 28951
rect 34238 28948 34244 28960
rect 34199 28920 34244 28948
rect 33873 28911 33931 28917
rect 34238 28908 34244 28920
rect 34296 28908 34302 28960
rect 38654 28908 38660 28960
rect 38712 28948 38718 28960
rect 38749 28951 38807 28957
rect 38749 28948 38761 28951
rect 38712 28920 38761 28948
rect 38712 28908 38718 28920
rect 38749 28917 38761 28920
rect 38795 28948 38807 28951
rect 38930 28948 38936 28960
rect 38795 28920 38936 28948
rect 38795 28917 38807 28920
rect 38749 28911 38807 28917
rect 38930 28908 38936 28920
rect 38988 28908 38994 28960
rect 39390 28948 39396 28960
rect 39351 28920 39396 28948
rect 39390 28908 39396 28920
rect 39448 28908 39454 28960
rect 40218 28948 40224 28960
rect 40179 28920 40224 28948
rect 40218 28908 40224 28920
rect 40276 28948 40282 28960
rect 40880 28948 40908 28979
rect 41693 28951 41751 28957
rect 41693 28948 41705 28951
rect 40276 28920 41705 28948
rect 40276 28908 40282 28920
rect 41693 28917 41705 28920
rect 41739 28948 41751 28951
rect 41877 28951 41935 28957
rect 41877 28948 41889 28951
rect 41739 28920 41889 28948
rect 41739 28917 41751 28920
rect 41693 28911 41751 28917
rect 41877 28917 41889 28920
rect 41923 28917 41935 28951
rect 42076 28948 42104 29047
rect 47210 29044 47216 29056
rect 47268 29044 47274 29096
rect 42429 29019 42487 29025
rect 42429 28985 42441 29019
rect 42475 28985 42487 29019
rect 44634 29016 44640 29028
rect 44595 28988 44640 29016
rect 42429 28979 42487 28985
rect 42444 28948 42472 28979
rect 44634 28976 44640 28988
rect 44692 28976 44698 29028
rect 42076 28920 42472 28948
rect 41877 28911 41935 28917
rect 42518 28908 42524 28960
rect 42576 28948 42582 28960
rect 43349 28951 43407 28957
rect 43349 28948 43361 28951
rect 42576 28920 43361 28948
rect 42576 28908 42582 28920
rect 43349 28917 43361 28920
rect 43395 28917 43407 28951
rect 43349 28911 43407 28917
rect 1104 28858 48852 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 48852 28858
rect 1104 28784 48852 28806
rect 13078 28704 13084 28756
rect 13136 28744 13142 28756
rect 13265 28747 13323 28753
rect 13265 28744 13277 28747
rect 13136 28716 13277 28744
rect 13136 28704 13142 28716
rect 13265 28713 13277 28716
rect 13311 28744 13323 28747
rect 13633 28747 13691 28753
rect 13633 28744 13645 28747
rect 13311 28716 13645 28744
rect 13311 28713 13323 28716
rect 13265 28707 13323 28713
rect 13633 28713 13645 28716
rect 13679 28713 13691 28747
rect 13633 28707 13691 28713
rect 13648 28676 13676 28707
rect 13722 28704 13728 28756
rect 13780 28744 13786 28756
rect 14829 28747 14887 28753
rect 14829 28744 14841 28747
rect 13780 28716 14841 28744
rect 13780 28704 13786 28716
rect 14829 28713 14841 28716
rect 14875 28713 14887 28747
rect 14829 28707 14887 28713
rect 15286 28704 15292 28756
rect 15344 28744 15350 28756
rect 15473 28747 15531 28753
rect 15473 28744 15485 28747
rect 15344 28716 15485 28744
rect 15344 28704 15350 28716
rect 15473 28713 15485 28716
rect 15519 28713 15531 28747
rect 16390 28744 16396 28756
rect 15473 28707 15531 28713
rect 15580 28716 16396 28744
rect 13814 28676 13820 28688
rect 13648 28648 13820 28676
rect 13814 28636 13820 28648
rect 13872 28676 13878 28688
rect 15580 28676 15608 28716
rect 16390 28704 16396 28716
rect 16448 28744 16454 28756
rect 18414 28744 18420 28756
rect 16448 28716 17816 28744
rect 18375 28716 18420 28744
rect 16448 28704 16454 28716
rect 15930 28676 15936 28688
rect 13872 28648 15608 28676
rect 15891 28648 15936 28676
rect 13872 28636 13878 28648
rect 15930 28636 15936 28648
rect 15988 28636 15994 28688
rect 17788 28620 17816 28716
rect 18414 28704 18420 28716
rect 18472 28704 18478 28756
rect 19150 28744 19156 28756
rect 19111 28716 19156 28744
rect 19150 28704 19156 28716
rect 19208 28704 19214 28756
rect 21266 28704 21272 28756
rect 21324 28744 21330 28756
rect 21361 28747 21419 28753
rect 21361 28744 21373 28747
rect 21324 28716 21373 28744
rect 21324 28704 21330 28716
rect 21361 28713 21373 28716
rect 21407 28713 21419 28747
rect 22830 28744 22836 28756
rect 21361 28707 21419 28713
rect 22710 28716 22836 28744
rect 18046 28676 18052 28688
rect 18007 28648 18052 28676
rect 18046 28636 18052 28648
rect 18104 28676 18110 28688
rect 18693 28679 18751 28685
rect 18693 28676 18705 28679
rect 18104 28648 18705 28676
rect 18104 28636 18110 28648
rect 18693 28645 18705 28648
rect 18739 28645 18751 28679
rect 18693 28639 18751 28645
rect 14185 28611 14243 28617
rect 14185 28577 14197 28611
rect 14231 28608 14243 28611
rect 14231 28580 14412 28608
rect 14231 28577 14243 28580
rect 14185 28571 14243 28577
rect 14384 28552 14412 28580
rect 17218 28568 17224 28620
rect 17276 28608 17282 28620
rect 17313 28611 17371 28617
rect 17313 28608 17325 28611
rect 17276 28580 17325 28608
rect 17276 28568 17282 28580
rect 17313 28577 17325 28580
rect 17359 28577 17371 28611
rect 17770 28608 17776 28620
rect 17731 28580 17776 28608
rect 17313 28571 17371 28577
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 19153 28611 19211 28617
rect 19153 28577 19165 28611
rect 19199 28608 19211 28611
rect 19242 28608 19248 28620
rect 19199 28580 19248 28608
rect 19199 28577 19211 28580
rect 19153 28571 19211 28577
rect 19242 28568 19248 28580
rect 19300 28568 19306 28620
rect 19334 28568 19340 28620
rect 19392 28608 19398 28620
rect 19429 28611 19487 28617
rect 19429 28608 19441 28611
rect 19392 28580 19441 28608
rect 19392 28568 19398 28580
rect 19429 28577 19441 28580
rect 19475 28608 19487 28611
rect 20898 28608 20904 28620
rect 19475 28580 20024 28608
rect 20859 28580 20904 28608
rect 19475 28577 19487 28580
rect 19429 28571 19487 28577
rect 14366 28500 14372 28552
rect 14424 28500 14430 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 15838 28540 15844 28552
rect 15528 28512 15844 28540
rect 15528 28500 15534 28512
rect 15838 28500 15844 28512
rect 15896 28500 15902 28552
rect 16482 28540 16488 28552
rect 16443 28512 16488 28540
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 14369 28407 14427 28413
rect 14369 28373 14381 28407
rect 14415 28404 14427 28407
rect 17218 28404 17224 28416
rect 14415 28376 17224 28404
rect 14415 28373 14427 28376
rect 14369 28367 14427 28373
rect 17218 28364 17224 28376
rect 17276 28364 17282 28416
rect 19996 28413 20024 28580
rect 20898 28568 20904 28580
rect 20956 28568 20962 28620
rect 22557 28611 22615 28617
rect 22557 28577 22569 28611
rect 22603 28608 22615 28611
rect 22710 28608 22738 28716
rect 22830 28704 22836 28716
rect 22888 28704 22894 28756
rect 24210 28704 24216 28756
rect 24268 28744 24274 28756
rect 25866 28744 25872 28756
rect 24268 28716 25872 28744
rect 24268 28704 24274 28716
rect 25866 28704 25872 28716
rect 25924 28704 25930 28756
rect 26234 28704 26240 28756
rect 26292 28744 26298 28756
rect 26651 28747 26709 28753
rect 26651 28744 26663 28747
rect 26292 28716 26663 28744
rect 26292 28704 26298 28716
rect 26651 28713 26663 28716
rect 26697 28713 26709 28747
rect 28258 28744 28264 28756
rect 28219 28716 28264 28744
rect 26651 28707 26709 28713
rect 28258 28704 28264 28716
rect 28316 28704 28322 28756
rect 29365 28747 29423 28753
rect 29365 28713 29377 28747
rect 29411 28744 29423 28747
rect 29454 28744 29460 28756
rect 29411 28716 29460 28744
rect 29411 28713 29423 28716
rect 29365 28707 29423 28713
rect 29454 28704 29460 28716
rect 29512 28704 29518 28756
rect 30006 28704 30012 28756
rect 30064 28744 30070 28756
rect 30193 28747 30251 28753
rect 30193 28744 30205 28747
rect 30064 28716 30205 28744
rect 30064 28704 30070 28716
rect 30193 28713 30205 28716
rect 30239 28713 30251 28747
rect 32214 28744 32220 28756
rect 32175 28716 32220 28744
rect 30193 28707 30251 28713
rect 32214 28704 32220 28716
rect 32272 28704 32278 28756
rect 33321 28747 33379 28753
rect 33321 28713 33333 28747
rect 33367 28744 33379 28747
rect 33502 28744 33508 28756
rect 33367 28716 33508 28744
rect 33367 28713 33379 28716
rect 33321 28707 33379 28713
rect 33502 28704 33508 28716
rect 33560 28704 33566 28756
rect 34241 28747 34299 28753
rect 34241 28713 34253 28747
rect 34287 28744 34299 28747
rect 34514 28744 34520 28756
rect 34287 28716 34520 28744
rect 34287 28713 34299 28716
rect 34241 28707 34299 28713
rect 34514 28704 34520 28716
rect 34572 28704 34578 28756
rect 35342 28744 35348 28756
rect 35303 28716 35348 28744
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 36633 28747 36691 28753
rect 36633 28713 36645 28747
rect 36679 28744 36691 28747
rect 37642 28744 37648 28756
rect 36679 28716 37648 28744
rect 36679 28713 36691 28716
rect 36633 28707 36691 28713
rect 37642 28704 37648 28716
rect 37700 28704 37706 28756
rect 37921 28747 37979 28753
rect 37921 28713 37933 28747
rect 37967 28744 37979 28747
rect 38286 28744 38292 28756
rect 37967 28716 38292 28744
rect 37967 28713 37979 28716
rect 37921 28707 37979 28713
rect 38286 28704 38292 28716
rect 38344 28704 38350 28756
rect 38378 28704 38384 28756
rect 38436 28744 38442 28756
rect 38749 28747 38807 28753
rect 38749 28744 38761 28747
rect 38436 28716 38761 28744
rect 38436 28704 38442 28716
rect 38749 28713 38761 28716
rect 38795 28713 38807 28747
rect 38749 28707 38807 28713
rect 38930 28704 38936 28756
rect 38988 28744 38994 28756
rect 40218 28744 40224 28756
rect 38988 28716 40224 28744
rect 38988 28704 38994 28716
rect 40218 28704 40224 28716
rect 40276 28704 40282 28756
rect 41506 28744 41512 28756
rect 41467 28716 41512 28744
rect 41506 28704 41512 28716
rect 41564 28704 41570 28756
rect 42334 28704 42340 28756
rect 42392 28744 42398 28756
rect 42613 28747 42671 28753
rect 42613 28744 42625 28747
rect 42392 28716 42625 28744
rect 42392 28704 42398 28716
rect 42613 28713 42625 28716
rect 42659 28713 42671 28747
rect 44542 28744 44548 28756
rect 44503 28716 44548 28744
rect 42613 28707 42671 28713
rect 44542 28704 44548 28716
rect 44600 28704 44606 28756
rect 44818 28704 44824 28756
rect 44876 28744 44882 28756
rect 45005 28747 45063 28753
rect 45005 28744 45017 28747
rect 44876 28716 45017 28744
rect 44876 28704 44882 28716
rect 45005 28713 45017 28716
rect 45051 28713 45063 28747
rect 45005 28707 45063 28713
rect 24851 28679 24909 28685
rect 24851 28645 24863 28679
rect 24897 28676 24909 28679
rect 26142 28676 26148 28688
rect 24897 28648 26148 28676
rect 24897 28645 24909 28648
rect 24851 28639 24909 28645
rect 26142 28636 26148 28648
rect 26200 28636 26206 28688
rect 30098 28676 30104 28688
rect 30011 28648 30104 28676
rect 22603 28580 22738 28608
rect 22833 28611 22891 28617
rect 22603 28577 22615 28580
rect 22557 28571 22615 28577
rect 22833 28577 22845 28611
rect 22879 28608 22891 28611
rect 23474 28608 23480 28620
rect 22879 28580 23480 28608
rect 22879 28577 22891 28580
rect 22833 28571 22891 28577
rect 23474 28568 23480 28580
rect 23532 28608 23538 28620
rect 26580 28611 26638 28617
rect 23532 28580 24348 28608
rect 23532 28568 23538 28580
rect 22738 28540 22744 28552
rect 22699 28512 22744 28540
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 24320 28484 24348 28580
rect 26580 28577 26592 28611
rect 26626 28608 26638 28611
rect 26694 28608 26700 28620
rect 26626 28580 26700 28608
rect 26626 28577 26638 28580
rect 26580 28571 26638 28577
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 26970 28568 26976 28620
rect 27028 28608 27034 28620
rect 28166 28608 28172 28620
rect 27028 28580 28172 28608
rect 27028 28568 27034 28580
rect 28166 28568 28172 28580
rect 28224 28568 28230 28620
rect 28350 28568 28356 28620
rect 28408 28608 28414 28620
rect 28629 28611 28687 28617
rect 28629 28608 28641 28611
rect 28408 28580 28641 28608
rect 28408 28568 28414 28580
rect 28629 28577 28641 28580
rect 28675 28577 28687 28611
rect 28629 28571 28687 28577
rect 29362 28568 29368 28620
rect 29420 28608 29426 28620
rect 30024 28617 30052 28648
rect 30098 28636 30104 28648
rect 30156 28676 30162 28688
rect 32030 28676 32036 28688
rect 30156 28648 32036 28676
rect 30156 28636 30162 28648
rect 32030 28636 32036 28648
rect 32088 28636 32094 28688
rect 33686 28676 33692 28688
rect 33599 28648 33692 28676
rect 33686 28636 33692 28648
rect 33744 28676 33750 28688
rect 37660 28676 37688 28704
rect 39758 28676 39764 28688
rect 33744 28648 34523 28676
rect 37660 28648 39068 28676
rect 39719 28648 39764 28676
rect 33744 28636 33750 28648
rect 29641 28611 29699 28617
rect 29641 28608 29653 28611
rect 29420 28580 29653 28608
rect 29420 28568 29426 28580
rect 29641 28577 29653 28580
rect 29687 28577 29699 28611
rect 29641 28571 29699 28577
rect 30009 28611 30067 28617
rect 30009 28577 30021 28611
rect 30055 28577 30067 28611
rect 31018 28608 31024 28620
rect 30931 28580 31024 28608
rect 30009 28571 30067 28577
rect 31018 28568 31024 28580
rect 31076 28608 31082 28620
rect 31386 28608 31392 28620
rect 31076 28580 31392 28608
rect 31076 28568 31082 28580
rect 31386 28568 31392 28580
rect 31444 28568 31450 28620
rect 32401 28611 32459 28617
rect 32401 28577 32413 28611
rect 32447 28608 32459 28611
rect 32490 28608 32496 28620
rect 32447 28580 32496 28608
rect 32447 28577 32459 28580
rect 32401 28571 32459 28577
rect 32490 28568 32496 28580
rect 32548 28568 32554 28620
rect 32674 28608 32680 28620
rect 32635 28580 32680 28608
rect 32674 28568 32680 28580
rect 32732 28568 32738 28620
rect 34330 28608 34336 28620
rect 34291 28580 34336 28608
rect 34330 28568 34336 28580
rect 34388 28568 34394 28620
rect 34495 28617 34523 28648
rect 34480 28611 34538 28617
rect 34480 28577 34492 28611
rect 34526 28608 34538 28611
rect 35250 28608 35256 28620
rect 34526 28580 35256 28608
rect 34526 28577 34538 28580
rect 34480 28571 34538 28577
rect 35250 28568 35256 28580
rect 35308 28568 35314 28620
rect 36078 28608 36084 28620
rect 36039 28580 36084 28608
rect 36078 28568 36084 28580
rect 36136 28568 36142 28620
rect 36449 28611 36507 28617
rect 36449 28577 36461 28611
rect 36495 28608 36507 28611
rect 37090 28608 37096 28620
rect 36495 28580 37096 28608
rect 36495 28577 36507 28580
rect 36449 28571 36507 28577
rect 37090 28568 37096 28580
rect 37148 28568 37154 28620
rect 37734 28608 37740 28620
rect 37695 28580 37740 28608
rect 37734 28568 37740 28580
rect 37792 28568 37798 28620
rect 39040 28617 39068 28648
rect 39758 28636 39764 28648
rect 39816 28636 39822 28688
rect 41414 28636 41420 28688
rect 41472 28676 41478 28688
rect 41785 28679 41843 28685
rect 41785 28676 41797 28679
rect 41472 28648 41797 28676
rect 41472 28636 41478 28648
rect 41785 28645 41797 28648
rect 41831 28676 41843 28679
rect 42058 28676 42064 28688
rect 41831 28648 42064 28676
rect 41831 28645 41843 28648
rect 41785 28639 41843 28645
rect 42058 28636 42064 28648
rect 42116 28636 42122 28688
rect 39025 28611 39083 28617
rect 39025 28577 39037 28611
rect 39071 28608 39083 28611
rect 39298 28608 39304 28620
rect 39071 28580 39304 28608
rect 39071 28577 39083 28580
rect 39025 28571 39083 28577
rect 39298 28568 39304 28580
rect 39356 28568 39362 28620
rect 39574 28608 39580 28620
rect 39535 28580 39580 28608
rect 39574 28568 39580 28580
rect 39632 28568 39638 28620
rect 40586 28608 40592 28620
rect 40547 28580 40592 28608
rect 40586 28568 40592 28580
rect 40644 28568 40650 28620
rect 42337 28611 42395 28617
rect 42337 28577 42349 28611
rect 42383 28608 42395 28611
rect 43070 28608 43076 28620
rect 42383 28580 43076 28608
rect 42383 28577 42395 28580
rect 42337 28571 42395 28577
rect 43070 28568 43076 28580
rect 43128 28608 43134 28620
rect 43384 28611 43442 28617
rect 43384 28608 43396 28611
rect 43128 28580 43396 28608
rect 43128 28568 43134 28580
rect 43384 28577 43396 28580
rect 43430 28577 43442 28611
rect 43384 28571 43442 28577
rect 45624 28611 45682 28617
rect 45624 28577 45636 28611
rect 45670 28608 45682 28611
rect 45738 28608 45744 28620
rect 45670 28580 45744 28608
rect 45670 28577 45682 28580
rect 45624 28571 45682 28577
rect 45738 28568 45744 28580
rect 45796 28568 45802 28620
rect 46569 28611 46627 28617
rect 46569 28577 46581 28611
rect 46615 28608 46627 28611
rect 47118 28608 47124 28620
rect 46615 28580 47124 28608
rect 46615 28577 46627 28580
rect 46569 28571 46627 28577
rect 47118 28568 47124 28580
rect 47176 28568 47182 28620
rect 24486 28540 24492 28552
rect 24447 28512 24492 28540
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 30466 28500 30472 28552
rect 30524 28540 30530 28552
rect 30561 28543 30619 28549
rect 30561 28540 30573 28543
rect 30524 28512 30573 28540
rect 30524 28500 30530 28512
rect 30561 28509 30573 28512
rect 30607 28540 30619 28543
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 30607 28512 31585 28540
rect 30607 28509 30619 28512
rect 30561 28503 30619 28509
rect 31573 28509 31585 28512
rect 31619 28540 31631 28543
rect 31662 28540 31668 28552
rect 31619 28512 31668 28540
rect 31619 28509 31631 28512
rect 31573 28503 31631 28509
rect 31662 28500 31668 28512
rect 31720 28540 31726 28552
rect 32692 28540 32720 28568
rect 31720 28512 32720 28540
rect 31720 28500 31726 28512
rect 34054 28500 34060 28552
rect 34112 28540 34118 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34112 28512 34713 28540
rect 34112 28500 34118 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 41693 28543 41751 28549
rect 41693 28509 41705 28543
rect 41739 28540 41751 28543
rect 41782 28540 41788 28552
rect 41739 28512 41788 28540
rect 41739 28509 41751 28512
rect 41693 28503 41751 28509
rect 41782 28500 41788 28512
rect 41840 28500 41846 28552
rect 23198 28432 23204 28484
rect 23256 28472 23262 28484
rect 24210 28472 24216 28484
rect 23256 28444 24216 28472
rect 23256 28432 23262 28444
rect 24210 28432 24216 28444
rect 24268 28432 24274 28484
rect 24302 28432 24308 28484
rect 24360 28472 24366 28484
rect 31205 28475 31263 28481
rect 31205 28472 31217 28475
rect 24360 28444 31217 28472
rect 24360 28432 24366 28444
rect 31205 28441 31217 28444
rect 31251 28441 31263 28475
rect 34606 28472 34612 28484
rect 34567 28444 34612 28472
rect 31205 28435 31263 28441
rect 34606 28432 34612 28444
rect 34664 28432 34670 28484
rect 19981 28407 20039 28413
rect 19981 28373 19993 28407
rect 20027 28404 20039 28407
rect 21082 28404 21088 28416
rect 20027 28376 21088 28404
rect 20027 28373 20039 28376
rect 19981 28367 20039 28373
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 21450 28364 21456 28416
rect 21508 28404 21514 28416
rect 21821 28407 21879 28413
rect 21821 28404 21833 28407
rect 21508 28376 21833 28404
rect 21508 28364 21514 28376
rect 21821 28373 21833 28376
rect 21867 28373 21879 28407
rect 25406 28404 25412 28416
rect 25367 28376 25412 28404
rect 21821 28367 21879 28373
rect 25406 28364 25412 28376
rect 25464 28364 25470 28416
rect 34698 28364 34704 28416
rect 34756 28404 34762 28416
rect 34793 28407 34851 28413
rect 34793 28404 34805 28407
rect 34756 28376 34805 28404
rect 34756 28364 34762 28376
rect 34793 28373 34805 28376
rect 34839 28373 34851 28407
rect 38470 28404 38476 28416
rect 38431 28376 38476 28404
rect 34793 28367 34851 28373
rect 38470 28364 38476 28376
rect 38528 28364 38534 28416
rect 40727 28407 40785 28413
rect 40727 28373 40739 28407
rect 40773 28404 40785 28407
rect 40954 28404 40960 28416
rect 40773 28376 40960 28404
rect 40773 28373 40785 28376
rect 40727 28367 40785 28373
rect 40954 28364 40960 28376
rect 41012 28364 41018 28416
rect 41138 28404 41144 28416
rect 41099 28376 41144 28404
rect 41138 28364 41144 28376
rect 41196 28364 41202 28416
rect 43162 28364 43168 28416
rect 43220 28404 43226 28416
rect 43487 28407 43545 28413
rect 43487 28404 43499 28407
rect 43220 28376 43499 28404
rect 43220 28364 43226 28376
rect 43487 28373 43499 28376
rect 43533 28373 43545 28407
rect 45370 28404 45376 28416
rect 45331 28376 45376 28404
rect 43487 28367 43545 28373
rect 45370 28364 45376 28376
rect 45428 28364 45434 28416
rect 45695 28407 45753 28413
rect 45695 28373 45707 28407
rect 45741 28404 45753 28407
rect 46109 28407 46167 28413
rect 46109 28404 46121 28407
rect 45741 28376 46121 28404
rect 45741 28373 45753 28376
rect 45695 28367 45753 28373
rect 46109 28373 46121 28376
rect 46155 28404 46167 28407
rect 46198 28404 46204 28416
rect 46155 28376 46204 28404
rect 46155 28373 46167 28376
rect 46109 28367 46167 28373
rect 46198 28364 46204 28376
rect 46256 28364 46262 28416
rect 46750 28404 46756 28416
rect 46711 28376 46756 28404
rect 46750 28364 46756 28376
rect 46808 28364 46814 28416
rect 47121 28407 47179 28413
rect 47121 28373 47133 28407
rect 47167 28404 47179 28407
rect 47210 28404 47216 28416
rect 47167 28376 47216 28404
rect 47167 28373 47179 28376
rect 47121 28367 47179 28373
rect 47210 28364 47216 28376
rect 47268 28404 47274 28416
rect 48222 28404 48228 28416
rect 47268 28376 48228 28404
rect 47268 28364 47274 28376
rect 48222 28364 48228 28376
rect 48280 28364 48286 28416
rect 1104 28314 48852 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 48852 28314
rect 1104 28240 48852 28262
rect 14093 28203 14151 28209
rect 14093 28169 14105 28203
rect 14139 28200 14151 28203
rect 14366 28200 14372 28212
rect 14139 28172 14372 28200
rect 14139 28169 14151 28172
rect 14093 28163 14151 28169
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 15470 28200 15476 28212
rect 15431 28172 15476 28200
rect 15470 28160 15476 28172
rect 15528 28160 15534 28212
rect 15841 28203 15899 28209
rect 15841 28169 15853 28203
rect 15887 28200 15899 28203
rect 15930 28200 15936 28212
rect 15887 28172 15936 28200
rect 15887 28169 15899 28172
rect 15841 28163 15899 28169
rect 15930 28160 15936 28172
rect 15988 28160 15994 28212
rect 17770 28200 17776 28212
rect 17731 28172 17776 28200
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 18601 28203 18659 28209
rect 18601 28169 18613 28203
rect 18647 28200 18659 28203
rect 19334 28200 19340 28212
rect 18647 28172 19340 28200
rect 18647 28169 18659 28172
rect 18601 28163 18659 28169
rect 14200 28036 18000 28064
rect 13630 27996 13636 28008
rect 13543 27968 13636 27996
rect 13630 27956 13636 27968
rect 13688 27996 13694 28008
rect 14200 28005 14228 28036
rect 14185 27999 14243 28005
rect 14185 27996 14197 27999
rect 13688 27968 14197 27996
rect 13688 27956 13694 27968
rect 14185 27965 14197 27968
rect 14231 27965 14243 27999
rect 14185 27959 14243 27965
rect 14645 27999 14703 28005
rect 14645 27965 14657 27999
rect 14691 27965 14703 27999
rect 14645 27959 14703 27965
rect 16301 27999 16359 28005
rect 16301 27965 16313 27999
rect 16347 27996 16359 27999
rect 16666 27996 16672 28008
rect 16347 27968 16672 27996
rect 16347 27965 16359 27968
rect 16301 27959 16359 27965
rect 13357 27931 13415 27937
rect 13357 27897 13369 27931
rect 13403 27928 13415 27931
rect 13722 27928 13728 27940
rect 13403 27900 13728 27928
rect 13403 27897 13415 27900
rect 13357 27891 13415 27897
rect 13722 27888 13728 27900
rect 13780 27928 13786 27940
rect 14660 27928 14688 27959
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 16945 27999 17003 28005
rect 16945 27965 16957 27999
rect 16991 27996 17003 27999
rect 17494 27996 17500 28008
rect 16991 27968 17500 27996
rect 16991 27965 17003 27968
rect 16945 27959 17003 27965
rect 17494 27956 17500 27968
rect 17552 27956 17558 28008
rect 17126 27928 17132 27940
rect 13780 27900 14688 27928
rect 17087 27900 17132 27928
rect 13780 27888 13786 27900
rect 17126 27888 17132 27900
rect 17184 27888 17190 27940
rect 17972 27928 18000 28036
rect 18049 27999 18107 28005
rect 18049 27965 18061 27999
rect 18095 27996 18107 27999
rect 18616 27996 18644 28163
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 20898 28200 20904 28212
rect 20859 28172 20904 28200
rect 20898 28160 20904 28172
rect 20956 28160 20962 28212
rect 22830 28200 22836 28212
rect 22791 28172 22836 28200
rect 22830 28160 22836 28172
rect 22888 28160 22894 28212
rect 28166 28160 28172 28212
rect 28224 28200 28230 28212
rect 28997 28203 29055 28209
rect 28997 28200 29009 28203
rect 28224 28172 29009 28200
rect 28224 28160 28230 28172
rect 28997 28169 29009 28172
rect 29043 28169 29055 28203
rect 30098 28200 30104 28212
rect 30059 28172 30104 28200
rect 28997 28163 29055 28169
rect 30098 28160 30104 28172
rect 30156 28160 30162 28212
rect 31018 28200 31024 28212
rect 30979 28172 31024 28200
rect 31018 28160 31024 28172
rect 31076 28160 31082 28212
rect 31389 28203 31447 28209
rect 31389 28169 31401 28203
rect 31435 28200 31447 28203
rect 31846 28200 31852 28212
rect 31435 28172 31852 28200
rect 31435 28169 31447 28172
rect 31389 28163 31447 28169
rect 31846 28160 31852 28172
rect 31904 28200 31910 28212
rect 32398 28200 32404 28212
rect 31904 28172 32404 28200
rect 31904 28160 31910 28172
rect 32398 28160 32404 28172
rect 32456 28160 32462 28212
rect 32674 28160 32680 28212
rect 32732 28200 32738 28212
rect 33413 28203 33471 28209
rect 33413 28200 33425 28203
rect 32732 28172 33425 28200
rect 32732 28160 32738 28172
rect 33413 28169 33425 28172
rect 33459 28169 33471 28203
rect 34054 28200 34060 28212
rect 34015 28172 34060 28200
rect 33413 28163 33471 28169
rect 34054 28160 34060 28172
rect 34112 28160 34118 28212
rect 34425 28203 34483 28209
rect 34425 28169 34437 28203
rect 34471 28200 34483 28203
rect 34606 28200 34612 28212
rect 34471 28172 34612 28200
rect 34471 28169 34483 28172
rect 34425 28163 34483 28169
rect 34606 28160 34612 28172
rect 34664 28160 34670 28212
rect 35069 28203 35127 28209
rect 35069 28169 35081 28203
rect 35115 28200 35127 28203
rect 35250 28200 35256 28212
rect 35115 28172 35256 28200
rect 35115 28169 35127 28172
rect 35069 28163 35127 28169
rect 35250 28160 35256 28172
rect 35308 28160 35314 28212
rect 36173 28203 36231 28209
rect 36173 28169 36185 28203
rect 36219 28200 36231 28203
rect 36354 28200 36360 28212
rect 36219 28172 36360 28200
rect 36219 28169 36231 28172
rect 36173 28163 36231 28169
rect 36354 28160 36360 28172
rect 36412 28160 36418 28212
rect 37182 28160 37188 28212
rect 37240 28200 37246 28212
rect 37461 28203 37519 28209
rect 37461 28200 37473 28203
rect 37240 28172 37473 28200
rect 37240 28160 37246 28172
rect 37461 28169 37473 28172
rect 37507 28169 37519 28203
rect 37461 28163 37519 28169
rect 39298 28160 39304 28212
rect 39356 28200 39362 28212
rect 39393 28203 39451 28209
rect 39393 28200 39405 28203
rect 39356 28172 39405 28200
rect 39356 28160 39362 28172
rect 39393 28169 39405 28172
rect 39439 28169 39451 28203
rect 39393 28163 39451 28169
rect 39574 28160 39580 28212
rect 39632 28200 39638 28212
rect 39761 28203 39819 28209
rect 39761 28200 39773 28203
rect 39632 28172 39773 28200
rect 39632 28160 39638 28172
rect 39761 28169 39773 28172
rect 39807 28169 39819 28203
rect 39761 28163 39819 28169
rect 40218 28160 40224 28212
rect 40276 28200 40282 28212
rect 40586 28200 40592 28212
rect 40276 28172 40592 28200
rect 40276 28160 40282 28172
rect 40586 28160 40592 28172
rect 40644 28200 40650 28212
rect 40681 28203 40739 28209
rect 40681 28200 40693 28203
rect 40644 28172 40693 28200
rect 40644 28160 40650 28172
rect 40681 28169 40693 28172
rect 40727 28169 40739 28203
rect 42058 28200 42064 28212
rect 42019 28172 42064 28200
rect 40681 28163 40739 28169
rect 42058 28160 42064 28172
rect 42116 28160 42122 28212
rect 43070 28160 43076 28212
rect 43128 28200 43134 28212
rect 43441 28203 43499 28209
rect 43441 28200 43453 28203
rect 43128 28172 43453 28200
rect 43128 28160 43134 28172
rect 43441 28169 43453 28172
rect 43487 28169 43499 28203
rect 43441 28163 43499 28169
rect 44223 28203 44281 28209
rect 44223 28169 44235 28203
rect 44269 28200 44281 28203
rect 45370 28200 45376 28212
rect 44269 28172 45376 28200
rect 44269 28169 44281 28172
rect 44223 28163 44281 28169
rect 45370 28160 45376 28172
rect 45428 28160 45434 28212
rect 18969 28135 19027 28141
rect 18969 28101 18981 28135
rect 19015 28132 19027 28135
rect 19242 28132 19248 28144
rect 19015 28104 19248 28132
rect 19015 28101 19027 28104
rect 18969 28095 19027 28101
rect 19242 28092 19248 28104
rect 19300 28092 19306 28144
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28064 19855 28067
rect 22848 28064 22876 28160
rect 28258 28092 28264 28144
rect 28316 28132 28322 28144
rect 30653 28135 30711 28141
rect 30653 28132 30665 28135
rect 28316 28104 30665 28132
rect 28316 28092 28322 28104
rect 30653 28101 30665 28104
rect 30699 28101 30711 28135
rect 30653 28095 30711 28101
rect 33137 28135 33195 28141
rect 33137 28101 33149 28135
rect 33183 28132 33195 28135
rect 33318 28132 33324 28144
rect 33183 28104 33324 28132
rect 33183 28101 33195 28104
rect 33137 28095 33195 28101
rect 33318 28092 33324 28104
rect 33376 28092 33382 28144
rect 36449 28135 36507 28141
rect 36449 28101 36461 28135
rect 36495 28132 36507 28135
rect 39482 28132 39488 28144
rect 36495 28104 39488 28132
rect 36495 28101 36507 28104
rect 36449 28095 36507 28101
rect 39482 28092 39488 28104
rect 39540 28092 39546 28144
rect 41874 28092 41880 28144
rect 41932 28132 41938 28144
rect 42429 28135 42487 28141
rect 42429 28132 42441 28135
rect 41932 28104 42441 28132
rect 41932 28092 41938 28104
rect 42429 28101 42441 28104
rect 42475 28101 42487 28135
rect 42429 28095 42487 28101
rect 24486 28064 24492 28076
rect 19843 28036 22876 28064
rect 24399 28036 24492 28064
rect 19843 28033 19855 28036
rect 19797 28027 19855 28033
rect 20180 28005 20208 28036
rect 24486 28024 24492 28036
rect 24544 28064 24550 28076
rect 25133 28067 25191 28073
rect 25133 28064 25145 28067
rect 24544 28036 25145 28064
rect 24544 28024 24550 28036
rect 25133 28033 25145 28036
rect 25179 28033 25191 28067
rect 25133 28027 25191 28033
rect 26050 28024 26056 28076
rect 26108 28064 26114 28076
rect 26326 28064 26332 28076
rect 26108 28036 26332 28064
rect 26108 28024 26114 28036
rect 26326 28024 26332 28036
rect 26384 28064 26390 28076
rect 28077 28067 28135 28073
rect 26384 28036 26601 28064
rect 26384 28024 26390 28036
rect 18095 27968 18644 27996
rect 20165 27999 20223 28005
rect 18095 27965 18107 27968
rect 18049 27959 18107 27965
rect 20165 27965 20177 27999
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27996 20499 27999
rect 21082 27996 21088 28008
rect 20487 27968 21088 27996
rect 20487 27965 20499 27968
rect 20441 27959 20499 27965
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 21637 27999 21695 28005
rect 21637 27996 21649 27999
rect 21192 27968 21649 27996
rect 21192 27928 21220 27968
rect 21637 27965 21649 27968
rect 21683 27996 21695 27999
rect 21818 27996 21824 28008
rect 21683 27968 21824 27996
rect 21683 27965 21695 27968
rect 21637 27959 21695 27965
rect 21818 27956 21824 27968
rect 21876 27956 21882 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 22646 27996 22652 28008
rect 22327 27968 22652 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 17972 27900 21220 27928
rect 21450 27888 21456 27940
rect 21508 27928 21514 27940
rect 22296 27928 22324 27959
rect 22646 27956 22652 27968
rect 22704 27956 22710 28008
rect 23474 27956 23480 28008
rect 23532 27996 23538 28008
rect 24029 27999 24087 28005
rect 24029 27996 24041 27999
rect 23532 27968 24041 27996
rect 23532 27956 23538 27968
rect 24029 27965 24041 27968
rect 24075 27996 24087 27999
rect 24118 27996 24124 28008
rect 24075 27968 24124 27996
rect 24075 27965 24087 27968
rect 24029 27959 24087 27965
rect 24118 27956 24124 27968
rect 24176 27956 24182 28008
rect 24302 27996 24308 28008
rect 24263 27968 24308 27996
rect 24302 27956 24308 27968
rect 24360 27956 24366 28008
rect 25682 27996 25688 28008
rect 25643 27968 25688 27996
rect 25682 27956 25688 27968
rect 25740 27956 25746 28008
rect 26573 27996 26601 28036
rect 28077 28033 28089 28067
rect 28123 28064 28135 28067
rect 28350 28064 28356 28076
rect 28123 28036 28356 28064
rect 28123 28033 28135 28036
rect 28077 28027 28135 28033
rect 28350 28024 28356 28036
rect 28408 28024 28414 28076
rect 31478 28064 31484 28076
rect 31439 28036 31484 28064
rect 31478 28024 31484 28036
rect 31536 28024 31542 28076
rect 39022 28064 39028 28076
rect 38626 28036 39028 28064
rect 28204 27999 28262 28005
rect 28204 27996 28216 27999
rect 26573 27968 28216 27996
rect 28204 27965 28216 27968
rect 28250 27996 28262 27999
rect 28629 27999 28687 28005
rect 28629 27996 28641 27999
rect 28250 27968 28641 27996
rect 28250 27965 28262 27968
rect 28204 27959 28262 27965
rect 28629 27965 28641 27968
rect 28675 27965 28687 27999
rect 28629 27959 28687 27965
rect 29178 27956 29184 28008
rect 29236 27996 29242 28008
rect 29308 27999 29366 28005
rect 29308 27996 29320 27999
rect 29236 27968 29320 27996
rect 29236 27956 29242 27968
rect 29308 27965 29320 27968
rect 29354 27996 29366 27999
rect 29733 27999 29791 28005
rect 29733 27996 29745 27999
rect 29354 27968 29745 27996
rect 29354 27965 29366 27968
rect 29308 27959 29366 27965
rect 29733 27965 29745 27968
rect 29779 27965 29791 27999
rect 30466 27996 30472 28008
rect 30427 27968 30472 27996
rect 29733 27959 29791 27965
rect 30466 27956 30472 27968
rect 30524 27956 30530 28008
rect 30834 27956 30840 28008
rect 30892 27996 30898 28008
rect 30892 27968 32076 27996
rect 30892 27956 30898 27968
rect 32048 27940 32076 27968
rect 33042 27956 33048 28008
rect 33100 27996 33106 28008
rect 33229 27999 33287 28005
rect 33229 27996 33241 27999
rect 33100 27968 33241 27996
rect 33100 27956 33106 27968
rect 33229 27965 33241 27968
rect 33275 27965 33287 27999
rect 35320 27999 35378 28005
rect 35320 27996 35332 27999
rect 33229 27959 33287 27965
rect 35303 27965 35332 27996
rect 35366 27996 35378 27999
rect 36265 27999 36323 28005
rect 35366 27968 35848 27996
rect 35366 27965 35378 27968
rect 35303 27959 35378 27965
rect 21508 27900 22324 27928
rect 24857 27931 24915 27937
rect 21508 27888 21514 27900
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25593 27931 25651 27937
rect 25593 27928 25605 27931
rect 24903 27900 25605 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25593 27897 25605 27900
rect 25639 27928 25651 27931
rect 26047 27931 26105 27937
rect 26047 27928 26059 27931
rect 25639 27900 26059 27928
rect 25639 27897 25651 27900
rect 25593 27891 25651 27897
rect 26047 27897 26059 27900
rect 26093 27928 26105 27931
rect 26142 27928 26148 27940
rect 26093 27900 26148 27928
rect 26093 27897 26105 27900
rect 26047 27891 26105 27897
rect 26142 27888 26148 27900
rect 26200 27888 26206 27940
rect 28307 27931 28365 27937
rect 28307 27897 28319 27931
rect 28353 27928 28365 27931
rect 30926 27928 30932 27940
rect 28353 27900 30932 27928
rect 28353 27897 28365 27900
rect 28307 27891 28365 27897
rect 30926 27888 30932 27900
rect 30984 27888 30990 27940
rect 31734 27931 31792 27937
rect 31734 27897 31746 27931
rect 31780 27928 31792 27931
rect 31846 27928 31852 27940
rect 31780 27900 31852 27928
rect 31780 27897 31792 27900
rect 31734 27891 31792 27897
rect 31846 27888 31852 27900
rect 31904 27888 31910 27940
rect 32030 27888 32036 27940
rect 32088 27928 32094 27940
rect 35303 27928 35331 27959
rect 32088 27900 35331 27928
rect 32088 27888 32094 27900
rect 14458 27860 14464 27872
rect 14419 27832 14464 27860
rect 14458 27820 14464 27832
rect 14516 27820 14522 27872
rect 17218 27820 17224 27872
rect 17276 27860 17282 27872
rect 17405 27863 17463 27869
rect 17405 27860 17417 27863
rect 17276 27832 17417 27860
rect 17276 27820 17282 27832
rect 17405 27829 17417 27832
rect 17451 27829 17463 27863
rect 18230 27860 18236 27872
rect 18191 27832 18236 27860
rect 17405 27823 17463 27829
rect 18230 27820 18236 27832
rect 18288 27820 18294 27872
rect 19978 27860 19984 27872
rect 19939 27832 19984 27860
rect 19978 27820 19984 27832
rect 20036 27820 20042 27872
rect 21910 27860 21916 27872
rect 21871 27832 21916 27860
rect 21910 27820 21916 27832
rect 21968 27820 21974 27872
rect 26602 27860 26608 27872
rect 26563 27832 26608 27860
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 26694 27820 26700 27872
rect 26752 27860 26758 27872
rect 26973 27863 27031 27869
rect 26973 27860 26985 27863
rect 26752 27832 26985 27860
rect 26752 27820 26758 27832
rect 26973 27829 26985 27832
rect 27019 27860 27031 27863
rect 28074 27860 28080 27872
rect 27019 27832 28080 27860
rect 27019 27829 27031 27832
rect 26973 27823 27031 27829
rect 28074 27820 28080 27832
rect 28132 27820 28138 27872
rect 29270 27820 29276 27872
rect 29328 27860 29334 27872
rect 29411 27863 29469 27869
rect 29411 27860 29423 27863
rect 29328 27832 29423 27860
rect 29328 27820 29334 27832
rect 29411 27829 29423 27832
rect 29457 27829 29469 27863
rect 29411 27823 29469 27829
rect 30558 27820 30564 27872
rect 30616 27860 30622 27872
rect 32401 27863 32459 27869
rect 32401 27860 32413 27863
rect 30616 27832 32413 27860
rect 30616 27820 30622 27832
rect 32401 27829 32413 27832
rect 32447 27829 32459 27863
rect 32401 27823 32459 27829
rect 32490 27820 32496 27872
rect 32548 27860 32554 27872
rect 32769 27863 32827 27869
rect 32769 27860 32781 27863
rect 32548 27832 32781 27860
rect 32548 27820 32554 27832
rect 32769 27829 32781 27832
rect 32815 27860 32827 27863
rect 32950 27860 32956 27872
rect 32815 27832 32956 27860
rect 32815 27829 32827 27832
rect 32769 27823 32827 27829
rect 32950 27820 32956 27832
rect 33008 27820 33014 27872
rect 35391 27863 35449 27869
rect 35391 27829 35403 27863
rect 35437 27860 35449 27863
rect 35618 27860 35624 27872
rect 35437 27832 35624 27860
rect 35437 27829 35449 27832
rect 35391 27823 35449 27829
rect 35618 27820 35624 27832
rect 35676 27820 35682 27872
rect 35820 27869 35848 27968
rect 36265 27965 36277 27999
rect 36311 27996 36323 27999
rect 36725 27999 36783 28005
rect 36725 27996 36737 27999
rect 36311 27968 36737 27996
rect 36311 27965 36323 27968
rect 36265 27959 36323 27965
rect 36725 27965 36737 27968
rect 36771 27996 36783 27999
rect 37182 27996 37188 28008
rect 36771 27968 37188 27996
rect 36771 27965 36783 27968
rect 36725 27959 36783 27965
rect 37182 27956 37188 27968
rect 37240 27956 37246 28008
rect 37277 27999 37335 28005
rect 37277 27965 37289 27999
rect 37323 27996 37335 27999
rect 37550 27996 37556 28008
rect 37323 27968 37556 27996
rect 37323 27965 37335 27968
rect 37277 27959 37335 27965
rect 37550 27956 37556 27968
rect 37608 27996 37614 28008
rect 38105 27999 38163 28005
rect 38105 27996 38117 27999
rect 37608 27968 38117 27996
rect 37608 27956 37614 27968
rect 38105 27965 38117 27968
rect 38151 27965 38163 27999
rect 38470 27996 38476 28008
rect 38431 27968 38476 27996
rect 38105 27959 38163 27965
rect 38470 27956 38476 27968
rect 38528 27996 38534 28008
rect 38626 27996 38654 28036
rect 39022 28024 39028 28036
rect 39080 28024 39086 28076
rect 39117 28067 39175 28073
rect 39117 28033 39129 28067
rect 39163 28064 39175 28067
rect 44358 28064 44364 28076
rect 39163 28036 44364 28064
rect 39163 28033 39175 28036
rect 39117 28027 39175 28033
rect 44358 28024 44364 28036
rect 44416 28024 44422 28076
rect 46198 28064 46204 28076
rect 46159 28036 46204 28064
rect 46198 28024 46204 28036
rect 46256 28024 46262 28076
rect 46474 28064 46480 28076
rect 46435 28036 46480 28064
rect 46474 28024 46480 28036
rect 46532 28024 46538 28076
rect 38528 27968 38654 27996
rect 38528 27956 38534 27968
rect 38746 27956 38752 28008
rect 38804 27996 38810 28008
rect 38933 27999 38991 28005
rect 38933 27996 38945 27999
rect 38804 27968 38945 27996
rect 38804 27956 38810 27968
rect 38933 27965 38945 27968
rect 38979 27996 38991 27999
rect 39390 27996 39396 28008
rect 38979 27968 39396 27996
rect 38979 27965 38991 27968
rect 38933 27959 38991 27965
rect 39390 27956 39396 27968
rect 39448 27956 39454 28008
rect 42648 27999 42706 28005
rect 42648 27996 42660 27999
rect 41867 27968 42660 27996
rect 41138 27928 41144 27940
rect 41099 27900 41144 27928
rect 41138 27888 41144 27900
rect 41196 27888 41202 27940
rect 41230 27888 41236 27940
rect 41288 27928 41294 27940
rect 41288 27900 41333 27928
rect 41288 27888 41294 27900
rect 35805 27863 35863 27869
rect 35805 27829 35817 27863
rect 35851 27860 35863 27863
rect 36170 27860 36176 27872
rect 35851 27832 36176 27860
rect 35851 27829 35863 27832
rect 35805 27823 35863 27829
rect 36170 27820 36176 27832
rect 36228 27820 36234 27872
rect 37090 27860 37096 27872
rect 37051 27832 37096 27860
rect 37090 27820 37096 27832
rect 37148 27820 37154 27872
rect 37734 27820 37740 27872
rect 37792 27860 37798 27872
rect 37829 27863 37887 27869
rect 37829 27860 37841 27863
rect 37792 27832 37841 27860
rect 37792 27820 37798 27832
rect 37829 27829 37841 27832
rect 37875 27860 37887 27863
rect 38838 27860 38844 27872
rect 37875 27832 38844 27860
rect 37875 27829 37887 27832
rect 37829 27823 37887 27829
rect 38838 27820 38844 27832
rect 38896 27820 38902 27872
rect 40034 27820 40040 27872
rect 40092 27860 40098 27872
rect 41867 27860 41895 27968
rect 42648 27965 42660 27968
rect 42694 27996 42706 27999
rect 43073 27999 43131 28005
rect 43073 27996 43085 27999
rect 42694 27968 43085 27996
rect 42694 27965 42706 27968
rect 42648 27959 42706 27965
rect 43073 27965 43085 27968
rect 43119 27965 43131 27999
rect 43073 27959 43131 27965
rect 44152 27999 44210 28005
rect 44152 27965 44164 27999
rect 44198 27996 44210 27999
rect 44450 27996 44456 28008
rect 44198 27968 44456 27996
rect 44198 27965 44210 27968
rect 44152 27959 44210 27965
rect 44450 27956 44456 27968
rect 44508 27996 44514 28008
rect 44634 27996 44640 28008
rect 44508 27968 44640 27996
rect 44508 27956 44514 27968
rect 44634 27956 44640 27968
rect 44692 27956 44698 28008
rect 41969 27931 42027 27937
rect 41969 27897 41981 27931
rect 42015 27928 42027 27931
rect 42058 27928 42064 27940
rect 42015 27900 42064 27928
rect 42015 27897 42027 27900
rect 41969 27891 42027 27897
rect 42058 27888 42064 27900
rect 42116 27928 42122 27940
rect 42116 27900 45876 27928
rect 42116 27888 42122 27900
rect 40092 27832 41895 27860
rect 40092 27820 40098 27832
rect 42518 27820 42524 27872
rect 42576 27860 42582 27872
rect 42751 27863 42809 27869
rect 42751 27860 42763 27863
rect 42576 27832 42763 27860
rect 42576 27820 42582 27832
rect 42751 27829 42763 27832
rect 42797 27829 42809 27863
rect 44634 27860 44640 27872
rect 44595 27832 44640 27860
rect 42751 27823 42809 27829
rect 44634 27820 44640 27832
rect 44692 27820 44698 27872
rect 45649 27863 45707 27869
rect 45649 27829 45661 27863
rect 45695 27860 45707 27863
rect 45738 27860 45744 27872
rect 45695 27832 45744 27860
rect 45695 27829 45707 27832
rect 45649 27823 45707 27829
rect 45738 27820 45744 27832
rect 45796 27820 45802 27872
rect 45848 27860 45876 27900
rect 46198 27888 46204 27940
rect 46256 27928 46262 27940
rect 46293 27931 46351 27937
rect 46293 27928 46305 27931
rect 46256 27900 46305 27928
rect 46256 27888 46262 27900
rect 46293 27897 46305 27900
rect 46339 27897 46351 27931
rect 46293 27891 46351 27897
rect 46474 27860 46480 27872
rect 45848 27832 46480 27860
rect 46474 27820 46480 27832
rect 46532 27820 46538 27872
rect 47118 27860 47124 27872
rect 47079 27832 47124 27860
rect 47118 27820 47124 27832
rect 47176 27820 47182 27872
rect 1104 27770 48852 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 48852 27770
rect 1104 27696 48852 27718
rect 15378 27656 15384 27668
rect 15339 27628 15384 27656
rect 15378 27616 15384 27628
rect 15436 27616 15442 27668
rect 16666 27616 16672 27668
rect 16724 27656 16730 27668
rect 22373 27659 22431 27665
rect 16724 27628 21036 27656
rect 16724 27616 16730 27628
rect 19334 27588 19340 27600
rect 19295 27560 19340 27588
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 14182 27520 14188 27532
rect 14143 27492 14188 27520
rect 14182 27480 14188 27492
rect 14240 27480 14246 27532
rect 14550 27480 14556 27532
rect 14608 27520 14614 27532
rect 15565 27523 15623 27529
rect 15565 27520 15577 27523
rect 14608 27492 15577 27520
rect 14608 27480 14614 27492
rect 15565 27489 15577 27492
rect 15611 27520 15623 27523
rect 15746 27520 15752 27532
rect 15611 27492 15752 27520
rect 15611 27489 15623 27492
rect 15565 27483 15623 27489
rect 15746 27480 15752 27492
rect 15804 27480 15810 27532
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27520 15899 27523
rect 17218 27520 17224 27532
rect 15887 27492 16436 27520
rect 17179 27492 17224 27520
rect 15887 27489 15899 27492
rect 15841 27483 15899 27489
rect 16408 27464 16436 27492
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 17494 27480 17500 27532
rect 17552 27520 17558 27532
rect 17589 27523 17647 27529
rect 17589 27520 17601 27523
rect 17552 27492 17601 27520
rect 17552 27480 17558 27492
rect 17589 27489 17601 27492
rect 17635 27520 17647 27523
rect 18230 27520 18236 27532
rect 17635 27492 18236 27520
rect 17635 27489 17647 27492
rect 17589 27483 17647 27489
rect 18230 27480 18236 27492
rect 18288 27480 18294 27532
rect 19061 27523 19119 27529
rect 19061 27489 19073 27523
rect 19107 27520 19119 27523
rect 19150 27520 19156 27532
rect 19107 27492 19156 27520
rect 19107 27489 19119 27492
rect 19061 27483 19119 27489
rect 19150 27480 19156 27492
rect 19208 27480 19214 27532
rect 21008 27529 21036 27628
rect 22373 27625 22385 27659
rect 22419 27656 22431 27659
rect 23845 27659 23903 27665
rect 23845 27656 23857 27659
rect 22419 27628 23857 27656
rect 22419 27625 22431 27628
rect 22373 27619 22431 27625
rect 23845 27625 23857 27628
rect 23891 27656 23903 27659
rect 24302 27656 24308 27668
rect 23891 27628 24308 27656
rect 23891 27625 23903 27628
rect 23845 27619 23903 27625
rect 24302 27616 24308 27628
rect 24360 27616 24366 27668
rect 26510 27616 26516 27668
rect 26568 27656 26574 27668
rect 26605 27659 26663 27665
rect 26605 27656 26617 27659
rect 26568 27628 26617 27656
rect 26568 27616 26574 27628
rect 26605 27625 26617 27628
rect 26651 27625 26663 27659
rect 26605 27619 26663 27625
rect 29270 27616 29276 27668
rect 29328 27656 29334 27668
rect 29365 27659 29423 27665
rect 29365 27656 29377 27659
rect 29328 27628 29377 27656
rect 29328 27616 29334 27628
rect 29365 27625 29377 27628
rect 29411 27625 29423 27659
rect 31478 27656 31484 27668
rect 31439 27628 31484 27656
rect 29365 27619 29423 27625
rect 31478 27616 31484 27628
rect 31536 27616 31542 27668
rect 31662 27616 31668 27668
rect 31720 27656 31726 27668
rect 31849 27659 31907 27665
rect 31849 27656 31861 27659
rect 31720 27628 31861 27656
rect 31720 27616 31726 27628
rect 31849 27625 31861 27628
rect 31895 27625 31907 27659
rect 32490 27656 32496 27668
rect 32451 27628 32496 27656
rect 31849 27619 31907 27625
rect 32490 27616 32496 27628
rect 32548 27616 32554 27668
rect 33042 27616 33048 27668
rect 33100 27656 33106 27668
rect 33321 27659 33379 27665
rect 33321 27656 33333 27659
rect 33100 27628 33333 27656
rect 33100 27616 33106 27628
rect 33321 27625 33333 27628
rect 33367 27625 33379 27659
rect 33321 27619 33379 27625
rect 34422 27616 34428 27668
rect 34480 27656 34486 27668
rect 34885 27659 34943 27665
rect 34885 27656 34897 27659
rect 34480 27628 34897 27656
rect 34480 27616 34486 27628
rect 34885 27625 34897 27628
rect 34931 27625 34943 27659
rect 38470 27656 38476 27668
rect 34885 27619 34943 27625
rect 35728 27628 38476 27656
rect 22919 27591 22977 27597
rect 22919 27557 22931 27591
rect 22965 27588 22977 27591
rect 23014 27588 23020 27600
rect 22965 27560 23020 27588
rect 22965 27557 22977 27560
rect 22919 27551 22977 27557
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 25593 27591 25651 27597
rect 25593 27557 25605 27591
rect 25639 27588 25651 27591
rect 25682 27588 25688 27600
rect 25639 27560 25688 27588
rect 25639 27557 25651 27560
rect 25593 27551 25651 27557
rect 25682 27548 25688 27560
rect 25740 27588 25746 27600
rect 25869 27591 25927 27597
rect 25869 27588 25881 27591
rect 25740 27560 25881 27588
rect 25740 27548 25746 27560
rect 25869 27557 25881 27560
rect 25915 27557 25927 27591
rect 25869 27551 25927 27557
rect 28531 27591 28589 27597
rect 28531 27557 28543 27591
rect 28577 27588 28589 27591
rect 28718 27588 28724 27600
rect 28577 27560 28724 27588
rect 28577 27557 28589 27560
rect 28531 27551 28589 27557
rect 28718 27548 28724 27560
rect 28776 27548 28782 27600
rect 30558 27588 30564 27600
rect 30519 27560 30564 27588
rect 30558 27548 30564 27560
rect 30616 27548 30622 27600
rect 35728 27588 35756 27628
rect 38470 27616 38476 27628
rect 38528 27616 38534 27668
rect 38746 27656 38752 27668
rect 38707 27628 38752 27656
rect 38746 27616 38752 27628
rect 38804 27616 38810 27668
rect 38930 27616 38936 27668
rect 38988 27656 38994 27668
rect 39482 27656 39488 27668
rect 38988 27628 39488 27656
rect 38988 27616 38994 27628
rect 39482 27616 39488 27628
rect 39540 27656 39546 27668
rect 39577 27659 39635 27665
rect 39577 27656 39589 27659
rect 39540 27628 39589 27656
rect 39540 27616 39546 27628
rect 39577 27625 39589 27628
rect 39623 27625 39635 27659
rect 39577 27619 39635 27625
rect 41141 27659 41199 27665
rect 41141 27625 41153 27659
rect 41187 27656 41199 27659
rect 41230 27656 41236 27668
rect 41187 27628 41236 27656
rect 41187 27625 41199 27628
rect 41141 27619 41199 27625
rect 41230 27616 41236 27628
rect 41288 27656 41294 27668
rect 41288 27628 41920 27656
rect 41288 27616 41294 27628
rect 34164 27560 35756 27588
rect 35805 27591 35863 27597
rect 34164 27532 34192 27560
rect 35805 27557 35817 27591
rect 35851 27588 35863 27591
rect 35894 27588 35900 27600
rect 35851 27560 35900 27588
rect 35851 27557 35863 27560
rect 35805 27551 35863 27557
rect 35894 27548 35900 27560
rect 35952 27548 35958 27600
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 21082 27520 21088 27532
rect 21039 27492 21088 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 21450 27520 21456 27532
rect 21411 27492 21456 27520
rect 21450 27480 21456 27492
rect 21508 27480 21514 27532
rect 22557 27523 22615 27529
rect 22557 27489 22569 27523
rect 22603 27520 22615 27523
rect 22738 27520 22744 27532
rect 22603 27492 22744 27520
rect 22603 27489 22615 27492
rect 22557 27483 22615 27489
rect 22738 27480 22744 27492
rect 22796 27480 22802 27532
rect 24854 27520 24860 27532
rect 24815 27492 24860 27520
rect 24854 27480 24860 27492
rect 24912 27480 24918 27532
rect 25317 27523 25375 27529
rect 25317 27489 25329 27523
rect 25363 27489 25375 27523
rect 25317 27483 25375 27489
rect 16390 27412 16396 27464
rect 16448 27452 16454 27464
rect 16485 27455 16543 27461
rect 16485 27452 16497 27455
rect 16448 27424 16497 27452
rect 16448 27412 16454 27424
rect 16485 27421 16497 27424
rect 16531 27452 16543 27455
rect 17512 27452 17540 27480
rect 16531 27424 17540 27452
rect 17773 27455 17831 27461
rect 16531 27421 16543 27424
rect 16485 27415 16543 27421
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 18046 27452 18052 27464
rect 17819 27424 18052 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 21726 27452 21732 27464
rect 21687 27424 21732 27452
rect 21726 27412 21732 27424
rect 21784 27412 21790 27464
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 22704 27424 24685 27452
rect 22704 27412 22710 27424
rect 24673 27421 24685 27424
rect 24719 27452 24731 27455
rect 25332 27452 25360 27483
rect 26418 27480 26424 27532
rect 26476 27520 26482 27532
rect 26513 27523 26571 27529
rect 26513 27520 26525 27523
rect 26476 27492 26525 27520
rect 26476 27480 26482 27492
rect 26513 27489 26525 27492
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 26973 27523 27031 27529
rect 26973 27489 26985 27523
rect 27019 27489 27031 27523
rect 26973 27483 27031 27489
rect 32125 27523 32183 27529
rect 32125 27489 32137 27523
rect 32171 27520 32183 27523
rect 32214 27520 32220 27532
rect 32171 27492 32220 27520
rect 32171 27489 32183 27492
rect 32125 27483 32183 27489
rect 25498 27452 25504 27464
rect 24719 27424 25504 27452
rect 24719 27421 24731 27424
rect 24673 27415 24731 27421
rect 25498 27412 25504 27424
rect 25556 27452 25562 27464
rect 26988 27452 27016 27483
rect 32214 27480 32220 27492
rect 32272 27480 32278 27532
rect 34146 27520 34152 27532
rect 34107 27492 34152 27520
rect 34146 27480 34152 27492
rect 34204 27480 34210 27532
rect 34330 27520 34336 27532
rect 34291 27492 34336 27520
rect 34330 27480 34336 27492
rect 34388 27480 34394 27532
rect 38102 27480 38108 27532
rect 38160 27520 38166 27532
rect 38197 27523 38255 27529
rect 38197 27520 38209 27523
rect 38160 27492 38209 27520
rect 38160 27480 38166 27492
rect 38197 27489 38209 27492
rect 38243 27520 38255 27523
rect 38764 27520 38792 27616
rect 40954 27548 40960 27600
rect 41012 27588 41018 27600
rect 41782 27588 41788 27600
rect 41012 27560 41788 27588
rect 41012 27548 41018 27560
rect 41782 27548 41788 27560
rect 41840 27548 41846 27600
rect 41892 27597 41920 27628
rect 43898 27616 43904 27668
rect 43956 27656 43962 27668
rect 43956 27628 46612 27656
rect 43956 27616 43962 27628
rect 41877 27591 41935 27597
rect 41877 27557 41889 27591
rect 41923 27588 41935 27591
rect 41966 27588 41972 27600
rect 41923 27560 41972 27588
rect 41923 27557 41935 27560
rect 41877 27551 41935 27557
rect 41966 27548 41972 27560
rect 42024 27548 42030 27600
rect 44450 27548 44456 27600
rect 44508 27588 44514 27600
rect 44866 27591 44924 27597
rect 44866 27588 44878 27591
rect 44508 27560 44878 27588
rect 44508 27548 44514 27560
rect 44866 27557 44878 27560
rect 44912 27557 44924 27591
rect 46198 27588 46204 27600
rect 46111 27560 46204 27588
rect 44866 27551 44924 27557
rect 38243 27492 38792 27520
rect 38243 27489 38255 27492
rect 38197 27483 38255 27489
rect 43254 27480 43260 27532
rect 43312 27520 43318 27532
rect 43384 27523 43442 27529
rect 43384 27520 43396 27523
rect 43312 27492 43396 27520
rect 43312 27480 43318 27492
rect 43384 27489 43396 27492
rect 43430 27489 43442 27523
rect 43384 27483 43442 27489
rect 44358 27480 44364 27532
rect 44416 27520 44422 27532
rect 44545 27523 44603 27529
rect 44545 27520 44557 27523
rect 44416 27492 44557 27520
rect 44416 27480 44422 27492
rect 44545 27489 44557 27492
rect 44591 27489 44603 27523
rect 44545 27483 44603 27489
rect 25556 27424 27016 27452
rect 28169 27455 28227 27461
rect 25556 27412 25562 27424
rect 28169 27421 28181 27455
rect 28215 27452 28227 27455
rect 28350 27452 28356 27464
rect 28215 27424 28356 27452
rect 28215 27421 28227 27424
rect 28169 27415 28227 27421
rect 28350 27412 28356 27424
rect 28408 27412 28414 27464
rect 30466 27452 30472 27464
rect 30427 27424 30472 27452
rect 30466 27412 30472 27424
rect 30524 27412 30530 27464
rect 34422 27452 34428 27464
rect 34383 27424 34428 27452
rect 34422 27412 34428 27424
rect 34480 27412 34486 27464
rect 35710 27452 35716 27464
rect 35671 27424 35716 27452
rect 35710 27412 35716 27424
rect 35768 27412 35774 27464
rect 36354 27452 36360 27464
rect 36315 27424 36360 27452
rect 36354 27412 36360 27424
rect 36412 27412 36418 27464
rect 39209 27455 39267 27461
rect 39209 27421 39221 27455
rect 39255 27452 39267 27455
rect 39574 27452 39580 27464
rect 39255 27424 39580 27452
rect 39255 27421 39267 27424
rect 39209 27415 39267 27421
rect 39574 27412 39580 27424
rect 39632 27412 39638 27464
rect 42429 27455 42487 27461
rect 42429 27421 42441 27455
rect 42475 27452 42487 27455
rect 43714 27452 43720 27464
rect 42475 27424 43720 27452
rect 42475 27421 42487 27424
rect 42429 27415 42487 27421
rect 43714 27412 43720 27424
rect 43772 27412 43778 27464
rect 23842 27344 23848 27396
rect 23900 27384 23906 27396
rect 29178 27384 29184 27396
rect 23900 27356 29184 27384
rect 23900 27344 23906 27356
rect 29178 27344 29184 27356
rect 29236 27344 29242 27396
rect 31018 27384 31024 27396
rect 30979 27356 31024 27384
rect 31018 27344 31024 27356
rect 31076 27344 31082 27396
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 14366 27316 14372 27328
rect 13412 27288 14372 27316
rect 13412 27276 13418 27288
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 19886 27276 19892 27328
rect 19944 27316 19950 27328
rect 19981 27319 20039 27325
rect 19981 27316 19993 27319
rect 19944 27288 19993 27316
rect 19944 27276 19950 27288
rect 19981 27285 19993 27288
rect 20027 27285 20039 27319
rect 19981 27279 20039 27285
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 29086 27316 29092 27328
rect 23532 27288 23577 27316
rect 29047 27288 29092 27316
rect 23532 27276 23538 27288
rect 29086 27276 29092 27288
rect 29144 27276 29150 27328
rect 31110 27276 31116 27328
rect 31168 27316 31174 27328
rect 33045 27319 33103 27325
rect 33045 27316 33057 27319
rect 31168 27288 33057 27316
rect 31168 27276 31174 27288
rect 33045 27285 33057 27288
rect 33091 27285 33103 27319
rect 35250 27316 35256 27328
rect 35211 27288 35256 27316
rect 33045 27279 33103 27285
rect 35250 27276 35256 27288
rect 35308 27276 35314 27328
rect 36722 27316 36728 27328
rect 36683 27288 36728 27316
rect 36722 27276 36728 27288
rect 36780 27276 36786 27328
rect 38381 27319 38439 27325
rect 38381 27285 38393 27319
rect 38427 27316 38439 27319
rect 39390 27316 39396 27328
rect 38427 27288 39396 27316
rect 38427 27285 38439 27288
rect 38381 27279 38439 27285
rect 39390 27276 39396 27288
rect 39448 27276 39454 27328
rect 40126 27316 40132 27328
rect 40087 27288 40132 27316
rect 40126 27276 40132 27288
rect 40184 27276 40190 27328
rect 40494 27316 40500 27328
rect 40455 27288 40500 27316
rect 40494 27276 40500 27288
rect 40552 27276 40558 27328
rect 43254 27276 43260 27328
rect 43312 27316 43318 27328
rect 43487 27319 43545 27325
rect 43487 27316 43499 27319
rect 43312 27288 43499 27316
rect 43312 27276 43318 27288
rect 43487 27285 43499 27288
rect 43533 27285 43545 27319
rect 43487 27279 43545 27285
rect 45465 27319 45523 27325
rect 45465 27285 45477 27319
rect 45511 27316 45523 27319
rect 45830 27316 45836 27328
rect 45511 27288 45836 27316
rect 45511 27285 45523 27288
rect 45465 27279 45523 27285
rect 45830 27276 45836 27288
rect 45888 27316 45894 27328
rect 46124 27325 46152 27560
rect 46198 27548 46204 27560
rect 46256 27588 46262 27600
rect 46477 27591 46535 27597
rect 46477 27588 46489 27591
rect 46256 27560 46489 27588
rect 46256 27548 46262 27560
rect 46477 27557 46489 27560
rect 46523 27557 46535 27591
rect 46584 27588 46612 27628
rect 47029 27591 47087 27597
rect 47029 27588 47041 27591
rect 46584 27560 47041 27588
rect 46477 27551 46535 27557
rect 47029 27557 47041 27560
rect 47075 27557 47087 27591
rect 47029 27551 47087 27557
rect 46382 27452 46388 27464
rect 46343 27424 46388 27452
rect 46382 27412 46388 27424
rect 46440 27412 46446 27464
rect 46109 27319 46167 27325
rect 46109 27316 46121 27319
rect 45888 27288 46121 27316
rect 45888 27276 45894 27288
rect 46109 27285 46121 27288
rect 46155 27285 46167 27319
rect 46109 27279 46167 27285
rect 1104 27226 48852 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 48852 27226
rect 1104 27152 48852 27174
rect 13722 27112 13728 27124
rect 13683 27084 13728 27112
rect 13722 27072 13728 27084
rect 13780 27112 13786 27124
rect 14734 27112 14740 27124
rect 13780 27084 14740 27112
rect 13780 27072 13786 27084
rect 14734 27072 14740 27084
rect 14792 27072 14798 27124
rect 17494 27112 17500 27124
rect 17455 27084 17500 27112
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 21082 27112 21088 27124
rect 21043 27084 21088 27112
rect 21082 27072 21088 27084
rect 21140 27072 21146 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 23385 27115 23443 27121
rect 23385 27112 23397 27115
rect 22796 27084 23397 27112
rect 22796 27072 22802 27084
rect 23385 27081 23397 27084
rect 23431 27081 23443 27115
rect 26418 27112 26424 27124
rect 26379 27084 26424 27112
rect 23385 27075 23443 27081
rect 26418 27072 26424 27084
rect 26476 27112 26482 27124
rect 26789 27115 26847 27121
rect 26789 27112 26801 27115
rect 26476 27084 26801 27112
rect 26476 27072 26482 27084
rect 26789 27081 26801 27084
rect 26835 27081 26847 27115
rect 28718 27112 28724 27124
rect 28631 27084 28724 27112
rect 26789 27075 26847 27081
rect 28718 27072 28724 27084
rect 28776 27112 28782 27124
rect 30101 27115 30159 27121
rect 30101 27112 30113 27115
rect 28776 27084 30113 27112
rect 28776 27072 28782 27084
rect 30101 27081 30113 27084
rect 30147 27081 30159 27115
rect 30101 27075 30159 27081
rect 30377 27115 30435 27121
rect 30377 27081 30389 27115
rect 30423 27112 30435 27115
rect 30558 27112 30564 27124
rect 30423 27084 30564 27112
rect 30423 27081 30435 27084
rect 30377 27075 30435 27081
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 38102 27112 38108 27124
rect 38063 27084 38108 27112
rect 38102 27072 38108 27084
rect 38160 27072 38166 27124
rect 41782 27072 41788 27124
rect 41840 27112 41846 27124
rect 42061 27115 42119 27121
rect 42061 27112 42073 27115
rect 41840 27084 42073 27112
rect 41840 27072 41846 27084
rect 42061 27081 42073 27084
rect 42107 27081 42119 27115
rect 42061 27075 42119 27081
rect 43070 27072 43076 27124
rect 43128 27112 43134 27124
rect 43346 27112 43352 27124
rect 43128 27084 43352 27112
rect 43128 27072 43134 27084
rect 43346 27072 43352 27084
rect 43404 27112 43410 27124
rect 44177 27115 44235 27121
rect 44177 27112 44189 27115
rect 43404 27084 44189 27112
rect 43404 27072 43410 27084
rect 44177 27081 44189 27084
rect 44223 27081 44235 27115
rect 44177 27075 44235 27081
rect 45143 27115 45201 27121
rect 45143 27081 45155 27115
rect 45189 27112 45201 27115
rect 46382 27112 46388 27124
rect 45189 27084 46388 27112
rect 45189 27081 45201 27084
rect 45143 27075 45201 27081
rect 46382 27072 46388 27084
rect 46440 27112 46446 27124
rect 47489 27115 47547 27121
rect 47489 27112 47501 27115
rect 46440 27084 47501 27112
rect 46440 27072 46446 27084
rect 47489 27081 47501 27084
rect 47535 27081 47547 27115
rect 47489 27075 47547 27081
rect 22922 27004 22928 27056
rect 22980 27044 22986 27056
rect 24213 27047 24271 27053
rect 24213 27044 24225 27047
rect 22980 27016 24225 27044
rect 22980 27004 22986 27016
rect 24213 27013 24225 27016
rect 24259 27013 24271 27047
rect 24213 27007 24271 27013
rect 24581 27047 24639 27053
rect 24581 27013 24593 27047
rect 24627 27044 24639 27047
rect 29086 27044 29092 27056
rect 24627 27016 27568 27044
rect 29047 27016 29092 27044
rect 24627 27013 24639 27016
rect 24581 27007 24639 27013
rect 14826 26976 14832 26988
rect 14787 26948 14832 26976
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26976 17187 26979
rect 17218 26976 17224 26988
rect 17175 26948 17224 26976
rect 17175 26945 17187 26948
rect 17129 26939 17187 26945
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 18046 26976 18052 26988
rect 18007 26948 18052 26976
rect 18046 26936 18052 26948
rect 18104 26936 18110 26988
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26976 19855 26979
rect 19978 26976 19984 26988
rect 19843 26948 19984 26976
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 21821 26979 21879 26985
rect 21821 26945 21833 26979
rect 21867 26976 21879 26979
rect 21910 26976 21916 26988
rect 21867 26948 21916 26976
rect 21867 26945 21879 26948
rect 21821 26939 21879 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 14366 26908 14372 26920
rect 14327 26880 14372 26908
rect 14366 26868 14372 26880
rect 14424 26868 14430 26920
rect 14734 26908 14740 26920
rect 14695 26880 14740 26908
rect 14734 26868 14740 26880
rect 14792 26868 14798 26920
rect 15102 26868 15108 26920
rect 15160 26908 15166 26920
rect 15749 26911 15807 26917
rect 15749 26908 15761 26911
rect 15160 26880 15761 26908
rect 15160 26868 15166 26880
rect 15749 26877 15761 26880
rect 15795 26908 15807 26911
rect 16114 26908 16120 26920
rect 15795 26880 16120 26908
rect 15795 26877 15807 26880
rect 15749 26871 15807 26877
rect 16114 26868 16120 26880
rect 16172 26868 16178 26920
rect 16390 26908 16396 26920
rect 16351 26880 16396 26908
rect 16390 26868 16396 26880
rect 16448 26868 16454 26920
rect 16574 26868 16580 26920
rect 16632 26908 16638 26920
rect 21082 26908 21088 26920
rect 16632 26880 21088 26908
rect 16632 26868 16638 26880
rect 21082 26868 21088 26880
rect 21140 26868 21146 26920
rect 24029 26911 24087 26917
rect 24029 26877 24041 26911
rect 24075 26908 24087 26911
rect 24596 26908 24624 27007
rect 24854 26976 24860 26988
rect 24815 26948 24860 26976
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 25590 26976 25596 26988
rect 25551 26948 25596 26976
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25038 26908 25044 26920
rect 24075 26880 24624 26908
rect 24999 26880 25044 26908
rect 24075 26877 24087 26880
rect 24029 26871 24087 26877
rect 25038 26868 25044 26880
rect 25096 26868 25102 26920
rect 25498 26908 25504 26920
rect 25459 26880 25504 26908
rect 25498 26868 25504 26880
rect 25556 26868 25562 26920
rect 27540 26917 27568 27016
rect 29086 27004 29092 27016
rect 29144 27004 29150 27056
rect 29270 27004 29276 27056
rect 29328 27044 29334 27056
rect 31018 27044 31024 27056
rect 29328 27016 29408 27044
rect 29328 27004 29334 27016
rect 29380 26985 29408 27016
rect 29840 27016 31024 27044
rect 29840 26988 29868 27016
rect 31018 27004 31024 27016
rect 31076 27044 31082 27056
rect 31076 27016 31248 27044
rect 31076 27004 31082 27016
rect 29365 26979 29423 26985
rect 29365 26945 29377 26979
rect 29411 26945 29423 26979
rect 29822 26976 29828 26988
rect 29783 26948 29828 26976
rect 29365 26939 29423 26945
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 30926 26976 30932 26988
rect 30887 26948 30932 26976
rect 30926 26936 30932 26948
rect 30984 26936 30990 26988
rect 31220 26985 31248 27016
rect 31570 27004 31576 27056
rect 31628 27044 31634 27056
rect 32398 27044 32404 27056
rect 31628 27016 32404 27044
rect 31628 27004 31634 27016
rect 32398 27004 32404 27016
rect 32456 27044 32462 27056
rect 34146 27044 34152 27056
rect 32456 27016 34152 27044
rect 32456 27004 32462 27016
rect 34146 27004 34152 27016
rect 34204 27044 34210 27056
rect 34241 27047 34299 27053
rect 34241 27044 34253 27047
rect 34204 27016 34253 27044
rect 34204 27004 34210 27016
rect 34241 27013 34253 27016
rect 34287 27013 34299 27047
rect 34241 27007 34299 27013
rect 37277 27047 37335 27053
rect 37277 27013 37289 27047
rect 37323 27044 37335 27047
rect 37458 27044 37464 27056
rect 37323 27016 37464 27044
rect 37323 27013 37335 27016
rect 37277 27007 37335 27013
rect 37458 27004 37464 27016
rect 37516 27044 37522 27056
rect 45278 27044 45284 27056
rect 37516 27016 38516 27044
rect 37516 27004 37522 27016
rect 31205 26979 31263 26985
rect 31205 26945 31217 26979
rect 31251 26945 31263 26979
rect 33594 26976 33600 26988
rect 31205 26939 31263 26945
rect 33520 26948 33600 26976
rect 26605 26911 26663 26917
rect 26605 26877 26617 26911
rect 26651 26908 26663 26911
rect 27525 26911 27583 26917
rect 26651 26880 27108 26908
rect 26651 26877 26663 26880
rect 26605 26871 26663 26877
rect 18370 26843 18428 26849
rect 18370 26809 18382 26843
rect 18416 26840 18428 26843
rect 19245 26843 19303 26849
rect 19245 26840 19257 26843
rect 18416 26812 19257 26840
rect 18416 26809 18428 26812
rect 18370 26803 18428 26809
rect 19245 26809 19257 26812
rect 19291 26840 19303 26843
rect 19334 26840 19340 26852
rect 19291 26812 19340 26840
rect 19291 26809 19303 26812
rect 19245 26803 19303 26809
rect 14182 26772 14188 26784
rect 14143 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 15381 26775 15439 26781
rect 15381 26741 15393 26775
rect 15427 26772 15439 26775
rect 15746 26772 15752 26784
rect 15427 26744 15752 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 15930 26772 15936 26784
rect 15891 26744 15936 26772
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 17770 26772 17776 26784
rect 17731 26744 17776 26772
rect 17770 26732 17776 26744
rect 17828 26772 17834 26784
rect 18385 26772 18413 26803
rect 19334 26800 19340 26812
rect 19392 26840 19398 26852
rect 19613 26843 19671 26849
rect 19613 26840 19625 26843
rect 19392 26812 19625 26840
rect 19392 26800 19398 26812
rect 19613 26809 19625 26812
rect 19659 26840 19671 26843
rect 20118 26843 20176 26849
rect 20118 26840 20130 26843
rect 19659 26812 20130 26840
rect 19659 26809 19671 26812
rect 19613 26803 19671 26809
rect 20118 26809 20130 26812
rect 20164 26840 20176 26843
rect 21637 26843 21695 26849
rect 21637 26840 21649 26843
rect 20164 26812 21649 26840
rect 20164 26809 20176 26812
rect 20118 26803 20176 26809
rect 21637 26809 21649 26812
rect 21683 26840 21695 26843
rect 22002 26840 22008 26852
rect 21683 26812 22008 26840
rect 21683 26809 21695 26812
rect 21637 26803 21695 26809
rect 22002 26800 22008 26812
rect 22060 26840 22066 26852
rect 22142 26843 22200 26849
rect 22142 26840 22154 26843
rect 22060 26812 22154 26840
rect 22060 26800 22066 26812
rect 22142 26809 22154 26812
rect 22188 26840 22200 26843
rect 23014 26840 23020 26852
rect 22188 26812 23020 26840
rect 22188 26809 22200 26812
rect 22142 26803 22200 26809
rect 23014 26800 23020 26812
rect 23072 26800 23078 26852
rect 25056 26840 25084 26868
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25056 26812 26065 26840
rect 26053 26809 26065 26812
rect 26099 26840 26111 26843
rect 26970 26840 26976 26852
rect 26099 26812 26976 26840
rect 26099 26809 26111 26812
rect 26053 26803 26111 26809
rect 26970 26800 26976 26812
rect 27028 26800 27034 26852
rect 27080 26784 27108 26880
rect 27525 26877 27537 26911
rect 27571 26908 27583 26911
rect 27890 26908 27896 26920
rect 27571 26880 27896 26908
rect 27571 26877 27583 26880
rect 27525 26871 27583 26877
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 28169 26911 28227 26917
rect 28169 26877 28181 26911
rect 28215 26908 28227 26911
rect 28258 26908 28264 26920
rect 28215 26880 28264 26908
rect 28215 26877 28227 26880
rect 28169 26871 28227 26877
rect 28258 26868 28264 26880
rect 28316 26868 28322 26920
rect 32950 26868 32956 26920
rect 33008 26908 33014 26920
rect 33520 26917 33548 26948
rect 33594 26936 33600 26948
rect 33652 26936 33658 26988
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26976 34023 26979
rect 34885 26979 34943 26985
rect 34885 26976 34897 26979
rect 34011 26948 34897 26976
rect 34011 26945 34023 26948
rect 33965 26939 34023 26945
rect 34885 26945 34897 26948
rect 34931 26976 34943 26979
rect 35250 26976 35256 26988
rect 34931 26948 35256 26976
rect 34931 26945 34943 26948
rect 34885 26939 34943 26945
rect 35250 26936 35256 26948
rect 35308 26936 35314 26988
rect 36722 26976 36728 26988
rect 36683 26948 36728 26976
rect 36722 26936 36728 26948
rect 36780 26936 36786 26988
rect 38289 26979 38347 26985
rect 38289 26945 38301 26979
rect 38335 26976 38347 26979
rect 38378 26976 38384 26988
rect 38335 26948 38384 26976
rect 38335 26945 38347 26948
rect 38289 26939 38347 26945
rect 38378 26936 38384 26948
rect 38436 26936 38442 26988
rect 38488 26976 38516 27016
rect 45020 27016 45284 27044
rect 38565 26979 38623 26985
rect 38565 26976 38577 26979
rect 38488 26948 38577 26976
rect 38565 26945 38577 26948
rect 38611 26945 38623 26979
rect 38565 26939 38623 26945
rect 42705 26979 42763 26985
rect 42705 26945 42717 26979
rect 42751 26976 42763 26979
rect 43254 26976 43260 26988
rect 42751 26948 43260 26976
rect 42751 26945 42763 26948
rect 42705 26939 42763 26945
rect 43254 26936 43260 26948
rect 43312 26936 43318 26988
rect 43898 26976 43904 26988
rect 43859 26948 43904 26976
rect 43898 26936 43904 26948
rect 43956 26936 43962 26988
rect 33045 26911 33103 26917
rect 33045 26908 33057 26911
rect 33008 26880 33057 26908
rect 33008 26868 33014 26880
rect 33045 26877 33057 26880
rect 33091 26908 33103 26911
rect 33505 26911 33563 26917
rect 33505 26908 33517 26911
rect 33091 26880 33517 26908
rect 33091 26877 33103 26880
rect 33045 26871 33103 26877
rect 33505 26877 33517 26880
rect 33551 26877 33563 26911
rect 33505 26871 33563 26877
rect 33781 26911 33839 26917
rect 33781 26877 33793 26911
rect 33827 26908 33839 26911
rect 33870 26908 33876 26920
rect 33827 26880 33876 26908
rect 33827 26877 33839 26880
rect 33781 26871 33839 26877
rect 28350 26840 28356 26852
rect 28311 26812 28356 26840
rect 28350 26800 28356 26812
rect 28408 26800 28414 26852
rect 29086 26800 29092 26852
rect 29144 26840 29150 26852
rect 29434 26843 29492 26849
rect 29434 26840 29446 26843
rect 29144 26812 29446 26840
rect 29144 26800 29150 26812
rect 29434 26809 29446 26812
rect 29480 26809 29492 26843
rect 29434 26803 29492 26809
rect 30745 26843 30803 26849
rect 30745 26809 30757 26843
rect 30791 26840 30803 26843
rect 31021 26843 31079 26849
rect 31021 26840 31033 26843
rect 30791 26812 31033 26840
rect 30791 26809 30803 26812
rect 30745 26803 30803 26809
rect 31021 26809 31033 26812
rect 31067 26840 31079 26843
rect 31110 26840 31116 26852
rect 31067 26812 31116 26840
rect 31067 26809 31079 26812
rect 31021 26803 31079 26809
rect 31110 26800 31116 26812
rect 31168 26800 31174 26852
rect 32769 26843 32827 26849
rect 32769 26809 32781 26843
rect 32815 26840 32827 26843
rect 33796 26840 33824 26871
rect 33870 26868 33876 26880
rect 33928 26908 33934 26920
rect 34330 26908 34336 26920
rect 33928 26880 34336 26908
rect 33928 26868 33934 26880
rect 34330 26868 34336 26880
rect 34388 26868 34394 26920
rect 39666 26868 39672 26920
rect 39724 26908 39730 26920
rect 40494 26908 40500 26920
rect 39724 26880 40500 26908
rect 39724 26868 39730 26880
rect 40494 26868 40500 26880
rect 40552 26868 40558 26920
rect 45020 26917 45048 27016
rect 45278 27004 45284 27016
rect 45336 27004 45342 27056
rect 46750 27044 46756 27056
rect 46711 27016 46756 27044
rect 46750 27004 46756 27016
rect 46808 27004 46814 27056
rect 45020 26911 45098 26917
rect 45020 26880 45052 26911
rect 45040 26877 45052 26880
rect 45086 26877 45098 26911
rect 45040 26871 45098 26877
rect 35206 26843 35264 26849
rect 35206 26840 35218 26843
rect 32815 26812 33824 26840
rect 34164 26812 35218 26840
rect 32815 26809 32827 26812
rect 32769 26803 32827 26809
rect 18966 26772 18972 26784
rect 17828 26744 18413 26772
rect 18927 26744 18972 26772
rect 17828 26732 17834 26744
rect 18966 26732 18972 26744
rect 19024 26732 19030 26784
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 20717 26775 20775 26781
rect 20717 26772 20729 26775
rect 20312 26744 20729 26772
rect 20312 26732 20318 26744
rect 20717 26741 20729 26744
rect 20763 26741 20775 26775
rect 22738 26772 22744 26784
rect 22699 26744 22744 26772
rect 20717 26735 20775 26741
rect 22738 26732 22744 26744
rect 22796 26732 22802 26784
rect 27062 26772 27068 26784
rect 27023 26744 27068 26772
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 30101 26775 30159 26781
rect 30101 26741 30113 26775
rect 30147 26772 30159 26775
rect 32217 26775 32275 26781
rect 32217 26772 32229 26775
rect 30147 26744 32229 26772
rect 30147 26741 30159 26744
rect 30101 26735 30159 26741
rect 32217 26741 32229 26744
rect 32263 26772 32275 26775
rect 32490 26772 32496 26784
rect 32263 26744 32496 26772
rect 32263 26741 32275 26744
rect 32217 26735 32275 26741
rect 32490 26732 32496 26744
rect 32548 26772 32554 26784
rect 34164 26772 34192 26812
rect 34624 26781 34652 26812
rect 35206 26809 35218 26812
rect 35252 26809 35264 26843
rect 35206 26803 35264 26809
rect 35986 26800 35992 26852
rect 36044 26840 36050 26852
rect 36449 26843 36507 26849
rect 36449 26840 36461 26843
rect 36044 26812 36461 26840
rect 36044 26800 36050 26812
rect 36449 26809 36461 26812
rect 36495 26840 36507 26843
rect 36817 26843 36875 26849
rect 36817 26840 36829 26843
rect 36495 26812 36829 26840
rect 36495 26809 36507 26812
rect 36449 26803 36507 26809
rect 36817 26809 36829 26812
rect 36863 26809 36875 26843
rect 36817 26803 36875 26809
rect 37737 26843 37795 26849
rect 37737 26809 37749 26843
rect 37783 26840 37795 26843
rect 38381 26843 38439 26849
rect 38381 26840 38393 26843
rect 37783 26812 38393 26840
rect 37783 26809 37795 26812
rect 37737 26803 37795 26809
rect 38381 26809 38393 26812
rect 38427 26809 38439 26843
rect 38381 26803 38439 26809
rect 39301 26843 39359 26849
rect 39301 26809 39313 26843
rect 39347 26840 39359 26843
rect 39482 26840 39488 26852
rect 39347 26812 39488 26840
rect 39347 26809 39359 26812
rect 39301 26803 39359 26809
rect 32548 26744 34192 26772
rect 34609 26775 34667 26781
rect 32548 26732 32554 26744
rect 34609 26741 34621 26775
rect 34655 26741 34667 26775
rect 34609 26735 34667 26741
rect 35805 26775 35863 26781
rect 35805 26741 35817 26775
rect 35851 26772 35863 26775
rect 35894 26772 35900 26784
rect 35851 26744 35900 26772
rect 35851 26741 35863 26744
rect 35805 26735 35863 26741
rect 35894 26732 35900 26744
rect 35952 26772 35958 26784
rect 36173 26775 36231 26781
rect 36173 26772 36185 26775
rect 35952 26744 36185 26772
rect 35952 26732 35958 26744
rect 36173 26741 36185 26744
rect 36219 26772 36231 26775
rect 37752 26772 37780 26803
rect 39482 26800 39488 26812
rect 39540 26840 39546 26852
rect 40221 26843 40279 26849
rect 40221 26840 40233 26843
rect 39540 26812 40233 26840
rect 39540 26800 39546 26812
rect 40221 26809 40233 26812
rect 40267 26840 40279 26843
rect 40818 26843 40876 26849
rect 40818 26840 40830 26843
rect 40267 26812 40830 26840
rect 40267 26809 40279 26812
rect 40221 26803 40279 26809
rect 40818 26809 40830 26812
rect 40864 26809 40876 26843
rect 40818 26803 40876 26809
rect 43073 26843 43131 26849
rect 43073 26809 43085 26843
rect 43119 26840 43131 26843
rect 43349 26843 43407 26849
rect 43349 26840 43361 26843
rect 43119 26812 43361 26840
rect 43119 26809 43131 26812
rect 43073 26803 43131 26809
rect 43349 26809 43361 26812
rect 43395 26840 43407 26843
rect 43530 26840 43536 26852
rect 43395 26812 43536 26840
rect 43395 26809 43407 26812
rect 43349 26803 43407 26809
rect 43530 26800 43536 26812
rect 43588 26800 43594 26852
rect 43622 26800 43628 26852
rect 43680 26840 43686 26852
rect 44726 26840 44732 26852
rect 43680 26812 44732 26840
rect 43680 26800 43686 26812
rect 44726 26800 44732 26812
rect 44784 26800 44790 26852
rect 46198 26840 46204 26852
rect 46159 26812 46204 26840
rect 46198 26800 46204 26812
rect 46256 26800 46262 26852
rect 46293 26843 46351 26849
rect 46293 26809 46305 26843
rect 46339 26809 46351 26843
rect 46293 26803 46351 26809
rect 39574 26772 39580 26784
rect 36219 26744 37780 26772
rect 39535 26744 39580 26772
rect 36219 26741 36231 26744
rect 36173 26735 36231 26741
rect 39574 26732 39580 26744
rect 39632 26732 39638 26784
rect 41417 26775 41475 26781
rect 41417 26741 41429 26775
rect 41463 26772 41475 26775
rect 41785 26775 41843 26781
rect 41785 26772 41797 26775
rect 41463 26744 41797 26772
rect 41463 26741 41475 26744
rect 41417 26735 41475 26741
rect 41785 26741 41797 26744
rect 41831 26772 41843 26775
rect 41966 26772 41972 26784
rect 41831 26744 41972 26772
rect 41831 26741 41843 26744
rect 41785 26735 41843 26741
rect 41966 26732 41972 26744
rect 42024 26732 42030 26784
rect 44450 26732 44456 26784
rect 44508 26772 44514 26784
rect 44545 26775 44603 26781
rect 44545 26772 44557 26775
rect 44508 26744 44557 26772
rect 44508 26732 44514 26744
rect 44545 26741 44557 26744
rect 44591 26741 44603 26775
rect 44545 26735 44603 26741
rect 45278 26732 45284 26784
rect 45336 26772 45342 26784
rect 45465 26775 45523 26781
rect 45465 26772 45477 26775
rect 45336 26744 45477 26772
rect 45336 26732 45342 26744
rect 45465 26741 45477 26744
rect 45511 26741 45523 26775
rect 45830 26772 45836 26784
rect 45791 26744 45836 26772
rect 45465 26735 45523 26741
rect 45830 26732 45836 26744
rect 45888 26772 45894 26784
rect 46308 26772 46336 26803
rect 47121 26775 47179 26781
rect 47121 26772 47133 26775
rect 45888 26744 47133 26772
rect 45888 26732 45894 26744
rect 47121 26741 47133 26744
rect 47167 26741 47179 26775
rect 47121 26735 47179 26741
rect 1104 26682 48852 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 48852 26682
rect 1104 26608 48852 26630
rect 14734 26528 14740 26580
rect 14792 26568 14798 26580
rect 15105 26571 15163 26577
rect 15105 26568 15117 26571
rect 14792 26540 15117 26568
rect 14792 26528 14798 26540
rect 15105 26537 15117 26540
rect 15151 26568 15163 26571
rect 16390 26568 16396 26580
rect 15151 26540 16396 26568
rect 15151 26537 15163 26540
rect 15105 26531 15163 26537
rect 16390 26528 16396 26540
rect 16448 26568 16454 26580
rect 16485 26571 16543 26577
rect 16485 26568 16497 26571
rect 16448 26540 16497 26568
rect 16448 26528 16454 26540
rect 16485 26537 16497 26540
rect 16531 26537 16543 26571
rect 16485 26531 16543 26537
rect 17126 26528 17132 26580
rect 17184 26568 17190 26580
rect 18046 26568 18052 26580
rect 17184 26540 18052 26568
rect 17184 26528 17190 26540
rect 18046 26528 18052 26540
rect 18104 26528 18110 26580
rect 19150 26528 19156 26580
rect 19208 26568 19214 26580
rect 19337 26571 19395 26577
rect 19337 26568 19349 26571
rect 19208 26540 19349 26568
rect 19208 26528 19214 26540
rect 19337 26537 19349 26540
rect 19383 26537 19395 26571
rect 19337 26531 19395 26537
rect 19889 26571 19947 26577
rect 19889 26537 19901 26571
rect 19935 26568 19947 26571
rect 19978 26568 19984 26580
rect 19935 26540 19984 26568
rect 19935 26537 19947 26540
rect 19889 26531 19947 26537
rect 19978 26528 19984 26540
rect 20036 26528 20042 26580
rect 21450 26568 21456 26580
rect 21411 26540 21456 26568
rect 21450 26528 21456 26540
rect 21508 26528 21514 26580
rect 21910 26568 21916 26580
rect 21871 26540 21916 26568
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 27709 26571 27767 26577
rect 27709 26537 27721 26571
rect 27755 26568 27767 26571
rect 28258 26568 28264 26580
rect 27755 26540 28264 26568
rect 27755 26537 27767 26540
rect 27709 26531 27767 26537
rect 28258 26528 28264 26540
rect 28316 26528 28322 26580
rect 28350 26528 28356 26580
rect 28408 26568 28414 26580
rect 28445 26571 28503 26577
rect 28445 26568 28457 26571
rect 28408 26540 28457 26568
rect 28408 26528 28414 26540
rect 28445 26537 28457 26540
rect 28491 26537 28503 26571
rect 28445 26531 28503 26537
rect 29086 26528 29092 26580
rect 29144 26568 29150 26580
rect 29454 26568 29460 26580
rect 29144 26540 29460 26568
rect 29144 26528 29150 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 30147 26571 30205 26577
rect 30147 26537 30159 26571
rect 30193 26568 30205 26571
rect 30466 26568 30472 26580
rect 30193 26540 30472 26568
rect 30193 26537 30205 26540
rect 30147 26531 30205 26537
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 30926 26568 30932 26580
rect 30887 26540 30932 26568
rect 30926 26528 30932 26540
rect 30984 26528 30990 26580
rect 32214 26528 32220 26580
rect 32272 26568 32278 26580
rect 32677 26571 32735 26577
rect 32677 26568 32689 26571
rect 32272 26540 32689 26568
rect 32272 26528 32278 26540
rect 32677 26537 32689 26540
rect 32723 26537 32735 26571
rect 33413 26571 33471 26577
rect 33413 26568 33425 26571
rect 32677 26531 32735 26537
rect 33106 26540 33425 26568
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 14148 26472 15516 26500
rect 14148 26460 14154 26472
rect 15289 26435 15347 26441
rect 15289 26401 15301 26435
rect 15335 26432 15347 26435
rect 15378 26432 15384 26444
rect 15335 26404 15384 26432
rect 15335 26401 15347 26404
rect 15289 26395 15347 26401
rect 15378 26392 15384 26404
rect 15436 26392 15442 26444
rect 15488 26432 15516 26472
rect 15562 26460 15568 26512
rect 15620 26500 15626 26512
rect 18509 26503 18567 26509
rect 15620 26472 15665 26500
rect 15620 26460 15626 26472
rect 18509 26469 18521 26503
rect 18555 26500 18567 26503
rect 18874 26500 18880 26512
rect 18555 26472 18880 26500
rect 18555 26469 18567 26472
rect 18509 26463 18567 26469
rect 18874 26460 18880 26472
rect 18932 26460 18938 26512
rect 22002 26460 22008 26512
rect 22060 26500 22066 26512
rect 22694 26503 22752 26509
rect 22694 26500 22706 26503
rect 22060 26472 22706 26500
rect 22060 26460 22066 26472
rect 22694 26469 22706 26472
rect 22740 26469 22752 26503
rect 33106 26500 33134 26540
rect 33413 26537 33425 26540
rect 33459 26568 33471 26571
rect 33870 26568 33876 26580
rect 33459 26540 33876 26568
rect 33459 26537 33471 26540
rect 33413 26531 33471 26537
rect 33870 26528 33876 26540
rect 33928 26528 33934 26580
rect 34514 26528 34520 26580
rect 34572 26568 34578 26580
rect 34609 26571 34667 26577
rect 34609 26568 34621 26571
rect 34572 26540 34621 26568
rect 34572 26528 34578 26540
rect 34609 26537 34621 26540
rect 34655 26537 34667 26571
rect 34609 26531 34667 26537
rect 35986 26528 35992 26580
rect 36044 26568 36050 26580
rect 38059 26571 38117 26577
rect 36044 26540 36216 26568
rect 36044 26528 36050 26540
rect 22694 26463 22752 26469
rect 32232 26472 33134 26500
rect 17218 26432 17224 26444
rect 15488 26404 17224 26432
rect 17218 26392 17224 26404
rect 17276 26432 17282 26444
rect 17348 26435 17406 26441
rect 17348 26432 17360 26435
rect 17276 26404 17360 26432
rect 17276 26392 17282 26404
rect 17348 26401 17360 26404
rect 17394 26401 17406 26435
rect 17348 26395 17406 26401
rect 20968 26435 21026 26441
rect 20968 26401 20980 26435
rect 21014 26432 21026 26435
rect 21082 26432 21088 26444
rect 21014 26404 21088 26432
rect 21014 26401 21026 26404
rect 20968 26395 21026 26401
rect 21082 26392 21088 26404
rect 21140 26392 21146 26444
rect 21726 26392 21732 26444
rect 21784 26432 21790 26444
rect 22373 26435 22431 26441
rect 22373 26432 22385 26435
rect 21784 26404 22385 26432
rect 21784 26392 21790 26404
rect 22373 26401 22385 26404
rect 22419 26432 22431 26435
rect 22922 26432 22928 26444
rect 22419 26404 22928 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 22922 26392 22928 26404
rect 22980 26392 22986 26444
rect 23934 26392 23940 26444
rect 23992 26432 23998 26444
rect 24762 26432 24768 26444
rect 23992 26404 24768 26432
rect 23992 26392 23998 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 25225 26435 25283 26441
rect 25225 26401 25237 26435
rect 25271 26432 25283 26435
rect 25498 26432 25504 26444
rect 25271 26404 25504 26432
rect 25271 26401 25283 26404
rect 25225 26395 25283 26401
rect 25498 26392 25504 26404
rect 25556 26432 25562 26444
rect 25777 26435 25835 26441
rect 25777 26432 25789 26435
rect 25556 26404 25789 26432
rect 25556 26392 25562 26404
rect 25777 26401 25789 26404
rect 25823 26432 25835 26435
rect 26697 26435 26755 26441
rect 26697 26432 26709 26435
rect 25823 26404 26709 26432
rect 25823 26401 25835 26404
rect 25777 26395 25835 26401
rect 26697 26401 26709 26404
rect 26743 26401 26755 26435
rect 26697 26395 26755 26401
rect 27040 26435 27098 26441
rect 27040 26401 27052 26435
rect 27086 26432 27098 26435
rect 27154 26432 27160 26444
rect 27086 26404 27160 26432
rect 27086 26401 27098 26404
rect 27040 26395 27098 26401
rect 27154 26392 27160 26404
rect 27212 26392 27218 26444
rect 28902 26392 28908 26444
rect 28960 26432 28966 26444
rect 28997 26435 29055 26441
rect 28997 26432 29009 26435
rect 28960 26404 29009 26432
rect 28960 26392 28966 26404
rect 28997 26401 29009 26404
rect 29043 26401 29055 26435
rect 30006 26432 30012 26444
rect 29967 26404 30012 26432
rect 28997 26395 29055 26401
rect 18414 26364 18420 26376
rect 18375 26336 18420 26364
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18506 26324 18512 26376
rect 18564 26364 18570 26376
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18564 26336 18705 26364
rect 18564 26324 18570 26336
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 25314 26364 25320 26376
rect 25275 26336 25320 26364
rect 18693 26327 18751 26333
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 27893 26367 27951 26373
rect 27893 26333 27905 26367
rect 27939 26364 27951 26367
rect 28074 26364 28080 26376
rect 27939 26336 28080 26364
rect 27939 26333 27951 26336
rect 27893 26327 27951 26333
rect 28074 26324 28080 26336
rect 28132 26324 28138 26376
rect 29012 26364 29040 26395
rect 30006 26392 30012 26404
rect 30064 26392 30070 26444
rect 30926 26392 30932 26444
rect 30984 26432 30990 26444
rect 31056 26435 31114 26441
rect 31056 26432 31068 26435
rect 30984 26404 31068 26432
rect 30984 26392 30990 26404
rect 31056 26401 31068 26404
rect 31102 26432 31114 26435
rect 32030 26432 32036 26444
rect 31102 26404 32036 26432
rect 31102 26401 31114 26404
rect 31056 26395 31114 26401
rect 32030 26392 32036 26404
rect 32088 26392 32094 26444
rect 32122 26392 32128 26444
rect 32180 26432 32186 26444
rect 32232 26441 32260 26472
rect 35618 26460 35624 26512
rect 35676 26500 35682 26512
rect 36078 26500 36084 26512
rect 35676 26472 36084 26500
rect 35676 26460 35682 26472
rect 36078 26460 36084 26472
rect 36136 26460 36142 26512
rect 36188 26509 36216 26540
rect 38059 26537 38071 26571
rect 38105 26568 38117 26571
rect 41138 26568 41144 26580
rect 38105 26540 41144 26568
rect 38105 26537 38117 26540
rect 38059 26531 38117 26537
rect 41138 26528 41144 26540
rect 41196 26528 41202 26580
rect 43898 26568 43904 26580
rect 42444 26540 43904 26568
rect 36173 26503 36231 26509
rect 36173 26469 36185 26503
rect 36219 26469 36231 26503
rect 39666 26500 39672 26512
rect 39627 26472 39672 26500
rect 36173 26463 36231 26469
rect 39666 26460 39672 26472
rect 39724 26460 39730 26512
rect 41877 26503 41935 26509
rect 41877 26469 41889 26503
rect 41923 26500 41935 26503
rect 41966 26500 41972 26512
rect 41923 26472 41972 26500
rect 41923 26469 41935 26472
rect 41877 26463 41935 26469
rect 41966 26460 41972 26472
rect 42024 26460 42030 26512
rect 42444 26509 42472 26540
rect 43898 26528 43904 26540
rect 43956 26528 43962 26580
rect 44358 26528 44364 26580
rect 44416 26568 44422 26580
rect 44545 26571 44603 26577
rect 44545 26568 44557 26571
rect 44416 26540 44557 26568
rect 44416 26528 44422 26540
rect 44545 26537 44557 26540
rect 44591 26537 44603 26571
rect 44545 26531 44603 26537
rect 46198 26528 46204 26580
rect 46256 26568 46262 26580
rect 46661 26571 46719 26577
rect 46661 26568 46673 26571
rect 46256 26540 46673 26568
rect 46256 26528 46262 26540
rect 46661 26537 46673 26540
rect 46707 26537 46719 26571
rect 46661 26531 46719 26537
rect 46842 26528 46848 26580
rect 46900 26568 46906 26580
rect 49510 26568 49516 26580
rect 46900 26540 49516 26568
rect 46900 26528 46906 26540
rect 49510 26528 49516 26540
rect 49568 26528 49574 26580
rect 42429 26503 42487 26509
rect 42429 26469 42441 26503
rect 42475 26469 42487 26503
rect 43530 26500 43536 26512
rect 43491 26472 43536 26500
rect 42429 26463 42487 26469
rect 43530 26460 43536 26472
rect 43588 26460 43594 26512
rect 45830 26500 45836 26512
rect 45791 26472 45836 26500
rect 45830 26460 45836 26472
rect 45888 26460 45894 26512
rect 32217 26435 32275 26441
rect 32217 26432 32229 26435
rect 32180 26404 32229 26432
rect 32180 26392 32186 26404
rect 32217 26401 32229 26404
rect 32263 26401 32275 26435
rect 32217 26395 32275 26401
rect 33229 26435 33287 26441
rect 33229 26401 33241 26435
rect 33275 26432 33287 26435
rect 33318 26432 33324 26444
rect 33275 26404 33324 26432
rect 33275 26401 33287 26404
rect 33229 26395 33287 26401
rect 33318 26392 33324 26404
rect 33376 26432 33382 26444
rect 33962 26432 33968 26444
rect 33376 26404 33968 26432
rect 33376 26392 33382 26404
rect 33962 26392 33968 26404
rect 34020 26392 34026 26444
rect 34241 26435 34299 26441
rect 34241 26401 34253 26435
rect 34287 26432 34299 26435
rect 34422 26432 34428 26444
rect 34287 26404 34428 26432
rect 34287 26401 34299 26404
rect 34241 26395 34299 26401
rect 34422 26392 34428 26404
rect 34480 26392 34486 26444
rect 37829 26435 37887 26441
rect 37829 26401 37841 26435
rect 37875 26432 37887 26435
rect 38010 26432 38016 26444
rect 37875 26404 38016 26432
rect 37875 26401 37887 26404
rect 37829 26395 37887 26401
rect 38010 26392 38016 26404
rect 38068 26392 38074 26444
rect 38838 26392 38844 26444
rect 38896 26432 38902 26444
rect 38933 26435 38991 26441
rect 38933 26432 38945 26435
rect 38896 26404 38945 26432
rect 38896 26392 38902 26404
rect 38933 26401 38945 26404
rect 38979 26401 38991 26435
rect 39390 26432 39396 26444
rect 39351 26404 39396 26432
rect 38933 26395 38991 26401
rect 39390 26392 39396 26404
rect 39448 26392 39454 26444
rect 40532 26435 40590 26441
rect 40532 26401 40544 26435
rect 40578 26401 40590 26435
rect 40532 26395 40590 26401
rect 29546 26364 29552 26376
rect 29012 26336 29552 26364
rect 29546 26324 29552 26336
rect 29604 26364 29610 26376
rect 33042 26364 33048 26376
rect 29604 26336 33048 26364
rect 29604 26324 29610 26336
rect 33042 26324 33048 26336
rect 33100 26324 33106 26376
rect 36354 26364 36360 26376
rect 36315 26336 36360 26364
rect 36354 26324 36360 26336
rect 36412 26324 36418 26376
rect 39206 26324 39212 26376
rect 39264 26364 39270 26376
rect 40547 26364 40575 26395
rect 47118 26392 47124 26444
rect 47176 26432 47182 26444
rect 47248 26435 47306 26441
rect 47248 26432 47260 26435
rect 47176 26404 47260 26432
rect 47176 26392 47182 26404
rect 47248 26401 47260 26404
rect 47294 26401 47306 26435
rect 47248 26395 47306 26401
rect 40678 26364 40684 26376
rect 39264 26336 40684 26364
rect 39264 26324 39270 26336
rect 40678 26324 40684 26336
rect 40736 26324 40742 26376
rect 41601 26367 41659 26373
rect 41601 26333 41613 26367
rect 41647 26364 41659 26367
rect 41785 26367 41843 26373
rect 41785 26364 41797 26367
rect 41647 26336 41797 26364
rect 41647 26333 41659 26336
rect 41601 26327 41659 26333
rect 41785 26333 41797 26336
rect 41831 26364 41843 26367
rect 42518 26364 42524 26376
rect 41831 26336 42524 26364
rect 41831 26333 41843 26336
rect 41785 26327 41843 26333
rect 42518 26324 42524 26336
rect 42576 26324 42582 26376
rect 43441 26367 43499 26373
rect 43441 26333 43453 26367
rect 43487 26364 43499 26367
rect 43622 26364 43628 26376
rect 43487 26336 43628 26364
rect 43487 26333 43499 26336
rect 43441 26327 43499 26333
rect 43622 26324 43628 26336
rect 43680 26324 43686 26376
rect 43714 26324 43720 26376
rect 43772 26364 43778 26376
rect 43772 26336 43817 26364
rect 43772 26324 43778 26336
rect 44818 26324 44824 26376
rect 44876 26364 44882 26376
rect 45741 26367 45799 26373
rect 45741 26364 45753 26367
rect 44876 26336 45753 26364
rect 44876 26324 44882 26336
rect 45741 26333 45753 26336
rect 45787 26364 45799 26367
rect 47351 26367 47409 26373
rect 47351 26364 47363 26367
rect 45787 26336 47363 26364
rect 45787 26333 45799 26336
rect 45741 26327 45799 26333
rect 47351 26333 47363 26336
rect 47397 26333 47409 26367
rect 47351 26327 47409 26333
rect 32401 26299 32459 26305
rect 32401 26265 32413 26299
rect 32447 26296 32459 26299
rect 34146 26296 34152 26308
rect 32447 26268 34152 26296
rect 32447 26265 32459 26268
rect 32401 26259 32459 26265
rect 34146 26256 34152 26268
rect 34204 26256 34210 26308
rect 35161 26299 35219 26305
rect 35161 26265 35173 26299
rect 35207 26296 35219 26299
rect 35986 26296 35992 26308
rect 35207 26268 35992 26296
rect 35207 26265 35219 26268
rect 35161 26259 35219 26265
rect 35986 26256 35992 26268
rect 36044 26256 36050 26308
rect 45554 26256 45560 26308
rect 45612 26296 45618 26308
rect 46293 26299 46351 26305
rect 46293 26296 46305 26299
rect 45612 26268 46305 26296
rect 45612 26256 45618 26268
rect 46293 26265 46305 26268
rect 46339 26265 46351 26299
rect 46293 26259 46351 26265
rect 14366 26228 14372 26240
rect 14327 26200 14372 26228
rect 14366 26188 14372 26200
rect 14424 26188 14430 26240
rect 16209 26231 16267 26237
rect 16209 26197 16221 26231
rect 16255 26228 16267 26231
rect 16390 26228 16396 26240
rect 16255 26200 16396 26228
rect 16255 26197 16267 26200
rect 16209 26191 16267 26197
rect 16390 26188 16396 26200
rect 16448 26188 16454 26240
rect 17451 26231 17509 26237
rect 17451 26197 17463 26231
rect 17497 26228 17509 26231
rect 17954 26228 17960 26240
rect 17497 26200 17960 26228
rect 17497 26197 17509 26200
rect 17451 26191 17509 26197
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 20070 26188 20076 26240
rect 20128 26228 20134 26240
rect 21039 26231 21097 26237
rect 21039 26228 21051 26231
rect 20128 26200 21051 26228
rect 20128 26188 20134 26200
rect 21039 26197 21051 26200
rect 21085 26197 21097 26231
rect 22186 26228 22192 26240
rect 22147 26200 22192 26228
rect 21039 26191 21097 26197
rect 22186 26188 22192 26200
rect 22244 26188 22250 26240
rect 23290 26228 23296 26240
rect 23251 26200 23296 26228
rect 23290 26188 23296 26200
rect 23348 26188 23354 26240
rect 27111 26231 27169 26237
rect 27111 26197 27123 26231
rect 27157 26228 27169 26231
rect 27522 26228 27528 26240
rect 27157 26200 27528 26228
rect 27157 26197 27169 26200
rect 27111 26191 27169 26197
rect 27522 26188 27528 26200
rect 27580 26188 27586 26240
rect 28123 26231 28181 26237
rect 28123 26197 28135 26231
rect 28169 26228 28181 26231
rect 28994 26228 29000 26240
rect 28169 26200 29000 26228
rect 28169 26197 28181 26200
rect 28123 26191 28181 26197
rect 28994 26188 29000 26200
rect 29052 26188 29058 26240
rect 29135 26231 29193 26237
rect 29135 26197 29147 26231
rect 29181 26228 29193 26231
rect 29270 26228 29276 26240
rect 29181 26200 29276 26228
rect 29181 26197 29193 26200
rect 29135 26191 29193 26197
rect 29270 26188 29276 26200
rect 29328 26188 29334 26240
rect 31159 26231 31217 26237
rect 31159 26197 31171 26231
rect 31205 26228 31217 26231
rect 33226 26228 33232 26240
rect 31205 26200 33232 26228
rect 31205 26197 31217 26200
rect 31159 26191 31217 26197
rect 33226 26188 33232 26200
rect 33284 26188 33290 26240
rect 35618 26228 35624 26240
rect 35579 26200 35624 26228
rect 35618 26188 35624 26200
rect 35676 26188 35682 26240
rect 38378 26228 38384 26240
rect 38339 26200 38384 26228
rect 38378 26188 38384 26200
rect 38436 26188 38442 26240
rect 40635 26231 40693 26237
rect 40635 26197 40647 26231
rect 40681 26228 40693 26231
rect 40957 26231 41015 26237
rect 40957 26228 40969 26231
rect 40681 26200 40969 26228
rect 40681 26197 40693 26200
rect 40635 26191 40693 26197
rect 40957 26197 40969 26200
rect 41003 26228 41015 26231
rect 41046 26228 41052 26240
rect 41003 26200 41052 26228
rect 41003 26197 41015 26200
rect 40957 26191 41015 26197
rect 41046 26188 41052 26200
rect 41104 26188 41110 26240
rect 1104 26138 48852 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 48852 26138
rect 1104 26064 48852 26086
rect 15378 25984 15384 26036
rect 15436 26024 15442 26036
rect 16393 26027 16451 26033
rect 16393 26024 16405 26027
rect 15436 25996 16405 26024
rect 15436 25984 15442 25996
rect 16393 25993 16405 25996
rect 16439 25993 16451 26027
rect 16393 25987 16451 25993
rect 16853 26027 16911 26033
rect 16853 25993 16865 26027
rect 16899 26024 16911 26027
rect 18414 26024 18420 26036
rect 16899 25996 18420 26024
rect 16899 25993 16911 25996
rect 16853 25987 16911 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 18966 25984 18972 26036
rect 19024 26024 19030 26036
rect 19245 26027 19303 26033
rect 19245 26024 19257 26027
rect 19024 25996 19257 26024
rect 19024 25984 19030 25996
rect 19245 25993 19257 25996
rect 19291 25993 19303 26027
rect 19245 25987 19303 25993
rect 19886 25984 19892 26036
rect 19944 26024 19950 26036
rect 21361 26027 21419 26033
rect 21361 26024 21373 26027
rect 19944 25996 21373 26024
rect 19944 25984 19950 25996
rect 21361 25993 21373 25996
rect 21407 26024 21419 26027
rect 21726 26024 21732 26036
rect 21407 25996 21732 26024
rect 21407 25993 21419 25996
rect 21361 25987 21419 25993
rect 21726 25984 21732 25996
rect 21784 25984 21790 26036
rect 22922 26024 22928 26036
rect 22883 25996 22928 26024
rect 22922 25984 22928 25996
rect 22980 25984 22986 26036
rect 24762 26024 24768 26036
rect 24723 25996 24768 26024
rect 24762 25984 24768 25996
rect 24820 25984 24826 26036
rect 28074 26024 28080 26036
rect 27987 25996 28080 26024
rect 28074 25984 28080 25996
rect 28132 26024 28138 26036
rect 31846 26024 31852 26036
rect 28132 25996 31852 26024
rect 28132 25984 28138 25996
rect 31846 25984 31852 25996
rect 31904 25984 31910 26036
rect 32122 26024 32128 26036
rect 32083 25996 32128 26024
rect 32122 25984 32128 25996
rect 32180 25984 32186 26036
rect 33318 26024 33324 26036
rect 33279 25996 33324 26024
rect 33318 25984 33324 25996
rect 33376 25984 33382 26036
rect 33919 26027 33977 26033
rect 33919 25993 33931 26027
rect 33965 26024 33977 26027
rect 35618 26024 35624 26036
rect 33965 25996 35624 26024
rect 33965 25993 33977 25996
rect 33919 25987 33977 25993
rect 35618 25984 35624 25996
rect 35676 25984 35682 26036
rect 36495 26027 36553 26033
rect 36495 25993 36507 26027
rect 36541 26024 36553 26027
rect 36722 26024 36728 26036
rect 36541 25996 36728 26024
rect 36541 25993 36553 25996
rect 36495 25987 36553 25993
rect 36722 25984 36728 25996
rect 36780 25984 36786 26036
rect 39390 25984 39396 26036
rect 39448 26024 39454 26036
rect 39577 26027 39635 26033
rect 39577 26024 39589 26027
rect 39448 25996 39589 26024
rect 39448 25984 39454 25996
rect 39577 25993 39589 25996
rect 39623 25993 39635 26027
rect 40678 26024 40684 26036
rect 40639 25996 40684 26024
rect 39577 25987 39635 25993
rect 40678 25984 40684 25996
rect 40736 25984 40742 26036
rect 41966 26024 41972 26036
rect 41927 25996 41972 26024
rect 41966 25984 41972 25996
rect 42024 25984 42030 26036
rect 42521 26027 42579 26033
rect 42521 25993 42533 26027
rect 42567 26024 42579 26027
rect 42889 26027 42947 26033
rect 42567 25996 42794 26024
rect 42567 25993 42579 25996
rect 42521 25987 42579 25993
rect 17954 25916 17960 25968
rect 18012 25956 18018 25968
rect 22186 25956 22192 25968
rect 18012 25928 22192 25956
rect 18012 25916 18018 25928
rect 14826 25888 14832 25900
rect 14787 25860 14832 25888
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 18046 25888 18052 25900
rect 18007 25860 18052 25888
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 20070 25888 20076 25900
rect 20031 25860 20076 25888
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20346 25888 20352 25900
rect 20307 25860 20352 25888
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 21652 25897 21680 25928
rect 22186 25916 22192 25928
rect 22244 25916 22250 25968
rect 24213 25959 24271 25965
rect 24213 25925 24225 25959
rect 24259 25956 24271 25959
rect 28092 25956 28120 25984
rect 28902 25956 28908 25968
rect 24259 25928 28120 25956
rect 28505 25928 28908 25956
rect 24259 25925 24271 25928
rect 24213 25919 24271 25925
rect 21637 25891 21695 25897
rect 21637 25857 21649 25891
rect 21683 25857 21695 25891
rect 21637 25851 21695 25857
rect 22002 25848 22008 25900
rect 22060 25888 22066 25900
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22060 25860 22569 25888
rect 22060 25848 22066 25860
rect 22557 25857 22569 25860
rect 22603 25888 22615 25891
rect 22741 25891 22799 25897
rect 22741 25888 22753 25891
rect 22603 25860 22753 25888
rect 22603 25857 22615 25860
rect 22557 25851 22615 25857
rect 22741 25857 22753 25860
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 17770 25820 17776 25832
rect 16040 25792 17776 25820
rect 16040 25761 16068 25792
rect 17770 25780 17776 25792
rect 17828 25780 17834 25832
rect 23658 25820 23664 25832
rect 23622 25792 23664 25820
rect 23658 25780 23664 25792
rect 23716 25829 23722 25832
rect 23716 25823 23770 25829
rect 23716 25789 23724 25823
rect 23758 25820 23770 25823
rect 24228 25820 24256 25919
rect 25590 25888 25596 25900
rect 25551 25860 25596 25888
rect 25590 25848 25596 25860
rect 25648 25848 25654 25900
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 28505 25888 28533 25928
rect 28902 25916 28908 25928
rect 28960 25956 28966 25968
rect 29089 25959 29147 25965
rect 29089 25956 29101 25959
rect 28960 25928 29101 25956
rect 28960 25916 28966 25928
rect 29089 25925 29101 25928
rect 29135 25925 29147 25959
rect 29089 25919 29147 25925
rect 30006 25916 30012 25968
rect 30064 25956 30070 25968
rect 30377 25959 30435 25965
rect 30377 25956 30389 25959
rect 30064 25928 30389 25956
rect 30064 25916 30070 25928
rect 30377 25925 30389 25928
rect 30423 25956 30435 25959
rect 33686 25956 33692 25968
rect 30423 25928 33692 25956
rect 30423 25925 30435 25928
rect 30377 25919 30435 25925
rect 33686 25916 33692 25928
rect 33744 25916 33750 25968
rect 42766 25956 42794 25996
rect 42889 25993 42901 26027
rect 42935 26024 42947 26027
rect 43257 26027 43315 26033
rect 43257 26024 43269 26027
rect 42935 25996 43269 26024
rect 42935 25993 42947 25996
rect 42889 25987 42947 25993
rect 43257 25993 43269 25996
rect 43303 26024 43315 26027
rect 43530 26024 43536 26036
rect 43303 25996 43536 26024
rect 43303 25993 43315 25996
rect 43257 25987 43315 25993
rect 43530 25984 43536 25996
rect 43588 25984 43594 26036
rect 44818 26024 44824 26036
rect 44779 25996 44824 26024
rect 44818 25984 44824 25996
rect 44876 25984 44882 26036
rect 45830 26024 45836 26036
rect 45791 25996 45836 26024
rect 45830 25984 45836 25996
rect 45888 25984 45894 26036
rect 46198 25984 46204 26036
rect 46256 26024 46262 26036
rect 46385 26027 46443 26033
rect 46385 26024 46397 26027
rect 46256 25996 46397 26024
rect 46256 25984 46262 25996
rect 46385 25993 46397 25996
rect 46431 25993 46443 26027
rect 46385 25987 46443 25993
rect 43622 25956 43628 25968
rect 33796 25928 36435 25956
rect 42766 25928 43628 25956
rect 26108 25860 28533 25888
rect 26108 25848 26114 25860
rect 28994 25848 29000 25900
rect 29052 25888 29058 25900
rect 29365 25891 29423 25897
rect 29365 25888 29377 25891
rect 29052 25860 29377 25888
rect 29052 25848 29058 25860
rect 29365 25857 29377 25860
rect 29411 25888 29423 25891
rect 29730 25888 29736 25900
rect 29411 25860 29736 25888
rect 29411 25857 29423 25860
rect 29365 25851 29423 25857
rect 29730 25848 29736 25860
rect 29788 25848 29794 25900
rect 31757 25891 31815 25897
rect 31757 25857 31769 25891
rect 31803 25888 31815 25891
rect 33796 25888 33824 25928
rect 34701 25891 34759 25897
rect 34701 25888 34713 25891
rect 31803 25860 33824 25888
rect 33863 25860 34713 25888
rect 31803 25857 31815 25860
rect 31757 25851 31815 25857
rect 23758 25792 24256 25820
rect 27065 25823 27123 25829
rect 23758 25789 23770 25792
rect 23716 25783 23770 25789
rect 27065 25789 27077 25823
rect 27111 25820 27123 25823
rect 27154 25820 27160 25832
rect 27111 25792 27160 25820
rect 27111 25789 27123 25792
rect 27065 25783 27123 25789
rect 23716 25780 23722 25783
rect 27154 25780 27160 25792
rect 27212 25820 27218 25832
rect 27982 25820 27988 25832
rect 27212 25792 27988 25820
rect 27212 25780 27218 25792
rect 27982 25780 27988 25792
rect 28040 25780 28046 25832
rect 28220 25823 28278 25829
rect 28220 25789 28232 25823
rect 28266 25820 28278 25823
rect 28718 25820 28724 25832
rect 28266 25792 28724 25820
rect 28266 25789 28278 25792
rect 28220 25783 28278 25789
rect 28718 25780 28724 25792
rect 28776 25780 28782 25832
rect 30190 25780 30196 25832
rect 30248 25820 30254 25832
rect 31272 25823 31330 25829
rect 31272 25820 31284 25823
rect 30248 25792 31284 25820
rect 30248 25780 30254 25792
rect 31272 25789 31284 25792
rect 31318 25820 31330 25823
rect 31772 25820 31800 25851
rect 31318 25792 31800 25820
rect 31318 25789 31330 25792
rect 31272 25783 31330 25789
rect 32030 25780 32036 25832
rect 32088 25820 32094 25832
rect 32252 25823 32310 25829
rect 32252 25820 32264 25823
rect 32088 25792 32264 25820
rect 32088 25780 32094 25792
rect 32252 25789 32264 25792
rect 32298 25820 32310 25823
rect 32674 25820 32680 25832
rect 32298 25792 32680 25820
rect 32298 25789 32310 25792
rect 32252 25783 32310 25789
rect 32674 25780 32680 25792
rect 32732 25780 32738 25832
rect 33042 25780 33048 25832
rect 33100 25820 33106 25832
rect 33863 25829 33891 25860
rect 34701 25857 34713 25860
rect 34747 25888 34759 25891
rect 34790 25888 34796 25900
rect 34747 25860 34796 25888
rect 34747 25857 34759 25860
rect 34701 25851 34759 25857
rect 34790 25848 34796 25860
rect 34848 25848 34854 25900
rect 36407 25829 36435 25928
rect 43622 25916 43628 25928
rect 43680 25956 43686 25968
rect 45051 25959 45109 25965
rect 45051 25956 45063 25959
rect 43680 25928 45063 25956
rect 43680 25916 43686 25928
rect 45051 25925 45063 25928
rect 45097 25925 45109 25959
rect 45051 25919 45109 25925
rect 37645 25891 37703 25897
rect 37645 25857 37657 25891
rect 37691 25888 37703 25891
rect 38933 25891 38991 25897
rect 37691 25860 38792 25888
rect 37691 25857 37703 25860
rect 37645 25851 37703 25857
rect 38764 25832 38792 25860
rect 38933 25857 38945 25891
rect 38979 25888 38991 25891
rect 39574 25888 39580 25900
rect 38979 25860 39580 25888
rect 38979 25857 38991 25860
rect 38933 25851 38991 25857
rect 39574 25848 39580 25860
rect 39632 25848 39638 25900
rect 41046 25888 41052 25900
rect 41007 25860 41052 25888
rect 41046 25848 41052 25860
rect 41104 25848 41110 25900
rect 41690 25888 41696 25900
rect 41603 25860 41696 25888
rect 41690 25848 41696 25860
rect 41748 25888 41754 25900
rect 42058 25888 42064 25900
rect 41748 25860 42064 25888
rect 41748 25848 41754 25860
rect 42058 25848 42064 25860
rect 42116 25848 42122 25900
rect 43441 25891 43499 25897
rect 43441 25857 43453 25891
rect 43487 25888 43499 25891
rect 43487 25860 44496 25888
rect 43487 25857 43499 25860
rect 43441 25851 43499 25857
rect 33848 25823 33906 25829
rect 33848 25820 33860 25823
rect 33100 25792 33860 25820
rect 33100 25780 33106 25792
rect 33848 25789 33860 25792
rect 33894 25789 33906 25823
rect 33848 25783 33906 25789
rect 34952 25823 35010 25829
rect 34952 25789 34964 25823
rect 34998 25820 35010 25823
rect 36407 25823 36482 25829
rect 34998 25792 35388 25820
rect 36407 25792 36436 25823
rect 34998 25789 35010 25792
rect 34952 25783 35010 25789
rect 15191 25755 15249 25761
rect 15191 25721 15203 25755
rect 15237 25721 15249 25755
rect 16025 25755 16083 25761
rect 16025 25752 16037 25755
rect 15191 25715 15249 25721
rect 15488 25724 16037 25752
rect 14737 25687 14795 25693
rect 14737 25653 14749 25687
rect 14783 25684 14795 25687
rect 15206 25684 15234 25715
rect 15488 25696 15516 25724
rect 16025 25721 16037 25724
rect 16071 25721 16083 25755
rect 16025 25715 16083 25721
rect 17218 25712 17224 25764
rect 17276 25752 17282 25764
rect 17405 25755 17463 25761
rect 17405 25752 17417 25755
rect 17276 25724 17417 25752
rect 17276 25712 17282 25724
rect 17405 25721 17417 25724
rect 17451 25721 17463 25755
rect 17788 25752 17816 25780
rect 18370 25755 18428 25761
rect 18370 25752 18382 25755
rect 17788 25724 18382 25752
rect 17405 25715 17463 25721
rect 18370 25721 18382 25724
rect 18416 25721 18428 25755
rect 18370 25715 18428 25721
rect 19889 25755 19947 25761
rect 19889 25721 19901 25755
rect 19935 25752 19947 25755
rect 20165 25755 20223 25761
rect 20165 25752 20177 25755
rect 19935 25724 20177 25752
rect 19935 25721 19947 25724
rect 19889 25715 19947 25721
rect 20165 25721 20177 25724
rect 20211 25752 20223 25755
rect 20254 25752 20260 25764
rect 20211 25724 20260 25752
rect 20211 25721 20223 25724
rect 20165 25715 20223 25721
rect 20254 25712 20260 25724
rect 20312 25712 20318 25764
rect 20346 25712 20352 25764
rect 20404 25752 20410 25764
rect 21726 25752 21732 25764
rect 20404 25724 21490 25752
rect 21687 25724 21732 25752
rect 20404 25712 20410 25724
rect 15470 25684 15476 25696
rect 14783 25656 15476 25684
rect 14783 25653 14795 25656
rect 14737 25647 14795 25653
rect 15470 25644 15476 25656
rect 15528 25644 15534 25696
rect 15746 25684 15752 25696
rect 15707 25656 15752 25684
rect 15746 25644 15752 25656
rect 15804 25644 15810 25696
rect 16945 25687 17003 25693
rect 16945 25653 16957 25687
rect 16991 25684 17003 25687
rect 17310 25684 17316 25696
rect 16991 25656 17316 25684
rect 16991 25653 17003 25656
rect 16945 25647 17003 25653
rect 17310 25644 17316 25656
rect 17368 25644 17374 25696
rect 18966 25684 18972 25696
rect 18927 25656 18972 25684
rect 18966 25644 18972 25656
rect 19024 25644 19030 25696
rect 21082 25684 21088 25696
rect 21043 25656 21088 25684
rect 21082 25644 21088 25656
rect 21140 25644 21146 25696
rect 21462 25684 21490 25724
rect 21726 25712 21732 25724
rect 21784 25712 21790 25764
rect 22281 25755 22339 25761
rect 22281 25721 22293 25755
rect 22327 25721 22339 25755
rect 22281 25715 22339 25721
rect 22296 25684 22324 25715
rect 22462 25712 22468 25764
rect 22520 25752 22526 25764
rect 23799 25755 23857 25761
rect 23799 25752 23811 25755
rect 22520 25724 23811 25752
rect 22520 25712 22526 25724
rect 23799 25721 23811 25724
rect 23845 25721 23857 25755
rect 25130 25752 25136 25764
rect 23799 25715 23857 25721
rect 24044 25724 25136 25752
rect 21462 25656 22324 25684
rect 22741 25687 22799 25693
rect 22741 25653 22753 25687
rect 22787 25684 22799 25687
rect 24044 25684 24072 25724
rect 25130 25712 25136 25724
rect 25188 25752 25194 25764
rect 25409 25755 25467 25761
rect 25409 25752 25421 25755
rect 25188 25724 25421 25752
rect 25188 25712 25194 25724
rect 25409 25721 25421 25724
rect 25455 25752 25467 25755
rect 25914 25755 25972 25761
rect 25914 25752 25926 25755
rect 25455 25724 25926 25752
rect 25455 25721 25467 25724
rect 25409 25715 25467 25721
rect 25914 25721 25926 25724
rect 25960 25752 25972 25755
rect 26878 25752 26884 25764
rect 25960 25724 26884 25752
rect 25960 25721 25972 25724
rect 25914 25715 25972 25721
rect 26878 25712 26884 25724
rect 26936 25712 26942 25764
rect 28307 25755 28365 25761
rect 28307 25721 28319 25755
rect 28353 25752 28365 25755
rect 28810 25752 28816 25764
rect 28353 25724 28816 25752
rect 28353 25721 28365 25724
rect 28307 25715 28365 25721
rect 28810 25712 28816 25724
rect 28868 25712 28874 25764
rect 28902 25712 28908 25764
rect 28960 25752 28966 25764
rect 29454 25752 29460 25764
rect 28960 25724 29460 25752
rect 28960 25712 28966 25724
rect 29454 25712 29460 25724
rect 29512 25712 29518 25764
rect 30006 25752 30012 25764
rect 29967 25724 30012 25752
rect 30006 25712 30012 25724
rect 30064 25712 30070 25764
rect 35360 25696 35388 25792
rect 36424 25789 36436 25792
rect 36470 25820 36482 25823
rect 38470 25820 38476 25832
rect 36470 25792 36952 25820
rect 38431 25792 38476 25820
rect 36470 25789 36482 25792
rect 36424 25783 36482 25789
rect 22787 25656 24072 25684
rect 26513 25687 26571 25693
rect 22787 25653 22799 25656
rect 22741 25647 22799 25653
rect 26513 25653 26525 25687
rect 26559 25684 26571 25687
rect 26694 25684 26700 25696
rect 26559 25656 26700 25684
rect 26559 25653 26571 25656
rect 26513 25647 26571 25653
rect 26694 25644 26700 25656
rect 26752 25644 26758 25696
rect 30926 25644 30932 25696
rect 30984 25684 30990 25696
rect 31021 25687 31079 25693
rect 31021 25684 31033 25687
rect 30984 25656 31033 25684
rect 30984 25644 30990 25656
rect 31021 25653 31033 25656
rect 31067 25653 31079 25687
rect 31021 25647 31079 25653
rect 31343 25687 31401 25693
rect 31343 25653 31355 25687
rect 31389 25684 31401 25687
rect 31662 25684 31668 25696
rect 31389 25656 31668 25684
rect 31389 25653 31401 25656
rect 31343 25647 31401 25653
rect 31662 25644 31668 25656
rect 31720 25644 31726 25696
rect 32122 25644 32128 25696
rect 32180 25684 32186 25696
rect 32355 25687 32413 25693
rect 32355 25684 32367 25687
rect 32180 25656 32367 25684
rect 32180 25644 32186 25656
rect 32355 25653 32367 25656
rect 32401 25653 32413 25687
rect 32355 25647 32413 25653
rect 34333 25687 34391 25693
rect 34333 25653 34345 25687
rect 34379 25684 34391 25687
rect 34514 25684 34520 25696
rect 34379 25656 34520 25684
rect 34379 25653 34391 25656
rect 34333 25647 34391 25653
rect 34514 25644 34520 25656
rect 34572 25644 34578 25696
rect 34790 25644 34796 25696
rect 34848 25684 34854 25696
rect 35023 25687 35081 25693
rect 35023 25684 35035 25687
rect 34848 25656 35035 25684
rect 34848 25644 34854 25656
rect 35023 25653 35035 25656
rect 35069 25653 35081 25687
rect 35342 25684 35348 25696
rect 35303 25656 35348 25684
rect 35023 25647 35081 25653
rect 35342 25644 35348 25656
rect 35400 25644 35406 25696
rect 35986 25684 35992 25696
rect 35947 25656 35992 25684
rect 35986 25644 35992 25656
rect 36044 25644 36050 25696
rect 36924 25693 36952 25792
rect 38470 25780 38476 25792
rect 38528 25780 38534 25832
rect 38746 25820 38752 25832
rect 38707 25792 38752 25820
rect 38746 25780 38752 25792
rect 38804 25780 38810 25832
rect 40126 25712 40132 25764
rect 40184 25752 40190 25764
rect 41046 25752 41052 25764
rect 40184 25724 41052 25752
rect 40184 25712 40190 25724
rect 41046 25712 41052 25724
rect 41104 25752 41110 25764
rect 41141 25755 41199 25761
rect 41141 25752 41153 25755
rect 41104 25724 41153 25752
rect 41104 25712 41110 25724
rect 41141 25721 41153 25724
rect 41187 25752 41199 25755
rect 43530 25752 43536 25764
rect 41187 25724 43536 25752
rect 41187 25721 41199 25724
rect 41141 25715 41199 25721
rect 43530 25712 43536 25724
rect 43588 25712 43594 25764
rect 44468 25761 44496 25860
rect 44726 25780 44732 25832
rect 44784 25820 44790 25832
rect 44948 25823 45006 25829
rect 44948 25820 44960 25823
rect 44784 25792 44960 25820
rect 44784 25780 44790 25792
rect 44948 25789 44960 25792
rect 44994 25820 45006 25823
rect 45370 25820 45376 25832
rect 44994 25792 45376 25820
rect 44994 25789 45006 25792
rect 44948 25783 45006 25789
rect 45370 25780 45376 25792
rect 45428 25780 45434 25832
rect 45462 25780 45468 25832
rect 45520 25820 45526 25832
rect 46144 25823 46202 25829
rect 46144 25820 46156 25823
rect 45520 25792 46156 25820
rect 45520 25780 45526 25792
rect 46144 25789 46156 25792
rect 46190 25820 46202 25823
rect 46569 25823 46627 25829
rect 46569 25820 46581 25823
rect 46190 25792 46581 25820
rect 46190 25789 46202 25792
rect 46144 25783 46202 25789
rect 46569 25789 46581 25792
rect 46615 25789 46627 25823
rect 46569 25783 46627 25789
rect 47026 25780 47032 25832
rect 47084 25820 47090 25832
rect 47156 25823 47214 25829
rect 47156 25820 47168 25823
rect 47084 25792 47168 25820
rect 47084 25780 47090 25792
rect 47156 25789 47168 25792
rect 47202 25820 47214 25823
rect 47949 25823 48007 25829
rect 47949 25820 47961 25823
rect 47202 25792 47961 25820
rect 47202 25789 47214 25792
rect 47156 25783 47214 25789
rect 47949 25789 47961 25792
rect 47995 25789 48007 25823
rect 47949 25783 48007 25789
rect 44085 25755 44143 25761
rect 44085 25721 44097 25755
rect 44131 25721 44143 25755
rect 44085 25715 44143 25721
rect 44453 25755 44511 25761
rect 44453 25721 44465 25755
rect 44499 25752 44511 25755
rect 47259 25755 47317 25761
rect 47259 25752 47271 25755
rect 44499 25724 47271 25752
rect 44499 25721 44511 25724
rect 44453 25715 44511 25721
rect 47259 25721 47271 25724
rect 47305 25721 47317 25755
rect 47259 25715 47317 25721
rect 36909 25687 36967 25693
rect 36909 25653 36921 25687
rect 36955 25684 36967 25687
rect 37274 25684 37280 25696
rect 36955 25656 37280 25684
rect 36955 25653 36967 25656
rect 36909 25647 36967 25653
rect 37274 25644 37280 25656
rect 37332 25644 37338 25696
rect 38010 25684 38016 25696
rect 37971 25656 38016 25684
rect 38010 25644 38016 25656
rect 38068 25644 38074 25696
rect 38838 25644 38844 25696
rect 38896 25684 38902 25696
rect 39209 25687 39267 25693
rect 39209 25684 39221 25687
rect 38896 25656 39221 25684
rect 38896 25644 38902 25656
rect 39209 25653 39221 25656
rect 39255 25653 39267 25687
rect 39209 25647 39267 25653
rect 43346 25644 43352 25696
rect 43404 25684 43410 25696
rect 44100 25684 44128 25715
rect 46566 25684 46572 25696
rect 43404 25656 46572 25684
rect 43404 25644 43410 25656
rect 46566 25644 46572 25656
rect 46624 25644 46630 25696
rect 46658 25644 46664 25696
rect 46716 25684 46722 25696
rect 47118 25684 47124 25696
rect 46716 25656 47124 25684
rect 46716 25644 46722 25656
rect 47118 25644 47124 25656
rect 47176 25684 47182 25696
rect 47581 25687 47639 25693
rect 47581 25684 47593 25687
rect 47176 25656 47593 25684
rect 47176 25644 47182 25656
rect 47581 25653 47593 25656
rect 47627 25653 47639 25687
rect 47581 25647 47639 25653
rect 1104 25594 48852 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 48852 25594
rect 1104 25520 48852 25542
rect 14826 25480 14832 25492
rect 14787 25452 14832 25480
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 15746 25440 15752 25492
rect 15804 25480 15810 25492
rect 16206 25480 16212 25492
rect 15804 25452 16212 25480
rect 15804 25440 15810 25452
rect 16206 25440 16212 25452
rect 16264 25480 16270 25492
rect 16485 25483 16543 25489
rect 16485 25480 16497 25483
rect 16264 25452 16497 25480
rect 16264 25440 16270 25452
rect 16485 25449 16497 25452
rect 16531 25449 16543 25483
rect 20070 25480 20076 25492
rect 20031 25452 20076 25480
rect 16485 25443 16543 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 21683 25483 21741 25489
rect 21683 25449 21695 25483
rect 21729 25480 21741 25483
rect 23661 25483 23719 25489
rect 23661 25480 23673 25483
rect 21729 25452 23673 25480
rect 21729 25449 21741 25452
rect 21683 25443 21741 25449
rect 23661 25449 23673 25452
rect 23707 25480 23719 25483
rect 23750 25480 23756 25492
rect 23707 25452 23756 25480
rect 23707 25449 23719 25452
rect 23661 25443 23719 25449
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 24765 25483 24823 25489
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 25498 25480 25504 25492
rect 24811 25452 25504 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 25869 25483 25927 25489
rect 25869 25480 25881 25483
rect 25648 25452 25881 25480
rect 25648 25440 25654 25452
rect 25869 25449 25881 25452
rect 25915 25449 25927 25483
rect 26878 25480 26884 25492
rect 26839 25452 26884 25480
rect 25869 25443 25927 25449
rect 26878 25440 26884 25452
rect 26936 25440 26942 25492
rect 29730 25480 29736 25492
rect 29691 25452 29736 25480
rect 29730 25440 29736 25452
rect 29788 25440 29794 25492
rect 31662 25440 31668 25492
rect 31720 25480 31726 25492
rect 31849 25483 31907 25489
rect 31849 25480 31861 25483
rect 31720 25452 31861 25480
rect 31720 25440 31726 25452
rect 31849 25449 31861 25452
rect 31895 25449 31907 25483
rect 31849 25443 31907 25449
rect 34333 25483 34391 25489
rect 34333 25449 34345 25483
rect 34379 25480 34391 25483
rect 34422 25480 34428 25492
rect 34379 25452 34428 25480
rect 34379 25449 34391 25452
rect 34333 25443 34391 25449
rect 15470 25372 15476 25424
rect 15528 25412 15534 25424
rect 15610 25415 15668 25421
rect 15610 25412 15622 25415
rect 15528 25384 15622 25412
rect 15528 25372 15534 25384
rect 15610 25381 15622 25384
rect 15656 25381 15668 25415
rect 15610 25375 15668 25381
rect 16390 25372 16396 25424
rect 16448 25412 16454 25424
rect 17126 25412 17132 25424
rect 16448 25384 17132 25412
rect 16448 25372 16454 25384
rect 17126 25372 17132 25384
rect 17184 25412 17190 25424
rect 17221 25415 17279 25421
rect 17221 25412 17233 25415
rect 17184 25384 17233 25412
rect 17184 25372 17190 25384
rect 17221 25381 17233 25384
rect 17267 25381 17279 25415
rect 17221 25375 17279 25381
rect 17310 25372 17316 25424
rect 17368 25412 17374 25424
rect 18690 25412 18696 25424
rect 17368 25384 18696 25412
rect 17368 25372 17374 25384
rect 18690 25372 18696 25384
rect 18748 25372 18754 25424
rect 18785 25415 18843 25421
rect 18785 25381 18797 25415
rect 18831 25412 18843 25415
rect 18966 25412 18972 25424
rect 18831 25384 18972 25412
rect 18831 25381 18843 25384
rect 18785 25375 18843 25381
rect 18966 25372 18972 25384
rect 19024 25372 19030 25424
rect 21082 25372 21088 25424
rect 21140 25412 21146 25424
rect 21910 25412 21916 25424
rect 21140 25384 21916 25412
rect 21140 25372 21146 25384
rect 21910 25372 21916 25384
rect 21968 25372 21974 25424
rect 22097 25415 22155 25421
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 22186 25412 22192 25424
rect 22143 25384 22192 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 22186 25372 22192 25384
rect 22244 25412 22250 25424
rect 22738 25412 22744 25424
rect 22244 25384 22744 25412
rect 22244 25372 22250 25384
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 25038 25412 25044 25424
rect 24999 25384 25044 25412
rect 25038 25372 25044 25384
rect 25096 25372 25102 25424
rect 28902 25412 28908 25424
rect 28863 25384 28908 25412
rect 28902 25372 28908 25384
rect 28960 25372 28966 25424
rect 30558 25372 30564 25424
rect 30616 25412 30622 25424
rect 30653 25415 30711 25421
rect 30653 25412 30665 25415
rect 30616 25384 30665 25412
rect 30616 25372 30622 25384
rect 30653 25381 30665 25384
rect 30699 25381 30711 25415
rect 30653 25375 30711 25381
rect 14918 25304 14924 25356
rect 14976 25344 14982 25356
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 14976 25316 15301 25344
rect 14976 25304 14982 25316
rect 15289 25313 15301 25316
rect 15335 25344 15347 25347
rect 15930 25344 15936 25356
rect 15335 25316 15936 25344
rect 15335 25313 15347 25316
rect 15289 25307 15347 25313
rect 15930 25304 15936 25316
rect 15988 25304 15994 25356
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 17862 25344 17868 25356
rect 17819 25316 17868 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 17862 25304 17868 25316
rect 17920 25344 17926 25356
rect 18506 25344 18512 25356
rect 17920 25316 18512 25344
rect 17920 25304 17926 25316
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 21453 25347 21511 25353
rect 21453 25344 21465 25347
rect 19484 25316 21465 25344
rect 19484 25304 19490 25316
rect 21453 25313 21465 25316
rect 21499 25344 21511 25347
rect 21542 25344 21548 25356
rect 21499 25316 21548 25344
rect 21499 25313 21511 25316
rect 21453 25307 21511 25313
rect 21542 25304 21548 25316
rect 21600 25304 21606 25356
rect 26510 25344 26516 25356
rect 26471 25316 26516 25344
rect 26510 25304 26516 25316
rect 26568 25304 26574 25356
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25276 17187 25279
rect 17402 25276 17408 25288
rect 17175 25248 17408 25276
rect 17175 25245 17187 25248
rect 17129 25239 17187 25245
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 18414 25236 18420 25288
rect 18472 25276 18478 25288
rect 18969 25279 19027 25285
rect 18969 25276 18981 25279
rect 18472 25248 18981 25276
rect 18472 25236 18478 25248
rect 18969 25245 18981 25248
rect 19015 25276 19027 25279
rect 20346 25276 20352 25288
rect 19015 25248 20352 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 22646 25276 22652 25288
rect 22607 25248 22652 25276
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 23293 25279 23351 25285
rect 23293 25245 23305 25279
rect 23339 25276 23351 25279
rect 23934 25276 23940 25288
rect 23339 25248 23940 25276
rect 23339 25245 23351 25248
rect 23293 25239 23351 25245
rect 23934 25236 23940 25248
rect 23992 25276 23998 25288
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 23992 25248 24961 25276
rect 23992 25236 23998 25248
rect 24949 25245 24961 25248
rect 24995 25245 25007 25279
rect 25590 25276 25596 25288
rect 25551 25248 25596 25276
rect 24949 25239 25007 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 28810 25276 28816 25288
rect 28771 25248 28816 25276
rect 28810 25236 28816 25248
rect 28868 25236 28874 25288
rect 29457 25279 29515 25285
rect 29457 25245 29469 25279
rect 29503 25276 29515 25279
rect 30374 25276 30380 25288
rect 29503 25248 30380 25276
rect 29503 25245 29515 25248
rect 29457 25239 29515 25245
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30558 25276 30564 25288
rect 30519 25248 30564 25276
rect 30558 25236 30564 25248
rect 30616 25236 30622 25288
rect 30837 25279 30895 25285
rect 30837 25245 30849 25279
rect 30883 25245 30895 25279
rect 31864 25276 31892 25443
rect 34422 25440 34428 25452
rect 34480 25440 34486 25492
rect 34701 25483 34759 25489
rect 34701 25449 34713 25483
rect 34747 25480 34759 25483
rect 34790 25480 34796 25492
rect 34747 25452 34796 25480
rect 34747 25449 34759 25452
rect 34701 25443 34759 25449
rect 34790 25440 34796 25452
rect 34848 25440 34854 25492
rect 36078 25480 36084 25492
rect 36039 25452 36084 25480
rect 36078 25440 36084 25452
rect 36136 25440 36142 25492
rect 36495 25483 36553 25489
rect 36495 25449 36507 25483
rect 36541 25480 36553 25483
rect 38378 25480 38384 25492
rect 36541 25452 38384 25480
rect 36541 25449 36553 25452
rect 36495 25443 36553 25449
rect 38378 25440 38384 25452
rect 38436 25440 38442 25492
rect 41046 25480 41052 25492
rect 41007 25452 41052 25480
rect 41046 25440 41052 25452
rect 41104 25440 41110 25492
rect 32306 25372 32312 25424
rect 32364 25412 32370 25424
rect 32364 25384 32409 25412
rect 32364 25372 32370 25384
rect 34606 25372 34612 25424
rect 34664 25412 34670 25424
rect 34977 25415 35035 25421
rect 34977 25412 34989 25415
rect 34664 25384 34989 25412
rect 34664 25372 34670 25384
rect 34977 25381 34989 25384
rect 35023 25412 35035 25415
rect 35894 25412 35900 25424
rect 35023 25384 35900 25412
rect 35023 25381 35035 25384
rect 34977 25375 35035 25381
rect 35894 25372 35900 25384
rect 35952 25372 35958 25424
rect 37182 25372 37188 25424
rect 37240 25412 37246 25424
rect 38286 25412 38292 25424
rect 37240 25384 38292 25412
rect 37240 25372 37246 25384
rect 38286 25372 38292 25384
rect 38344 25412 38350 25424
rect 41782 25412 41788 25424
rect 38344 25384 39252 25412
rect 41743 25384 41788 25412
rect 38344 25372 38350 25384
rect 33832 25347 33890 25353
rect 33832 25313 33844 25347
rect 33878 25344 33890 25347
rect 34238 25344 34244 25356
rect 33878 25316 34244 25344
rect 33878 25313 33890 25316
rect 33832 25307 33890 25313
rect 34238 25304 34244 25316
rect 34296 25304 34302 25356
rect 36262 25304 36268 25356
rect 36320 25344 36326 25356
rect 36392 25347 36450 25353
rect 36392 25344 36404 25347
rect 36320 25316 36404 25344
rect 36320 25304 36326 25316
rect 36392 25313 36404 25316
rect 36438 25313 36450 25347
rect 36392 25307 36450 25313
rect 37645 25347 37703 25353
rect 37645 25313 37657 25347
rect 37691 25344 37703 25347
rect 37826 25344 37832 25356
rect 37691 25316 37832 25344
rect 37691 25313 37703 25316
rect 37645 25307 37703 25313
rect 37826 25304 37832 25316
rect 37884 25304 37890 25356
rect 39224 25353 39252 25384
rect 41782 25372 41788 25384
rect 41840 25372 41846 25424
rect 43530 25412 43536 25424
rect 43491 25384 43536 25412
rect 43530 25372 43536 25384
rect 43588 25372 43594 25424
rect 45373 25415 45431 25421
rect 45373 25381 45385 25415
rect 45419 25412 45431 25415
rect 46290 25412 46296 25424
rect 45419 25384 46296 25412
rect 45419 25381 45431 25384
rect 45373 25375 45431 25381
rect 46290 25372 46296 25384
rect 46348 25372 46354 25424
rect 39209 25347 39267 25353
rect 39209 25313 39221 25347
rect 39255 25344 39267 25347
rect 39298 25344 39304 25356
rect 39255 25316 39304 25344
rect 39255 25313 39267 25316
rect 39209 25307 39267 25313
rect 39298 25304 39304 25316
rect 39356 25304 39362 25356
rect 39390 25304 39396 25356
rect 39448 25344 39454 25356
rect 39669 25347 39727 25353
rect 39669 25344 39681 25347
rect 39448 25316 39681 25344
rect 39448 25304 39454 25316
rect 39669 25313 39681 25316
rect 39715 25313 39727 25347
rect 39669 25307 39727 25313
rect 32217 25279 32275 25285
rect 32217 25276 32229 25279
rect 31864 25248 32229 25276
rect 30837 25239 30895 25245
rect 32217 25245 32229 25248
rect 32263 25245 32275 25279
rect 32490 25276 32496 25288
rect 32451 25248 32496 25276
rect 32217 25239 32275 25245
rect 16114 25168 16120 25220
rect 16172 25208 16178 25220
rect 16853 25211 16911 25217
rect 16853 25208 16865 25211
rect 16172 25180 16865 25208
rect 16172 25168 16178 25180
rect 16853 25177 16865 25180
rect 16899 25177 16911 25211
rect 30392 25208 30420 25236
rect 30852 25208 30880 25239
rect 32490 25236 32496 25248
rect 32548 25236 32554 25288
rect 33919 25279 33977 25285
rect 33919 25245 33931 25279
rect 33965 25276 33977 25279
rect 34885 25279 34943 25285
rect 34885 25276 34897 25279
rect 33965 25248 34897 25276
rect 33965 25245 33977 25248
rect 33919 25239 33977 25245
rect 34885 25245 34897 25248
rect 34931 25276 34943 25279
rect 35526 25276 35532 25288
rect 34931 25248 35532 25276
rect 34931 25245 34943 25248
rect 34885 25239 34943 25245
rect 35526 25236 35532 25248
rect 35584 25236 35590 25288
rect 38102 25236 38108 25288
rect 38160 25276 38166 25288
rect 38289 25279 38347 25285
rect 38289 25276 38301 25279
rect 38160 25248 38301 25276
rect 38160 25236 38166 25248
rect 38289 25245 38301 25248
rect 38335 25276 38347 25279
rect 38470 25276 38476 25288
rect 38335 25248 38476 25276
rect 38335 25245 38347 25248
rect 38289 25239 38347 25245
rect 38470 25236 38476 25248
rect 38528 25236 38534 25288
rect 39942 25276 39948 25288
rect 39903 25248 39948 25276
rect 39942 25236 39948 25248
rect 40000 25236 40006 25288
rect 41509 25279 41567 25285
rect 41509 25245 41521 25279
rect 41555 25276 41567 25279
rect 41690 25276 41696 25288
rect 41555 25248 41696 25276
rect 41555 25245 41567 25248
rect 41509 25239 41567 25245
rect 41690 25236 41696 25248
rect 41748 25236 41754 25288
rect 41966 25276 41972 25288
rect 41927 25248 41972 25276
rect 41966 25236 41972 25248
rect 42024 25276 42030 25288
rect 43438 25276 43444 25288
rect 42024 25248 42794 25276
rect 43399 25248 43444 25276
rect 42024 25236 42030 25248
rect 35434 25208 35440 25220
rect 30392 25180 30880 25208
rect 35395 25180 35440 25208
rect 16853 25171 16911 25177
rect 35434 25168 35440 25180
rect 35492 25168 35498 25220
rect 37875 25211 37933 25217
rect 37875 25177 37887 25211
rect 37921 25208 37933 25211
rect 38378 25208 38384 25220
rect 37921 25180 38384 25208
rect 37921 25177 37933 25180
rect 37875 25171 37933 25177
rect 38378 25168 38384 25180
rect 38436 25208 38442 25220
rect 38565 25211 38623 25217
rect 38565 25208 38577 25211
rect 38436 25180 38577 25208
rect 38436 25168 38442 25180
rect 38565 25177 38577 25180
rect 38611 25177 38623 25211
rect 42766 25208 42794 25248
rect 43438 25236 43444 25248
rect 43496 25236 43502 25288
rect 43717 25279 43775 25285
rect 43717 25245 43729 25279
rect 43763 25245 43775 25279
rect 45278 25276 45284 25288
rect 45239 25248 45284 25276
rect 43717 25239 43775 25245
rect 43622 25208 43628 25220
rect 42766 25180 43628 25208
rect 38565 25171 38623 25177
rect 43622 25168 43628 25180
rect 43680 25208 43686 25220
rect 43732 25208 43760 25239
rect 45278 25236 45284 25248
rect 45336 25236 45342 25288
rect 45554 25276 45560 25288
rect 45515 25248 45560 25276
rect 45554 25236 45560 25248
rect 45612 25236 45618 25288
rect 46198 25236 46204 25288
rect 46256 25276 46262 25288
rect 46753 25279 46811 25285
rect 46753 25276 46765 25279
rect 46256 25248 46765 25276
rect 46256 25236 46262 25248
rect 46753 25245 46765 25248
rect 46799 25245 46811 25279
rect 46753 25239 46811 25245
rect 43680 25180 43760 25208
rect 43680 25168 43686 25180
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16298 25140 16304 25152
rect 16255 25112 16304 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 18414 25140 18420 25152
rect 18375 25112 18420 25140
rect 18414 25100 18420 25112
rect 18472 25100 18478 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20349 25143 20407 25149
rect 20349 25140 20361 25143
rect 20036 25112 20361 25140
rect 20036 25100 20042 25112
rect 20349 25109 20361 25112
rect 20395 25109 20407 25143
rect 27430 25140 27436 25152
rect 27391 25112 27436 25140
rect 20349 25103 20407 25109
rect 27430 25100 27436 25112
rect 27488 25100 27494 25152
rect 30650 25100 30656 25152
rect 30708 25140 30714 25152
rect 32306 25140 32312 25152
rect 30708 25112 32312 25140
rect 30708 25100 30714 25112
rect 32306 25100 32312 25112
rect 32364 25100 32370 25152
rect 36906 25140 36912 25152
rect 36867 25112 36912 25140
rect 36906 25100 36912 25112
rect 36964 25100 36970 25152
rect 44542 25140 44548 25152
rect 44503 25112 44548 25140
rect 44542 25100 44548 25112
rect 44600 25100 44606 25152
rect 46290 25140 46296 25152
rect 46251 25112 46296 25140
rect 46290 25100 46296 25112
rect 46348 25100 46354 25152
rect 1104 25050 48852 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 48852 25050
rect 1104 24976 48852 24998
rect 14918 24936 14924 24948
rect 14879 24908 14924 24936
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 17126 24936 17132 24948
rect 17087 24908 17132 24936
rect 17126 24896 17132 24908
rect 17184 24896 17190 24948
rect 17402 24936 17408 24948
rect 17363 24908 17408 24936
rect 17402 24896 17408 24908
rect 17460 24936 17466 24948
rect 18598 24936 18604 24948
rect 17460 24908 18604 24936
rect 17460 24896 17466 24908
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 18690 24896 18696 24948
rect 18748 24936 18754 24948
rect 19337 24939 19395 24945
rect 19337 24936 19349 24939
rect 18748 24908 19349 24936
rect 18748 24896 18754 24908
rect 19337 24905 19349 24908
rect 19383 24905 19395 24939
rect 19337 24899 19395 24905
rect 19797 24939 19855 24945
rect 19797 24905 19809 24939
rect 19843 24936 19855 24939
rect 19886 24936 19892 24948
rect 19843 24908 19892 24936
rect 19843 24905 19855 24908
rect 19797 24899 19855 24905
rect 19886 24896 19892 24908
rect 19944 24936 19950 24948
rect 20070 24936 20076 24948
rect 19944 24908 20076 24936
rect 19944 24896 19950 24908
rect 20070 24896 20076 24908
rect 20128 24896 20134 24948
rect 23290 24896 23296 24948
rect 23348 24936 23354 24948
rect 23385 24939 23443 24945
rect 23385 24936 23397 24939
rect 23348 24908 23397 24936
rect 23348 24896 23354 24908
rect 23385 24905 23397 24908
rect 23431 24905 23443 24939
rect 25130 24936 25136 24948
rect 25091 24908 25136 24936
rect 23385 24899 23443 24905
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 26510 24896 26516 24948
rect 26568 24936 26574 24948
rect 28077 24939 28135 24945
rect 28077 24936 28089 24939
rect 26568 24908 28089 24936
rect 26568 24896 26574 24908
rect 28077 24905 28089 24908
rect 28123 24905 28135 24939
rect 28077 24899 28135 24905
rect 28813 24939 28871 24945
rect 28813 24905 28825 24939
rect 28859 24936 28871 24939
rect 28902 24936 28908 24948
rect 28859 24908 28908 24936
rect 28859 24905 28871 24908
rect 28813 24899 28871 24905
rect 28902 24896 28908 24908
rect 28960 24896 28966 24948
rect 30650 24896 30656 24948
rect 30708 24936 30714 24948
rect 31021 24939 31079 24945
rect 31021 24936 31033 24939
rect 30708 24908 31033 24936
rect 30708 24896 30714 24908
rect 31021 24905 31033 24908
rect 31067 24905 31079 24939
rect 31021 24899 31079 24905
rect 31110 24896 31116 24948
rect 31168 24936 31174 24948
rect 31297 24939 31355 24945
rect 31297 24936 31309 24939
rect 31168 24908 31309 24936
rect 31168 24896 31174 24908
rect 31297 24905 31309 24908
rect 31343 24936 31355 24939
rect 31389 24939 31447 24945
rect 31389 24936 31401 24939
rect 31343 24908 31401 24936
rect 31343 24905 31355 24908
rect 31297 24899 31355 24905
rect 31389 24905 31401 24908
rect 31435 24905 31447 24939
rect 31389 24899 31447 24905
rect 32306 24896 32312 24948
rect 32364 24936 32370 24948
rect 32585 24939 32643 24945
rect 32585 24936 32597 24939
rect 32364 24908 32597 24936
rect 32364 24896 32370 24908
rect 32585 24905 32597 24908
rect 32631 24936 32643 24939
rect 32953 24939 33011 24945
rect 32953 24936 32965 24939
rect 32631 24908 32965 24936
rect 32631 24905 32643 24908
rect 32585 24899 32643 24905
rect 32953 24905 32965 24908
rect 32999 24936 33011 24939
rect 33318 24936 33324 24948
rect 32999 24908 33324 24936
rect 32999 24905 33011 24908
rect 32953 24899 33011 24905
rect 33318 24896 33324 24908
rect 33376 24896 33382 24948
rect 34606 24936 34612 24948
rect 34567 24908 34612 24936
rect 34606 24896 34612 24908
rect 34664 24896 34670 24948
rect 37826 24936 37832 24948
rect 37787 24908 37832 24936
rect 37826 24896 37832 24908
rect 37884 24896 37890 24948
rect 39298 24936 39304 24948
rect 39259 24908 39304 24936
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 39390 24896 39396 24948
rect 39448 24936 39454 24948
rect 39669 24939 39727 24945
rect 39669 24936 39681 24939
rect 39448 24908 39681 24936
rect 39448 24896 39454 24908
rect 39669 24905 39681 24908
rect 39715 24905 39727 24939
rect 39669 24899 39727 24905
rect 43438 24896 43444 24948
rect 43496 24936 43502 24948
rect 43901 24939 43959 24945
rect 43901 24936 43913 24939
rect 43496 24908 43913 24936
rect 43496 24896 43502 24908
rect 43901 24905 43913 24908
rect 43947 24936 43959 24939
rect 45554 24936 45560 24948
rect 43947 24908 45560 24936
rect 43947 24905 43959 24908
rect 43901 24899 43959 24905
rect 45554 24896 45560 24908
rect 45612 24896 45618 24948
rect 16669 24871 16727 24877
rect 16669 24837 16681 24871
rect 16715 24868 16727 24871
rect 16758 24868 16764 24880
rect 16715 24840 16764 24868
rect 16715 24837 16727 24840
rect 16669 24831 16727 24837
rect 16758 24828 16764 24840
rect 16816 24868 16822 24880
rect 17862 24868 17868 24880
rect 16816 24840 17868 24868
rect 16816 24828 16822 24840
rect 17862 24828 17868 24840
rect 17920 24868 17926 24880
rect 18874 24868 18880 24880
rect 17920 24840 18880 24868
rect 17920 24828 17926 24840
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 24857 24871 24915 24877
rect 23446 24840 24808 24868
rect 15151 24803 15209 24809
rect 15151 24769 15163 24803
rect 15197 24800 15209 24803
rect 17773 24803 17831 24809
rect 17773 24800 17785 24803
rect 15197 24772 17785 24800
rect 15197 24769 15209 24772
rect 15151 24763 15209 24769
rect 17773 24769 17785 24772
rect 17819 24800 17831 24803
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 17819 24772 18429 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 18598 24760 18604 24812
rect 18656 24800 18662 24812
rect 18693 24803 18751 24809
rect 18693 24800 18705 24803
rect 18656 24772 18705 24800
rect 18656 24760 18662 24772
rect 18693 24769 18705 24772
rect 18739 24800 18751 24803
rect 19150 24800 19156 24812
rect 18739 24772 19156 24800
rect 18739 24769 18751 24772
rect 18693 24763 18751 24769
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 22370 24800 22376 24812
rect 22331 24772 22376 24800
rect 22370 24760 22376 24772
rect 22428 24800 22434 24812
rect 23446 24800 23474 24840
rect 23750 24800 23756 24812
rect 22428 24772 23474 24800
rect 23711 24772 23756 24800
rect 22428 24760 22434 24772
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 23934 24760 23940 24812
rect 23992 24800 23998 24812
rect 24029 24803 24087 24809
rect 24029 24800 24041 24803
rect 23992 24772 24041 24800
rect 23992 24760 23998 24772
rect 24029 24769 24041 24772
rect 24075 24769 24087 24803
rect 24029 24763 24087 24769
rect 15064 24735 15122 24741
rect 15064 24701 15076 24735
rect 15110 24732 15122 24735
rect 24780 24732 24808 24840
rect 24857 24837 24869 24871
rect 24903 24868 24915 24871
rect 25038 24868 25044 24880
rect 24903 24840 25044 24868
rect 24903 24837 24915 24840
rect 24857 24831 24915 24837
rect 25038 24828 25044 24840
rect 25096 24868 25102 24880
rect 26237 24871 26295 24877
rect 26237 24868 26249 24871
rect 25096 24840 26249 24868
rect 25096 24828 25102 24840
rect 26237 24837 26249 24840
rect 26283 24837 26295 24871
rect 26237 24831 26295 24837
rect 30006 24828 30012 24880
rect 30064 24868 30070 24880
rect 32217 24871 32275 24877
rect 32217 24868 32229 24871
rect 30064 24840 32229 24868
rect 30064 24828 30070 24840
rect 32217 24837 32229 24840
rect 32263 24868 32275 24871
rect 32490 24868 32496 24880
rect 32263 24840 32496 24868
rect 32263 24837 32275 24840
rect 32217 24831 32275 24837
rect 32490 24828 32496 24840
rect 32548 24828 32554 24880
rect 32674 24828 32680 24880
rect 32732 24868 32738 24880
rect 36262 24868 36268 24880
rect 32732 24840 36268 24868
rect 32732 24828 32738 24840
rect 36262 24828 36268 24840
rect 36320 24868 36326 24880
rect 36357 24871 36415 24877
rect 36357 24868 36369 24871
rect 36320 24840 36369 24868
rect 36320 24828 36326 24840
rect 36357 24837 36369 24840
rect 36403 24868 36415 24871
rect 39206 24868 39212 24880
rect 36403 24840 39212 24868
rect 36403 24837 36415 24840
rect 36357 24831 36415 24837
rect 39206 24828 39212 24840
rect 39264 24828 39270 24880
rect 40313 24871 40371 24877
rect 40313 24837 40325 24871
rect 40359 24868 40371 24871
rect 43990 24868 43996 24880
rect 40359 24840 43996 24868
rect 40359 24837 40371 24840
rect 40313 24831 40371 24837
rect 25314 24800 25320 24812
rect 25275 24772 25320 24800
rect 25314 24760 25320 24772
rect 25372 24760 25378 24812
rect 25590 24760 25596 24812
rect 25648 24800 25654 24812
rect 27246 24800 27252 24812
rect 25648 24772 27252 24800
rect 25648 24760 25654 24772
rect 27246 24760 27252 24772
rect 27304 24800 27310 24812
rect 27433 24803 27491 24809
rect 27433 24800 27445 24803
rect 27304 24772 27445 24800
rect 27304 24760 27310 24772
rect 27433 24769 27445 24772
rect 27479 24769 27491 24803
rect 30374 24800 30380 24812
rect 30335 24772 30380 24800
rect 27433 24763 27491 24769
rect 30374 24760 30380 24772
rect 30432 24760 30438 24812
rect 31662 24800 31668 24812
rect 31575 24772 31668 24800
rect 31662 24760 31668 24772
rect 31720 24800 31726 24812
rect 32122 24800 32128 24812
rect 31720 24772 32128 24800
rect 31720 24760 31726 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 33226 24800 33232 24812
rect 33187 24772 33232 24800
rect 33226 24760 33232 24772
rect 33284 24760 33290 24812
rect 33502 24800 33508 24812
rect 33463 24772 33508 24800
rect 33502 24760 33508 24772
rect 33560 24760 33566 24812
rect 34790 24760 34796 24812
rect 34848 24800 34854 24812
rect 34977 24803 35035 24809
rect 34977 24800 34989 24803
rect 34848 24772 34989 24800
rect 34848 24760 34854 24772
rect 34977 24769 34989 24772
rect 35023 24769 35035 24803
rect 35434 24800 35440 24812
rect 35395 24772 35440 24800
rect 34977 24763 35035 24769
rect 35434 24760 35440 24772
rect 35492 24760 35498 24812
rect 37458 24800 37464 24812
rect 37419 24772 37464 24800
rect 37458 24760 37464 24772
rect 37516 24800 37522 24812
rect 37642 24800 37648 24812
rect 37516 24772 37648 24800
rect 37516 24760 37522 24772
rect 37642 24760 37648 24772
rect 37700 24760 37706 24812
rect 38378 24800 38384 24812
rect 38339 24772 38384 24800
rect 38378 24760 38384 24772
rect 38436 24760 38442 24812
rect 38470 24760 38476 24812
rect 38528 24800 38534 24812
rect 40880 24809 40908 24840
rect 43990 24828 43996 24840
rect 44048 24868 44054 24880
rect 46750 24868 46756 24880
rect 44048 24840 44864 24868
rect 46711 24840 46756 24868
rect 44048 24828 44054 24840
rect 38657 24803 38715 24809
rect 38657 24800 38669 24803
rect 38528 24772 38669 24800
rect 38528 24760 38534 24772
rect 38657 24769 38669 24772
rect 38703 24769 38715 24803
rect 38657 24763 38715 24769
rect 40865 24803 40923 24809
rect 40865 24769 40877 24803
rect 40911 24769 40923 24803
rect 40865 24763 40923 24769
rect 41509 24803 41567 24809
rect 41509 24769 41521 24803
rect 41555 24800 41567 24803
rect 41966 24800 41972 24812
rect 41555 24772 41972 24800
rect 41555 24769 41567 24772
rect 41509 24763 41567 24769
rect 41966 24760 41972 24772
rect 42024 24760 42030 24812
rect 44542 24800 44548 24812
rect 44503 24772 44548 24800
rect 44542 24760 44548 24772
rect 44600 24760 44606 24812
rect 44836 24809 44864 24840
rect 46750 24828 46756 24840
rect 46808 24828 46814 24880
rect 44821 24803 44879 24809
rect 44821 24769 44833 24803
rect 44867 24769 44879 24803
rect 44821 24763 44879 24769
rect 45925 24803 45983 24809
rect 45925 24769 45937 24803
rect 45971 24800 45983 24803
rect 46198 24800 46204 24812
rect 45971 24772 46204 24800
rect 45971 24769 45983 24772
rect 45925 24763 45983 24769
rect 46198 24760 46204 24772
rect 46256 24760 46262 24812
rect 42337 24735 42395 24741
rect 15110 24704 15976 24732
rect 24780 24704 26372 24732
rect 15110 24701 15122 24704
rect 15064 24695 15122 24701
rect 15470 24596 15476 24608
rect 15431 24568 15476 24596
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15948 24605 15976 24704
rect 16114 24664 16120 24676
rect 16075 24636 16120 24664
rect 16114 24624 16120 24636
rect 16172 24624 16178 24676
rect 16206 24624 16212 24676
rect 16264 24664 16270 24676
rect 16264 24636 16309 24664
rect 16264 24624 16270 24636
rect 18414 24624 18420 24676
rect 18472 24664 18478 24676
rect 18509 24667 18567 24673
rect 18509 24664 18521 24667
rect 18472 24636 18521 24664
rect 18472 24624 18478 24636
rect 18509 24633 18521 24636
rect 18555 24664 18567 24667
rect 19334 24664 19340 24676
rect 18555 24636 19340 24664
rect 18555 24633 18567 24636
rect 18509 24627 18567 24633
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 19978 24664 19984 24676
rect 19438 24636 19984 24664
rect 15933 24599 15991 24605
rect 15933 24565 15945 24599
rect 15979 24596 15991 24599
rect 16022 24596 16028 24608
rect 15979 24568 16028 24596
rect 15979 24565 15991 24568
rect 15933 24559 15991 24565
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 18138 24556 18144 24608
rect 18196 24596 18202 24608
rect 19438 24596 19466 24636
rect 19978 24624 19984 24636
rect 20036 24624 20042 24676
rect 20070 24624 20076 24676
rect 20128 24664 20134 24676
rect 20622 24664 20628 24676
rect 20128 24636 20173 24664
rect 20583 24636 20628 24664
rect 20128 24624 20134 24636
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 21269 24667 21327 24673
rect 21269 24633 21281 24667
rect 21315 24664 21327 24667
rect 21450 24664 21456 24676
rect 21315 24636 21456 24664
rect 21315 24633 21327 24636
rect 21269 24627 21327 24633
rect 21450 24624 21456 24636
rect 21508 24664 21514 24676
rect 22097 24667 22155 24673
rect 22097 24664 22109 24667
rect 21508 24636 22109 24664
rect 21508 24624 21514 24636
rect 22097 24633 22109 24636
rect 22143 24633 22155 24667
rect 22097 24627 22155 24633
rect 22186 24624 22192 24676
rect 22244 24664 22250 24676
rect 22244 24636 22289 24664
rect 22244 24624 22250 24636
rect 23290 24624 23296 24676
rect 23348 24664 23354 24676
rect 23845 24667 23903 24673
rect 23348 24636 23474 24664
rect 23348 24624 23354 24636
rect 21542 24596 21548 24608
rect 18196 24568 19466 24596
rect 21503 24568 21548 24596
rect 18196 24556 18202 24568
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 22204 24596 22232 24624
rect 23017 24599 23075 24605
rect 23017 24596 23029 24599
rect 22204 24568 23029 24596
rect 23017 24565 23029 24568
rect 23063 24565 23075 24599
rect 23446 24596 23474 24636
rect 23845 24633 23857 24667
rect 23891 24633 23903 24667
rect 23845 24627 23903 24633
rect 23860 24596 23888 24627
rect 25130 24624 25136 24676
rect 25188 24664 25194 24676
rect 25638 24667 25696 24673
rect 25638 24664 25650 24667
rect 25188 24636 25650 24664
rect 25188 24624 25194 24636
rect 25638 24633 25650 24636
rect 25684 24633 25696 24667
rect 26344 24664 26372 24704
rect 42337 24701 42349 24735
rect 42383 24732 42395 24735
rect 42426 24732 42432 24744
rect 42383 24704 42432 24732
rect 42383 24701 42395 24704
rect 42337 24695 42395 24701
rect 42426 24692 42432 24704
rect 42484 24692 42490 24744
rect 27154 24664 27160 24676
rect 26344 24636 27160 24664
rect 25638 24627 25696 24633
rect 23446 24568 23888 24596
rect 25653 24596 25681 24627
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 27249 24667 27307 24673
rect 27249 24633 27261 24667
rect 27295 24664 27307 24667
rect 27430 24664 27436 24676
rect 27295 24636 27436 24664
rect 27295 24633 27307 24636
rect 27249 24627 27307 24633
rect 26513 24599 26571 24605
rect 26513 24596 26525 24599
rect 25653 24568 26525 24596
rect 23017 24559 23075 24565
rect 26513 24565 26525 24568
rect 26559 24596 26571 24599
rect 26878 24596 26884 24608
rect 26559 24568 26884 24596
rect 26559 24565 26571 24568
rect 26513 24559 26571 24565
rect 26878 24556 26884 24568
rect 26936 24556 26942 24608
rect 26973 24599 27031 24605
rect 26973 24565 26985 24599
rect 27019 24596 27031 24599
rect 27264 24596 27292 24627
rect 27430 24624 27436 24636
rect 27488 24624 27494 24676
rect 29549 24667 29607 24673
rect 29549 24633 29561 24667
rect 29595 24664 29607 24667
rect 30098 24664 30104 24676
rect 29595 24636 30104 24664
rect 29595 24633 29607 24636
rect 29549 24627 29607 24633
rect 30098 24624 30104 24636
rect 30156 24624 30162 24676
rect 30193 24667 30251 24673
rect 30193 24633 30205 24667
rect 30239 24664 30251 24667
rect 31297 24667 31355 24673
rect 31297 24664 31309 24667
rect 30239 24636 31309 24664
rect 30239 24633 30251 24636
rect 30193 24627 30251 24633
rect 31297 24633 31309 24636
rect 31343 24664 31355 24667
rect 31757 24667 31815 24673
rect 31757 24664 31769 24667
rect 31343 24636 31769 24664
rect 31343 24633 31355 24636
rect 31297 24627 31355 24633
rect 31757 24633 31769 24636
rect 31803 24664 31815 24667
rect 32306 24664 32312 24676
rect 31803 24636 32312 24664
rect 31803 24633 31815 24636
rect 31757 24627 31815 24633
rect 27019 24568 27292 24596
rect 29917 24599 29975 24605
rect 27019 24565 27031 24568
rect 26973 24559 27031 24565
rect 29917 24565 29929 24599
rect 29963 24596 29975 24599
rect 30208 24596 30236 24627
rect 32306 24624 32312 24636
rect 32364 24624 32370 24676
rect 33318 24664 33324 24676
rect 33279 24636 33324 24664
rect 33318 24624 33324 24636
rect 33376 24624 33382 24676
rect 34238 24664 34244 24676
rect 34199 24636 34244 24664
rect 34238 24624 34244 24636
rect 34296 24624 34302 24676
rect 35069 24667 35127 24673
rect 35069 24633 35081 24667
rect 35115 24664 35127 24667
rect 35986 24664 35992 24676
rect 35115 24636 35992 24664
rect 35115 24633 35127 24636
rect 35069 24627 35127 24633
rect 35986 24624 35992 24636
rect 36044 24664 36050 24676
rect 36044 24636 36492 24664
rect 36044 24624 36050 24636
rect 29963 24568 30236 24596
rect 36464 24596 36492 24636
rect 36630 24624 36636 24676
rect 36688 24664 36694 24676
rect 36817 24667 36875 24673
rect 36817 24664 36829 24667
rect 36688 24636 36829 24664
rect 36688 24624 36694 24636
rect 36817 24633 36829 24636
rect 36863 24633 36875 24667
rect 36817 24627 36875 24633
rect 36906 24624 36912 24676
rect 36964 24664 36970 24676
rect 38197 24667 38255 24673
rect 38197 24664 38209 24667
rect 36964 24636 37009 24664
rect 37108 24636 38209 24664
rect 36964 24624 36970 24636
rect 37108 24596 37136 24636
rect 38197 24633 38209 24636
rect 38243 24664 38255 24667
rect 38473 24667 38531 24673
rect 38473 24664 38485 24667
rect 38243 24636 38485 24664
rect 38243 24633 38255 24636
rect 38197 24627 38255 24633
rect 38473 24633 38485 24636
rect 38519 24633 38531 24667
rect 38473 24627 38531 24633
rect 40954 24624 40960 24676
rect 41012 24664 41018 24676
rect 42658 24667 42716 24673
rect 42658 24664 42670 24667
rect 41012 24636 41057 24664
rect 42168 24636 42670 24664
rect 41012 24624 41018 24636
rect 41782 24596 41788 24608
rect 36464 24568 37136 24596
rect 41743 24568 41788 24596
rect 29963 24565 29975 24568
rect 29917 24559 29975 24565
rect 41782 24556 41788 24568
rect 41840 24556 41846 24608
rect 42058 24556 42064 24608
rect 42116 24596 42122 24608
rect 42168 24605 42196 24636
rect 42658 24633 42670 24636
rect 42704 24633 42716 24667
rect 42658 24627 42716 24633
rect 44637 24667 44695 24673
rect 44637 24633 44649 24667
rect 44683 24633 44695 24667
rect 44637 24627 44695 24633
rect 45557 24667 45615 24673
rect 45557 24633 45569 24667
rect 45603 24664 45615 24667
rect 46290 24664 46296 24676
rect 45603 24636 46296 24664
rect 45603 24633 45615 24636
rect 45557 24627 45615 24633
rect 42153 24599 42211 24605
rect 42153 24596 42165 24599
rect 42116 24568 42165 24596
rect 42116 24556 42122 24568
rect 42153 24565 42165 24568
rect 42199 24565 42211 24599
rect 43254 24596 43260 24608
rect 43215 24568 43260 24596
rect 42153 24559 42211 24565
rect 43254 24556 43260 24568
rect 43312 24556 43318 24608
rect 43530 24596 43536 24608
rect 43491 24568 43536 24596
rect 43530 24556 43536 24568
rect 43588 24556 43594 24608
rect 44361 24599 44419 24605
rect 44361 24565 44373 24599
rect 44407 24596 44419 24599
rect 44652 24596 44680 24627
rect 45572 24596 45600 24627
rect 46290 24624 46296 24636
rect 46348 24624 46354 24676
rect 44407 24568 45600 24596
rect 44407 24565 44419 24568
rect 44361 24559 44419 24565
rect 1104 24506 48852 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 48852 24506
rect 1104 24432 48852 24454
rect 14323 24395 14381 24401
rect 14323 24361 14335 24395
rect 14369 24392 14381 24395
rect 18138 24392 18144 24404
rect 14369 24364 18144 24392
rect 14369 24361 14381 24364
rect 14323 24355 14381 24361
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 18230 24352 18236 24404
rect 18288 24392 18294 24404
rect 18693 24395 18751 24401
rect 18693 24392 18705 24395
rect 18288 24364 18705 24392
rect 18288 24352 18294 24364
rect 18693 24361 18705 24364
rect 18739 24392 18751 24395
rect 18966 24392 18972 24404
rect 18739 24364 18972 24392
rect 18739 24361 18751 24364
rect 18693 24355 18751 24361
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 19058 24352 19064 24404
rect 19116 24352 19122 24404
rect 22462 24392 22468 24404
rect 21836 24364 22468 24392
rect 16209 24327 16267 24333
rect 16209 24293 16221 24327
rect 16255 24324 16267 24327
rect 16298 24324 16304 24336
rect 16255 24296 16304 24324
rect 16255 24293 16267 24296
rect 16209 24287 16267 24293
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 16758 24324 16764 24336
rect 16719 24296 16764 24324
rect 16758 24284 16764 24296
rect 16816 24284 16822 24336
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 18192 24259 18250 24265
rect 18192 24256 18204 24259
rect 17920 24228 18204 24256
rect 17920 24216 17926 24228
rect 18192 24225 18204 24228
rect 18238 24256 18250 24259
rect 19076 24256 19104 24352
rect 21836 24336 21864 24364
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 22646 24352 22652 24404
rect 22704 24392 22710 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22704 24364 22753 24392
rect 22704 24352 22710 24364
rect 22741 24361 22753 24364
rect 22787 24361 22799 24395
rect 22741 24355 22799 24361
rect 25314 24352 25320 24404
rect 25372 24392 25378 24404
rect 25869 24395 25927 24401
rect 25869 24392 25881 24395
rect 25372 24364 25881 24392
rect 25372 24352 25378 24364
rect 25869 24361 25881 24364
rect 25915 24361 25927 24395
rect 25869 24355 25927 24361
rect 27154 24352 27160 24404
rect 27212 24392 27218 24404
rect 27525 24395 27583 24401
rect 27525 24392 27537 24395
rect 27212 24364 27537 24392
rect 27212 24352 27218 24364
rect 27525 24361 27537 24364
rect 27571 24361 27583 24395
rect 28534 24392 28540 24404
rect 28495 24364 28540 24392
rect 27525 24355 27583 24361
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 28810 24352 28816 24404
rect 28868 24392 28874 24404
rect 29365 24395 29423 24401
rect 29365 24392 29377 24395
rect 28868 24364 29377 24392
rect 28868 24352 28874 24364
rect 29365 24361 29377 24364
rect 29411 24361 29423 24395
rect 29365 24355 29423 24361
rect 30147 24395 30205 24401
rect 30147 24361 30159 24395
rect 30193 24392 30205 24395
rect 30558 24392 30564 24404
rect 30193 24364 30564 24392
rect 30193 24361 30205 24364
rect 30147 24355 30205 24361
rect 30558 24352 30564 24364
rect 30616 24352 30622 24404
rect 31662 24392 31668 24404
rect 31623 24364 31668 24392
rect 31662 24352 31668 24364
rect 31720 24352 31726 24404
rect 33226 24392 33232 24404
rect 33187 24364 33232 24392
rect 33226 24352 33232 24364
rect 33284 24352 33290 24404
rect 35526 24392 35532 24404
rect 35487 24364 35532 24392
rect 35526 24352 35532 24364
rect 35584 24352 35590 24404
rect 40405 24395 40463 24401
rect 40405 24361 40417 24395
rect 40451 24392 40463 24395
rect 41782 24392 41788 24404
rect 40451 24364 41788 24392
rect 40451 24361 40463 24364
rect 40405 24355 40463 24361
rect 41782 24352 41788 24364
rect 41840 24352 41846 24404
rect 42153 24395 42211 24401
rect 42153 24361 42165 24395
rect 42199 24392 42211 24395
rect 43530 24392 43536 24404
rect 42199 24364 43536 24392
rect 42199 24361 42211 24364
rect 42153 24355 42211 24361
rect 43530 24352 43536 24364
rect 43588 24352 43594 24404
rect 45189 24395 45247 24401
rect 45189 24361 45201 24395
rect 45235 24361 45247 24395
rect 45189 24355 45247 24361
rect 19334 24324 19340 24336
rect 19247 24296 19340 24324
rect 19334 24284 19340 24296
rect 19392 24324 19398 24336
rect 20070 24324 20076 24336
rect 19392 24296 20076 24324
rect 19392 24284 19398 24296
rect 20070 24284 20076 24296
rect 20128 24284 20134 24336
rect 21818 24324 21824 24336
rect 21731 24296 21824 24324
rect 21818 24284 21824 24296
rect 21876 24284 21882 24336
rect 21913 24327 21971 24333
rect 21913 24293 21925 24327
rect 21959 24324 21971 24327
rect 22186 24324 22192 24336
rect 21959 24296 22192 24324
rect 21959 24293 21971 24296
rect 21913 24287 21971 24293
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 23474 24284 23480 24336
rect 23532 24324 23538 24336
rect 25041 24327 25099 24333
rect 23532 24296 23577 24324
rect 23532 24284 23538 24296
rect 25041 24293 25053 24327
rect 25087 24324 25099 24327
rect 25406 24324 25412 24336
rect 25087 24296 25412 24324
rect 25087 24293 25099 24296
rect 25041 24287 25099 24293
rect 25406 24284 25412 24296
rect 25464 24284 25470 24336
rect 26694 24324 26700 24336
rect 26655 24296 26700 24324
rect 26694 24284 26700 24296
rect 26752 24284 26758 24336
rect 27246 24324 27252 24336
rect 27207 24296 27252 24324
rect 27246 24284 27252 24296
rect 27304 24284 27310 24336
rect 29270 24284 29276 24336
rect 29328 24324 29334 24336
rect 32214 24324 32220 24336
rect 29328 24296 32220 24324
rect 29328 24284 29334 24296
rect 32214 24284 32220 24296
rect 32272 24284 32278 24336
rect 32306 24284 32312 24336
rect 32364 24324 32370 24336
rect 32861 24327 32919 24333
rect 32364 24296 32409 24324
rect 32364 24284 32370 24296
rect 32861 24293 32873 24327
rect 32907 24324 32919 24327
rect 33502 24324 33508 24336
rect 32907 24296 33508 24324
rect 32907 24293 32919 24296
rect 32861 24287 32919 24293
rect 33502 24284 33508 24296
rect 33560 24284 33566 24336
rect 34514 24284 34520 24336
rect 34572 24324 34578 24336
rect 34654 24327 34712 24333
rect 34654 24324 34666 24327
rect 34572 24296 34666 24324
rect 34572 24284 34578 24296
rect 34654 24293 34666 24296
rect 34700 24293 34712 24327
rect 34654 24287 34712 24293
rect 35894 24284 35900 24336
rect 35952 24324 35958 24336
rect 36265 24327 36323 24333
rect 36265 24324 36277 24327
rect 35952 24296 36277 24324
rect 35952 24284 35958 24296
rect 36265 24293 36277 24296
rect 36311 24293 36323 24327
rect 36265 24287 36323 24293
rect 36446 24284 36452 24336
rect 36504 24324 36510 24336
rect 36504 24296 37044 24324
rect 36504 24284 36510 24296
rect 37016 24268 37044 24296
rect 39482 24284 39488 24336
rect 39540 24324 39546 24336
rect 39847 24327 39905 24333
rect 39847 24324 39859 24327
rect 39540 24296 39859 24324
rect 39540 24284 39546 24296
rect 39847 24293 39859 24296
rect 39893 24324 39905 24327
rect 40310 24324 40316 24336
rect 39893 24296 40316 24324
rect 39893 24293 39905 24296
rect 39847 24287 39905 24293
rect 40310 24284 40316 24296
rect 40368 24324 40374 24336
rect 41554 24327 41612 24333
rect 41554 24324 41566 24327
rect 40368 24296 41566 24324
rect 40368 24284 40374 24296
rect 41554 24293 41566 24296
rect 41600 24324 41612 24327
rect 42058 24324 42064 24336
rect 41600 24296 42064 24324
rect 41600 24293 41612 24296
rect 41554 24287 41612 24293
rect 42058 24284 42064 24296
rect 42116 24284 42122 24336
rect 44358 24284 44364 24336
rect 44416 24324 44422 24336
rect 44590 24327 44648 24333
rect 44590 24324 44602 24327
rect 44416 24296 44602 24324
rect 44416 24284 44422 24296
rect 44590 24293 44602 24296
rect 44636 24293 44648 24327
rect 45204 24324 45232 24355
rect 45278 24352 45284 24404
rect 45336 24392 45342 24404
rect 45462 24392 45468 24404
rect 45336 24364 45468 24392
rect 45336 24352 45342 24364
rect 45462 24352 45468 24364
rect 45520 24352 45526 24404
rect 45830 24324 45836 24336
rect 45204 24296 45836 24324
rect 44590 24287 44648 24293
rect 45830 24284 45836 24296
rect 45888 24324 45894 24336
rect 46201 24327 46259 24333
rect 46201 24324 46213 24327
rect 45888 24296 46213 24324
rect 45888 24284 45894 24296
rect 46201 24293 46213 24296
rect 46247 24324 46259 24327
rect 46290 24324 46296 24336
rect 46247 24296 46296 24324
rect 46247 24293 46259 24296
rect 46201 24287 46259 24293
rect 46290 24284 46296 24296
rect 46348 24284 46354 24336
rect 18238 24228 19104 24256
rect 18238 24225 18250 24228
rect 18192 24219 18250 24225
rect 27706 24216 27712 24268
rect 27764 24256 27770 24268
rect 30076 24259 30134 24265
rect 30076 24256 30088 24259
rect 27764 24228 30088 24256
rect 27764 24216 27770 24228
rect 30076 24225 30088 24228
rect 30122 24256 30134 24259
rect 30190 24256 30196 24268
rect 30122 24228 30196 24256
rect 30122 24225 30134 24228
rect 30076 24219 30134 24225
rect 30190 24216 30196 24228
rect 30248 24216 30254 24268
rect 31056 24259 31114 24265
rect 31056 24256 31068 24259
rect 30300 24228 31068 24256
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16117 24191 16175 24197
rect 16117 24188 16129 24191
rect 15979 24160 16129 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16117 24157 16129 24160
rect 16163 24188 16175 24191
rect 17034 24188 17040 24200
rect 16163 24160 17040 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 18279 24191 18337 24197
rect 18279 24157 18291 24191
rect 18325 24188 18337 24191
rect 19242 24188 19248 24200
rect 18325 24160 19248 24188
rect 18325 24157 18337 24160
rect 18279 24151 18337 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 19978 24188 19984 24200
rect 19935 24160 19984 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24188 22523 24191
rect 22738 24188 22744 24200
rect 22511 24160 22744 24188
rect 22511 24157 22523 24160
rect 22465 24151 22523 24157
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 23382 24188 23388 24200
rect 23343 24160 23388 24188
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 24946 24188 24952 24200
rect 24907 24160 24952 24188
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 16022 24080 16028 24132
rect 16080 24120 16086 24132
rect 20180 24120 20208 24148
rect 22922 24120 22928 24132
rect 16080 24092 22928 24120
rect 16080 24080 16086 24092
rect 22922 24080 22928 24092
rect 22980 24080 22986 24132
rect 23934 24120 23940 24132
rect 23895 24092 23940 24120
rect 23934 24080 23940 24092
rect 23992 24120 23998 24132
rect 24673 24123 24731 24129
rect 24673 24120 24685 24123
rect 23992 24092 24685 24120
rect 23992 24080 23998 24092
rect 24673 24089 24685 24092
rect 24719 24120 24731 24123
rect 25240 24120 25268 24151
rect 25866 24148 25872 24200
rect 25924 24188 25930 24200
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 25924 24160 26617 24188
rect 25924 24148 25930 24160
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 28166 24188 28172 24200
rect 28127 24160 28172 24188
rect 26605 24151 26663 24157
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 30300 24188 30328 24228
rect 31056 24225 31068 24228
rect 31102 24256 31114 24259
rect 31294 24256 31300 24268
rect 31102 24228 31300 24256
rect 31102 24225 31114 24228
rect 31056 24219 31114 24225
rect 31294 24216 31300 24228
rect 31352 24216 31358 24268
rect 33106 24228 35204 24256
rect 30069 24160 30328 24188
rect 24719 24092 25268 24120
rect 24719 24089 24731 24092
rect 24673 24083 24731 24089
rect 26326 24080 26332 24132
rect 26384 24120 26390 24132
rect 30069 24120 30097 24160
rect 26384 24092 30097 24120
rect 31159 24123 31217 24129
rect 26384 24080 26390 24092
rect 31159 24089 31171 24123
rect 31205 24120 31217 24123
rect 33106 24120 33134 24228
rect 34333 24191 34391 24197
rect 34333 24188 34345 24191
rect 31205 24092 33134 24120
rect 34164 24160 34345 24188
rect 31205 24089 31217 24092
rect 31159 24083 31217 24089
rect 18049 24055 18107 24061
rect 18049 24021 18061 24055
rect 18095 24052 18107 24055
rect 18138 24052 18144 24064
rect 18095 24024 18144 24052
rect 18095 24021 18107 24024
rect 18049 24015 18107 24021
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 20165 24055 20223 24061
rect 20165 24052 20177 24055
rect 19760 24024 20177 24052
rect 19760 24012 19766 24024
rect 20165 24021 20177 24024
rect 20211 24021 20223 24055
rect 29086 24052 29092 24064
rect 29047 24024 29092 24052
rect 20165 24015 20223 24021
rect 29086 24012 29092 24024
rect 29144 24012 29150 24064
rect 34054 24012 34060 24064
rect 34112 24052 34118 24064
rect 34164 24061 34192 24160
rect 34333 24157 34345 24160
rect 34379 24157 34391 24191
rect 35176 24188 35204 24228
rect 36998 24216 37004 24268
rect 37056 24256 37062 24268
rect 37918 24256 37924 24268
rect 37056 24228 37924 24256
rect 37056 24216 37062 24228
rect 37918 24216 37924 24228
rect 37976 24216 37982 24268
rect 38378 24216 38384 24268
rect 38436 24256 38442 24268
rect 38473 24259 38531 24265
rect 38473 24256 38485 24259
rect 38436 24228 38485 24256
rect 38436 24216 38442 24228
rect 38473 24225 38485 24228
rect 38519 24256 38531 24259
rect 39390 24256 39396 24268
rect 38519 24228 39396 24256
rect 38519 24225 38531 24228
rect 38473 24219 38531 24225
rect 39390 24216 39396 24228
rect 39448 24216 39454 24268
rect 36170 24188 36176 24200
rect 35176 24160 36176 24188
rect 34333 24151 34391 24157
rect 36170 24148 36176 24160
rect 36228 24148 36234 24200
rect 36630 24148 36636 24200
rect 36688 24188 36694 24200
rect 37093 24191 37151 24197
rect 37093 24188 37105 24191
rect 36688 24160 37105 24188
rect 36688 24148 36694 24160
rect 37093 24157 37105 24160
rect 37139 24157 37151 24191
rect 37093 24151 37151 24157
rect 38657 24191 38715 24197
rect 38657 24157 38669 24191
rect 38703 24188 38715 24191
rect 39482 24188 39488 24200
rect 38703 24160 39488 24188
rect 38703 24157 38715 24160
rect 38657 24151 38715 24157
rect 39482 24148 39488 24160
rect 39540 24148 39546 24200
rect 41230 24188 41236 24200
rect 41191 24160 41236 24188
rect 41230 24148 41236 24160
rect 41288 24148 41294 24200
rect 44266 24188 44272 24200
rect 44227 24160 44272 24188
rect 44266 24148 44272 24160
rect 44324 24148 44330 24200
rect 46106 24188 46112 24200
rect 46067 24160 46112 24188
rect 46106 24148 46112 24160
rect 46164 24148 46170 24200
rect 46474 24188 46480 24200
rect 46435 24160 46480 24188
rect 46474 24148 46480 24160
rect 46532 24148 46538 24200
rect 35250 24120 35256 24132
rect 35163 24092 35256 24120
rect 35250 24080 35256 24092
rect 35308 24120 35314 24132
rect 36725 24123 36783 24129
rect 35308 24092 36032 24120
rect 35308 24080 35314 24092
rect 34149 24055 34207 24061
rect 34149 24052 34161 24055
rect 34112 24024 34161 24052
rect 34112 24012 34118 24024
rect 34149 24021 34161 24024
rect 34195 24021 34207 24055
rect 35894 24052 35900 24064
rect 35855 24024 35900 24052
rect 34149 24015 34207 24021
rect 35894 24012 35900 24024
rect 35952 24012 35958 24064
rect 36004 24052 36032 24092
rect 36725 24089 36737 24123
rect 36771 24120 36783 24123
rect 37274 24120 37280 24132
rect 36771 24092 37280 24120
rect 36771 24089 36783 24092
rect 36725 24083 36783 24089
rect 37274 24080 37280 24092
rect 37332 24080 37338 24132
rect 36906 24052 36912 24064
rect 36004 24024 36912 24052
rect 36906 24012 36912 24024
rect 36964 24012 36970 24064
rect 40862 24052 40868 24064
rect 40823 24024 40868 24052
rect 40862 24012 40868 24024
rect 40920 24012 40926 24064
rect 42426 24052 42432 24064
rect 42387 24024 42432 24052
rect 42426 24012 42432 24024
rect 42484 24012 42490 24064
rect 42886 24012 42892 24064
rect 42944 24052 42950 24064
rect 44818 24052 44824 24064
rect 42944 24024 44824 24052
rect 42944 24012 42950 24024
rect 44818 24012 44824 24024
rect 44876 24052 44882 24064
rect 47026 24052 47032 24064
rect 44876 24024 47032 24052
rect 44876 24012 44882 24024
rect 47026 24012 47032 24024
rect 47084 24012 47090 24064
rect 1104 23962 48852 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 48852 23962
rect 1104 23888 48852 23910
rect 14090 23848 14096 23860
rect 14051 23820 14096 23848
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 15933 23851 15991 23857
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16298 23848 16304 23860
rect 15979 23820 16304 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 17862 23848 17868 23860
rect 17823 23820 17868 23848
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 19245 23851 19303 23857
rect 19245 23817 19257 23851
rect 19291 23848 19303 23851
rect 19334 23848 19340 23860
rect 19291 23820 19340 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20625 23851 20683 23857
rect 20625 23848 20637 23851
rect 20312 23820 20637 23848
rect 20312 23808 20318 23820
rect 20625 23817 20637 23820
rect 20671 23817 20683 23851
rect 21450 23848 21456 23860
rect 21411 23820 21456 23848
rect 20625 23811 20683 23817
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 22097 23851 22155 23857
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 22186 23848 22192 23860
rect 22143 23820 22192 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 22327 23851 22385 23857
rect 22327 23817 22339 23851
rect 22373 23848 22385 23851
rect 22646 23848 22652 23860
rect 22373 23820 22652 23848
rect 22373 23817 22385 23820
rect 22327 23811 22385 23817
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 22741 23851 22799 23857
rect 22741 23817 22753 23851
rect 22787 23848 22799 23851
rect 22830 23848 22836 23860
rect 22787 23820 22836 23848
rect 22787 23817 22799 23820
rect 22741 23811 22799 23817
rect 17034 23780 17040 23792
rect 16947 23752 17040 23780
rect 17034 23740 17040 23752
rect 17092 23780 17098 23792
rect 18693 23783 18751 23789
rect 18693 23780 18705 23783
rect 17092 23752 18705 23780
rect 17092 23740 17098 23752
rect 18693 23749 18705 23752
rect 18739 23780 18751 23783
rect 19978 23780 19984 23792
rect 18739 23752 19984 23780
rect 18739 23749 18751 23752
rect 18693 23743 18751 23749
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 14645 23715 14703 23721
rect 14645 23712 14657 23715
rect 14516 23684 14657 23712
rect 14516 23672 14522 23684
rect 14645 23681 14657 23684
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23712 16543 23715
rect 16666 23712 16672 23724
rect 16531 23684 16672 23712
rect 16531 23681 16543 23684
rect 16485 23675 16543 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 18138 23712 18144 23724
rect 18099 23684 18144 23712
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 19058 23672 19064 23724
rect 19116 23712 19122 23724
rect 19702 23712 19708 23724
rect 19116 23684 19708 23712
rect 19116 23672 19122 23684
rect 19702 23672 19708 23684
rect 19760 23672 19766 23724
rect 19794 23672 19800 23724
rect 19852 23712 19858 23724
rect 21637 23715 21695 23721
rect 21637 23712 21649 23715
rect 19852 23684 21649 23712
rect 19852 23672 19858 23684
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23644 15623 23647
rect 15838 23644 15844 23656
rect 15611 23616 15844 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 15838 23604 15844 23616
rect 15896 23644 15902 23656
rect 21259 23653 21287 23684
rect 21637 23681 21649 23684
rect 21683 23681 21695 23715
rect 21637 23675 21695 23681
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 15896 23616 16221 23644
rect 15896 23604 15902 23616
rect 16209 23613 16221 23616
rect 16255 23613 16267 23647
rect 21244 23647 21302 23653
rect 21244 23644 21256 23647
rect 21222 23616 21256 23644
rect 16209 23607 16267 23613
rect 21244 23613 21256 23616
rect 21290 23613 21302 23647
rect 21244 23607 21302 23613
rect 14553 23579 14611 23585
rect 14553 23545 14565 23579
rect 14599 23576 14611 23579
rect 14966 23579 15024 23585
rect 14966 23576 14978 23579
rect 14599 23548 14978 23576
rect 14599 23545 14611 23548
rect 14553 23539 14611 23545
rect 14966 23545 14978 23548
rect 15012 23576 15024 23579
rect 15470 23576 15476 23588
rect 15012 23548 15476 23576
rect 15012 23545 15024 23548
rect 14966 23539 15024 23545
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 16224 23576 16252 23607
rect 16577 23579 16635 23585
rect 16577 23576 16589 23579
rect 16224 23548 16589 23576
rect 16577 23545 16589 23548
rect 16623 23545 16635 23579
rect 17494 23576 17500 23588
rect 17407 23548 17500 23576
rect 16577 23539 16635 23545
rect 17494 23536 17500 23548
rect 17552 23576 17558 23588
rect 18230 23576 18236 23588
rect 17552 23548 18236 23576
rect 17552 23536 17558 23548
rect 18230 23536 18236 23548
rect 18288 23536 18294 23588
rect 19702 23576 19708 23588
rect 18385 23548 19708 23576
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 18385 23508 18413 23548
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 19797 23579 19855 23585
rect 19797 23545 19809 23579
rect 19843 23576 19855 23579
rect 20162 23576 20168 23588
rect 19843 23548 20168 23576
rect 19843 23545 19855 23548
rect 19797 23539 19855 23545
rect 20162 23536 20168 23548
rect 20220 23536 20226 23588
rect 20349 23579 20407 23585
rect 20349 23545 20361 23579
rect 20395 23545 20407 23579
rect 21259 23576 21287 23607
rect 21358 23604 21364 23656
rect 21416 23644 21422 23656
rect 22256 23647 22314 23653
rect 22256 23644 22268 23647
rect 21416 23616 22268 23644
rect 21416 23604 21422 23616
rect 22256 23613 22268 23616
rect 22302 23644 22314 23647
rect 22756 23644 22784 23811
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 23382 23808 23388 23860
rect 23440 23848 23446 23860
rect 23799 23851 23857 23857
rect 23799 23848 23811 23851
rect 23440 23820 23811 23848
rect 23440 23808 23446 23820
rect 23799 23817 23811 23820
rect 23845 23817 23857 23851
rect 23799 23811 23857 23817
rect 24857 23851 24915 23857
rect 24857 23817 24869 23851
rect 24903 23848 24915 23851
rect 25406 23848 25412 23860
rect 24903 23820 25412 23848
rect 24903 23817 24915 23820
rect 24857 23811 24915 23817
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 25866 23848 25872 23860
rect 25827 23820 25872 23848
rect 25866 23808 25872 23820
rect 25924 23808 25930 23860
rect 26326 23808 26332 23860
rect 26384 23848 26390 23860
rect 26421 23851 26479 23857
rect 26421 23848 26433 23851
rect 26384 23820 26433 23848
rect 26384 23808 26390 23820
rect 26421 23817 26433 23820
rect 26467 23817 26479 23851
rect 26421 23811 26479 23817
rect 26694 23808 26700 23860
rect 26752 23848 26758 23860
rect 26789 23851 26847 23857
rect 26789 23848 26801 23851
rect 26752 23820 26801 23848
rect 26752 23808 26758 23820
rect 26789 23817 26801 23820
rect 26835 23817 26847 23851
rect 26789 23811 26847 23817
rect 26878 23808 26884 23860
rect 26936 23848 26942 23860
rect 28534 23848 28540 23860
rect 26936 23820 28540 23848
rect 26936 23808 26942 23820
rect 28534 23808 28540 23820
rect 28592 23848 28598 23860
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 28592 23820 28641 23848
rect 28592 23808 28598 23820
rect 28629 23817 28641 23820
rect 28675 23817 28687 23851
rect 29086 23848 29092 23860
rect 29047 23820 29092 23848
rect 28629 23811 28687 23817
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 30098 23808 30104 23860
rect 30156 23848 30162 23860
rect 30975 23851 31033 23857
rect 30975 23848 30987 23851
rect 30156 23820 30987 23848
rect 30156 23808 30162 23820
rect 30975 23817 30987 23820
rect 31021 23817 31033 23851
rect 31294 23848 31300 23860
rect 31255 23820 31300 23848
rect 30975 23811 31033 23817
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 32214 23808 32220 23860
rect 32272 23848 32278 23860
rect 32493 23851 32551 23857
rect 32493 23848 32505 23851
rect 32272 23820 32505 23848
rect 32272 23808 32278 23820
rect 32493 23817 32505 23820
rect 32539 23817 32551 23851
rect 32493 23811 32551 23817
rect 32907 23851 32965 23857
rect 32907 23817 32919 23851
rect 32953 23848 32965 23851
rect 36630 23848 36636 23860
rect 32953 23820 36636 23848
rect 32953 23817 32965 23820
rect 32907 23811 32965 23817
rect 36630 23808 36636 23820
rect 36688 23808 36694 23860
rect 36725 23851 36783 23857
rect 36725 23817 36737 23851
rect 36771 23848 36783 23851
rect 36906 23848 36912 23860
rect 36771 23820 36912 23848
rect 36771 23817 36783 23820
rect 36725 23811 36783 23817
rect 36906 23808 36912 23820
rect 36964 23808 36970 23860
rect 37918 23848 37924 23860
rect 37879 23820 37924 23848
rect 37918 23808 37924 23820
rect 37976 23808 37982 23860
rect 38378 23848 38384 23860
rect 38339 23820 38384 23848
rect 38378 23808 38384 23820
rect 38436 23808 38442 23860
rect 41230 23808 41236 23860
rect 41288 23848 41294 23860
rect 42245 23851 42303 23857
rect 42245 23848 42257 23851
rect 41288 23820 42257 23848
rect 41288 23808 41294 23820
rect 42245 23817 42257 23820
rect 42291 23817 42303 23851
rect 42245 23811 42303 23817
rect 43073 23851 43131 23857
rect 43073 23817 43085 23851
rect 43119 23848 43131 23851
rect 43254 23848 43260 23860
rect 43119 23820 43260 23848
rect 43119 23817 43131 23820
rect 43073 23811 43131 23817
rect 43254 23808 43260 23820
rect 43312 23808 43318 23860
rect 44542 23808 44548 23860
rect 44600 23848 44606 23860
rect 44867 23851 44925 23857
rect 44867 23848 44879 23851
rect 44600 23820 44879 23848
rect 44600 23808 44606 23820
rect 44867 23817 44879 23820
rect 44913 23817 44925 23851
rect 45830 23848 45836 23860
rect 45791 23820 45836 23848
rect 44867 23811 44925 23817
rect 45830 23808 45836 23820
rect 45888 23808 45894 23860
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 22980 23752 24900 23780
rect 22980 23740 22986 23752
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23474 23712 23480 23724
rect 23431 23684 23480 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 22302 23616 22784 23644
rect 23728 23647 23786 23653
rect 22302 23613 22314 23616
rect 22256 23607 22314 23613
rect 23728 23613 23740 23647
rect 23774 23644 23786 23647
rect 24872 23644 24900 23752
rect 24946 23740 24952 23792
rect 25004 23780 25010 23792
rect 25087 23783 25145 23789
rect 25087 23780 25099 23783
rect 25004 23752 25099 23780
rect 25004 23740 25010 23752
rect 25087 23749 25099 23752
rect 25133 23749 25145 23783
rect 25087 23743 25145 23749
rect 25501 23783 25559 23789
rect 25501 23749 25513 23783
rect 25547 23780 25559 23783
rect 31757 23783 31815 23789
rect 25547 23752 30947 23780
rect 25547 23749 25559 23752
rect 25501 23743 25559 23749
rect 25016 23647 25074 23653
rect 25016 23644 25028 23647
rect 23774 23616 24164 23644
rect 24872 23616 25028 23644
rect 23774 23613 23786 23616
rect 23728 23607 23786 23613
rect 24136 23588 24164 23616
rect 25016 23613 25028 23616
rect 25062 23644 25074 23647
rect 25516 23644 25544 23743
rect 28166 23712 28172 23724
rect 28127 23684 28172 23712
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 29822 23712 29828 23724
rect 29783 23684 29828 23712
rect 29822 23672 29828 23684
rect 29880 23672 29886 23724
rect 30190 23672 30196 23724
rect 30248 23712 30254 23724
rect 30285 23715 30343 23721
rect 30285 23712 30297 23715
rect 30248 23684 30297 23712
rect 30248 23672 30254 23684
rect 30285 23681 30297 23684
rect 30331 23681 30343 23715
rect 30285 23675 30343 23681
rect 25062 23616 25544 23644
rect 26028 23647 26086 23653
rect 25062 23613 25074 23616
rect 25016 23607 25074 23613
rect 26028 23613 26040 23647
rect 26074 23644 26086 23647
rect 26326 23644 26332 23656
rect 26074 23616 26332 23644
rect 26074 23613 26086 23616
rect 26028 23607 26086 23613
rect 26326 23604 26332 23616
rect 26384 23604 26390 23656
rect 27338 23604 27344 23656
rect 27396 23644 27402 23656
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 27396 23616 27445 23644
rect 27396 23604 27402 23616
rect 27433 23613 27445 23616
rect 27479 23644 27491 23647
rect 27617 23647 27675 23653
rect 27617 23644 27629 23647
rect 27479 23616 27629 23644
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 27617 23613 27629 23616
rect 27663 23613 27675 23647
rect 27617 23607 27675 23613
rect 28077 23647 28135 23653
rect 28077 23613 28089 23647
rect 28123 23644 28135 23647
rect 28258 23644 28264 23656
rect 28123 23616 28264 23644
rect 28123 23613 28135 23616
rect 28077 23607 28135 23613
rect 28258 23604 28264 23616
rect 28316 23604 28322 23656
rect 30919 23653 30947 23752
rect 31757 23749 31769 23783
rect 31803 23780 31815 23783
rect 34238 23780 34244 23792
rect 31803 23752 34244 23780
rect 31803 23749 31815 23752
rect 31757 23743 31815 23749
rect 30904 23647 30962 23653
rect 30904 23613 30916 23647
rect 30950 23644 30962 23647
rect 31772 23644 31800 23743
rect 34238 23740 34244 23752
rect 34296 23740 34302 23792
rect 35894 23780 35900 23792
rect 34992 23752 35900 23780
rect 32217 23715 32275 23721
rect 32217 23681 32229 23715
rect 32263 23712 32275 23715
rect 32306 23712 32312 23724
rect 32263 23684 32312 23712
rect 32263 23681 32275 23684
rect 32217 23675 32275 23681
rect 32306 23672 32312 23684
rect 32364 23672 32370 23724
rect 34992 23721 35020 23752
rect 35894 23740 35900 23752
rect 35952 23740 35958 23792
rect 35986 23740 35992 23792
rect 36044 23780 36050 23792
rect 36081 23783 36139 23789
rect 36081 23780 36093 23783
rect 36044 23752 36093 23780
rect 36044 23740 36050 23752
rect 36081 23749 36093 23752
rect 36127 23749 36139 23783
rect 40034 23780 40040 23792
rect 36081 23743 36139 23749
rect 36407 23752 40040 23780
rect 33919 23715 33977 23721
rect 33919 23681 33931 23715
rect 33965 23712 33977 23715
rect 34977 23715 35035 23721
rect 34977 23712 34989 23715
rect 33965 23684 34989 23712
rect 33965 23681 33977 23684
rect 33919 23675 33977 23681
rect 34977 23681 34989 23684
rect 35023 23681 35035 23715
rect 35342 23712 35348 23724
rect 35303 23684 35348 23712
rect 34977 23675 35035 23681
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 30950 23616 31800 23644
rect 30950 23613 30962 23616
rect 30904 23607 30962 23613
rect 31846 23604 31852 23656
rect 31904 23644 31910 23656
rect 32836 23647 32894 23653
rect 32836 23644 32848 23647
rect 31904 23616 32848 23644
rect 31904 23604 31910 23616
rect 32836 23613 32848 23616
rect 32882 23644 32894 23647
rect 33229 23647 33287 23653
rect 33229 23644 33241 23647
rect 32882 23616 33241 23644
rect 32882 23613 32894 23616
rect 32836 23607 32894 23613
rect 33229 23613 33241 23616
rect 33275 23644 33287 23647
rect 33318 23644 33324 23656
rect 33275 23616 33324 23644
rect 33275 23613 33287 23616
rect 33229 23607 33287 23613
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 33816 23647 33874 23653
rect 33816 23613 33828 23647
rect 33862 23613 33874 23647
rect 33816 23607 33874 23613
rect 23842 23576 23848 23588
rect 21259 23548 23848 23576
rect 20349 23539 20407 23545
rect 15252 23480 18413 23508
rect 15252 23468 15258 23480
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 20364 23508 20392 23539
rect 23842 23536 23848 23548
rect 23900 23536 23906 23588
rect 24118 23536 24124 23588
rect 24176 23576 24182 23588
rect 24213 23579 24271 23585
rect 24213 23576 24225 23579
rect 24176 23548 24225 23576
rect 24176 23536 24182 23548
rect 24213 23545 24225 23548
rect 24259 23576 24271 23579
rect 27706 23576 27712 23588
rect 24259 23548 27712 23576
rect 24259 23545 24271 23548
rect 24213 23539 24271 23545
rect 27706 23536 27712 23548
rect 27764 23536 27770 23588
rect 29362 23576 29368 23588
rect 29323 23548 29368 23576
rect 29362 23536 29368 23548
rect 29420 23536 29426 23588
rect 29457 23579 29515 23585
rect 29457 23545 29469 23579
rect 29503 23545 29515 23579
rect 29457 23539 29515 23545
rect 19484 23480 20392 23508
rect 26099 23511 26157 23517
rect 19484 23468 19490 23480
rect 26099 23477 26111 23511
rect 26145 23508 26157 23511
rect 26326 23508 26332 23520
rect 26145 23480 26332 23508
rect 26145 23477 26157 23480
rect 26099 23471 26157 23477
rect 26326 23468 26332 23480
rect 26384 23468 26390 23520
rect 29086 23468 29092 23520
rect 29144 23508 29150 23520
rect 29472 23508 29500 23539
rect 33594 23536 33600 23588
rect 33652 23576 33658 23588
rect 33689 23579 33747 23585
rect 33689 23576 33701 23579
rect 33652 23548 33701 23576
rect 33652 23536 33658 23548
rect 33689 23545 33701 23548
rect 33735 23576 33747 23579
rect 33831 23576 33859 23607
rect 35069 23579 35127 23585
rect 33735 23548 34652 23576
rect 33735 23545 33747 23548
rect 33689 23539 33747 23545
rect 29638 23508 29644 23520
rect 29144 23480 29644 23508
rect 29144 23468 29150 23480
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 34425 23511 34483 23517
rect 34425 23477 34437 23511
rect 34471 23508 34483 23511
rect 34514 23508 34520 23520
rect 34471 23480 34520 23508
rect 34471 23477 34483 23480
rect 34425 23471 34483 23477
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 34624 23508 34652 23548
rect 35069 23545 35081 23579
rect 35115 23576 35127 23579
rect 35250 23576 35256 23588
rect 35115 23548 35256 23576
rect 35115 23545 35127 23548
rect 35069 23539 35127 23545
rect 35250 23536 35256 23548
rect 35308 23536 35314 23588
rect 36407 23508 36435 23752
rect 40034 23740 40040 23752
rect 40092 23740 40098 23792
rect 40862 23740 40868 23792
rect 40920 23780 40926 23792
rect 41601 23783 41659 23789
rect 41601 23780 41613 23783
rect 40920 23752 41613 23780
rect 40920 23740 40926 23752
rect 41601 23749 41613 23752
rect 41647 23749 41659 23783
rect 41601 23743 41659 23749
rect 46106 23740 46112 23792
rect 46164 23780 46170 23792
rect 46247 23783 46305 23789
rect 46247 23780 46259 23783
rect 46164 23752 46259 23780
rect 46164 23740 46170 23752
rect 46247 23749 46259 23752
rect 46293 23749 46305 23783
rect 46247 23743 46305 23749
rect 37274 23672 37280 23724
rect 37332 23712 37338 23724
rect 37553 23715 37611 23721
rect 37553 23712 37565 23715
rect 37332 23684 37565 23712
rect 37332 23672 37338 23684
rect 37553 23681 37565 23684
rect 37599 23712 37611 23715
rect 38470 23712 38476 23724
rect 37599 23684 38476 23712
rect 37599 23681 37611 23684
rect 37553 23675 37611 23681
rect 38470 23672 38476 23684
rect 38528 23672 38534 23724
rect 39942 23672 39948 23724
rect 40000 23712 40006 23724
rect 40678 23712 40684 23724
rect 40000 23684 40684 23712
rect 40000 23672 40006 23684
rect 40678 23672 40684 23684
rect 40736 23672 40742 23724
rect 42705 23715 42763 23721
rect 42705 23681 42717 23715
rect 42751 23712 42763 23715
rect 43257 23715 43315 23721
rect 43257 23712 43269 23715
rect 42751 23684 43269 23712
rect 42751 23681 42763 23684
rect 42705 23675 42763 23681
rect 43257 23681 43269 23684
rect 43303 23712 43315 23715
rect 43346 23712 43352 23724
rect 43303 23684 43352 23712
rect 43303 23681 43315 23684
rect 43257 23675 43315 23681
rect 43346 23672 43352 23684
rect 43404 23672 43410 23724
rect 43622 23712 43628 23724
rect 43583 23684 43628 23712
rect 43622 23672 43628 23684
rect 43680 23672 43686 23724
rect 45370 23672 45376 23724
rect 45428 23712 45434 23724
rect 45830 23712 45836 23724
rect 45428 23684 45836 23712
rect 45428 23672 45434 23684
rect 45830 23672 45836 23684
rect 45888 23672 45894 23724
rect 38654 23604 38660 23656
rect 38712 23644 38718 23656
rect 38841 23647 38899 23653
rect 38841 23644 38853 23647
rect 38712 23616 38853 23644
rect 38712 23604 38718 23616
rect 38841 23613 38853 23616
rect 38887 23613 38899 23647
rect 39390 23644 39396 23656
rect 39351 23616 39396 23644
rect 38841 23607 38899 23613
rect 39390 23604 39396 23616
rect 39448 23604 39454 23656
rect 39577 23647 39635 23653
rect 39577 23613 39589 23647
rect 39623 23644 39635 23647
rect 42426 23644 42432 23656
rect 39623 23616 42432 23644
rect 39623 23613 39635 23616
rect 39577 23607 39635 23613
rect 42426 23604 42432 23616
rect 42484 23604 42490 23656
rect 44796 23647 44854 23653
rect 44796 23613 44808 23647
rect 44842 23644 44854 23647
rect 45094 23644 45100 23656
rect 44842 23616 45100 23644
rect 44842 23613 44854 23616
rect 44796 23607 44854 23613
rect 45094 23604 45100 23616
rect 45152 23644 45158 23656
rect 45189 23647 45247 23653
rect 45189 23644 45201 23647
rect 45152 23616 45201 23644
rect 45152 23604 45158 23616
rect 45189 23613 45201 23616
rect 45235 23613 45247 23647
rect 45189 23607 45247 23613
rect 45646 23604 45652 23656
rect 45704 23644 45710 23656
rect 46144 23647 46202 23653
rect 46144 23644 46156 23647
rect 45704 23616 46156 23644
rect 45704 23604 45710 23616
rect 46144 23613 46156 23616
rect 46190 23644 46202 23647
rect 46569 23647 46627 23653
rect 46569 23644 46581 23647
rect 46190 23616 46581 23644
rect 46190 23613 46202 23616
rect 46144 23607 46202 23613
rect 46569 23613 46581 23616
rect 46615 23613 46627 23647
rect 46569 23607 46627 23613
rect 36906 23576 36912 23588
rect 36867 23548 36912 23576
rect 36906 23536 36912 23548
rect 36964 23536 36970 23588
rect 36998 23536 37004 23588
rect 37056 23576 37062 23588
rect 41002 23579 41060 23585
rect 37056 23548 37101 23576
rect 37056 23536 37062 23548
rect 41002 23545 41014 23579
rect 41048 23576 41060 23579
rect 41877 23579 41935 23585
rect 41877 23576 41889 23579
rect 41048 23548 41889 23576
rect 41048 23545 41060 23548
rect 41002 23539 41060 23545
rect 41877 23545 41889 23548
rect 41923 23545 41935 23579
rect 41877 23539 41935 23545
rect 38654 23508 38660 23520
rect 34624 23480 36435 23508
rect 38615 23480 38660 23508
rect 38654 23468 38660 23480
rect 38712 23468 38718 23520
rect 39945 23511 40003 23517
rect 39945 23477 39957 23511
rect 39991 23508 40003 23511
rect 40310 23508 40316 23520
rect 39991 23480 40316 23508
rect 39991 23477 40003 23480
rect 39945 23471 40003 23477
rect 40310 23468 40316 23480
rect 40368 23508 40374 23520
rect 41017 23508 41045 23539
rect 40368 23480 41045 23508
rect 41892 23508 41920 23539
rect 43346 23536 43352 23588
rect 43404 23576 43410 23588
rect 43404 23548 43449 23576
rect 43404 23536 43410 23548
rect 44269 23511 44327 23517
rect 44269 23508 44281 23511
rect 41892 23480 44281 23508
rect 40368 23468 40374 23480
rect 44269 23477 44281 23480
rect 44315 23508 44327 23511
rect 44358 23508 44364 23520
rect 44315 23480 44364 23508
rect 44315 23477 44327 23480
rect 44269 23471 44327 23477
rect 44358 23468 44364 23480
rect 44416 23468 44422 23520
rect 1104 23418 48852 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 48852 23418
rect 1104 23344 48852 23366
rect 14458 23264 14464 23316
rect 14516 23304 14522 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14516 23276 14657 23304
rect 14516 23264 14522 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 19242 23304 19248 23316
rect 14645 23267 14703 23273
rect 16408 23276 18828 23304
rect 19203 23276 19248 23304
rect 15838 23236 15844 23248
rect 15799 23208 15844 23236
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 16114 23196 16120 23248
rect 16172 23236 16178 23248
rect 16408 23245 16436 23276
rect 16393 23239 16451 23245
rect 16393 23236 16405 23239
rect 16172 23208 16405 23236
rect 16172 23196 16178 23208
rect 16393 23205 16405 23208
rect 16439 23205 16451 23239
rect 16393 23199 16451 23205
rect 18233 23239 18291 23245
rect 18233 23205 18245 23239
rect 18279 23236 18291 23239
rect 18322 23236 18328 23248
rect 18279 23208 18328 23236
rect 18279 23205 18291 23208
rect 18233 23199 18291 23205
rect 18322 23196 18328 23208
rect 18380 23196 18386 23248
rect 18800 23245 18828 23276
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 21818 23304 21824 23316
rect 21779 23276 21824 23304
rect 21818 23264 21824 23276
rect 21876 23264 21882 23316
rect 23382 23304 23388 23316
rect 23343 23276 23388 23304
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 24946 23304 24952 23316
rect 24907 23276 24952 23304
rect 24946 23264 24952 23276
rect 25004 23264 25010 23316
rect 28166 23304 28172 23316
rect 28127 23276 28172 23304
rect 28166 23264 28172 23276
rect 28224 23264 28230 23316
rect 33229 23307 33287 23313
rect 33229 23304 33241 23307
rect 32876 23276 33241 23304
rect 18785 23239 18843 23245
rect 18785 23205 18797 23239
rect 18831 23236 18843 23239
rect 20622 23236 20628 23248
rect 18831 23208 20628 23236
rect 18831 23205 18843 23208
rect 18785 23199 18843 23205
rect 20622 23196 20628 23208
rect 20680 23196 20686 23248
rect 22557 23239 22615 23245
rect 22557 23205 22569 23239
rect 22603 23236 22615 23239
rect 23290 23236 23296 23248
rect 22603 23208 23296 23236
rect 22603 23205 22615 23208
rect 22557 23199 22615 23205
rect 23290 23196 23296 23208
rect 23348 23196 23354 23248
rect 26418 23196 26424 23248
rect 26476 23236 26482 23248
rect 26602 23236 26608 23248
rect 26476 23208 26608 23236
rect 26476 23196 26482 23208
rect 26602 23196 26608 23208
rect 26660 23236 26666 23248
rect 26697 23239 26755 23245
rect 26697 23236 26709 23239
rect 26660 23208 26709 23236
rect 26660 23196 26666 23208
rect 26697 23205 26709 23208
rect 26743 23205 26755 23239
rect 27246 23236 27252 23248
rect 27207 23208 27252 23236
rect 26697 23199 26755 23205
rect 27246 23196 27252 23208
rect 27304 23196 27310 23248
rect 27522 23196 27528 23248
rect 27580 23236 27586 23248
rect 29546 23236 29552 23248
rect 27580 23208 29552 23236
rect 27580 23196 27586 23208
rect 29546 23196 29552 23208
rect 29604 23196 29610 23248
rect 29638 23196 29644 23248
rect 29696 23236 29702 23248
rect 29696 23208 29741 23236
rect 29696 23196 29702 23208
rect 31846 23196 31852 23248
rect 31904 23236 31910 23248
rect 32309 23239 32367 23245
rect 32309 23236 32321 23239
rect 31904 23208 32321 23236
rect 31904 23196 31910 23208
rect 32309 23205 32321 23208
rect 32355 23205 32367 23239
rect 32309 23199 32367 23205
rect 32490 23196 32496 23248
rect 32548 23236 32554 23248
rect 32876 23245 32904 23276
rect 33229 23273 33241 23276
rect 33275 23304 33287 23307
rect 33502 23304 33508 23316
rect 33275 23276 33508 23304
rect 33275 23273 33287 23276
rect 33229 23267 33287 23273
rect 33502 23264 33508 23276
rect 33560 23264 33566 23316
rect 34054 23304 34060 23316
rect 34015 23276 34060 23304
rect 34054 23264 34060 23276
rect 34112 23264 34118 23316
rect 34977 23307 35035 23313
rect 34977 23273 34989 23307
rect 35023 23304 35035 23307
rect 35250 23304 35256 23316
rect 35023 23276 35256 23304
rect 35023 23273 35035 23276
rect 34977 23267 35035 23273
rect 35250 23264 35256 23276
rect 35308 23264 35314 23316
rect 36170 23304 36176 23316
rect 36131 23276 36176 23304
rect 36170 23264 36176 23276
rect 36228 23264 36234 23316
rect 36679 23307 36737 23313
rect 36679 23273 36691 23307
rect 36725 23304 36737 23307
rect 36906 23304 36912 23316
rect 36725 23276 36912 23304
rect 36725 23273 36737 23276
rect 36679 23267 36737 23273
rect 36906 23264 36912 23276
rect 36964 23304 36970 23316
rect 37001 23307 37059 23313
rect 37001 23304 37013 23307
rect 36964 23276 37013 23304
rect 36964 23264 36970 23276
rect 37001 23273 37013 23276
rect 37047 23273 37059 23307
rect 37001 23267 37059 23273
rect 37090 23264 37096 23316
rect 37148 23304 37154 23316
rect 37148 23276 39344 23304
rect 37148 23264 37154 23276
rect 32861 23239 32919 23245
rect 32861 23236 32873 23239
rect 32548 23208 32873 23236
rect 32548 23196 32554 23208
rect 32861 23205 32873 23208
rect 32907 23205 32919 23239
rect 38838 23236 38844 23248
rect 32861 23199 32919 23205
rect 34072 23208 38844 23236
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23168 14151 23171
rect 14274 23168 14280 23180
rect 14139 23140 14280 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 19610 23168 19616 23180
rect 19571 23140 19616 23168
rect 19610 23128 19616 23140
rect 19668 23128 19674 23180
rect 21358 23168 21364 23180
rect 21319 23140 21364 23168
rect 21358 23128 21364 23140
rect 21416 23128 21422 23180
rect 23201 23171 23259 23177
rect 23201 23137 23213 23171
rect 23247 23168 23259 23171
rect 24004 23171 24062 23177
rect 24004 23168 24016 23171
rect 23247 23140 24016 23168
rect 23247 23137 23259 23140
rect 23201 23131 23259 23137
rect 24004 23137 24016 23140
rect 24050 23168 24062 23171
rect 24854 23168 24860 23180
rect 24050 23140 24860 23168
rect 24050 23137 24062 23140
rect 24004 23131 24062 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 25038 23128 25044 23180
rect 25096 23168 25102 23180
rect 25168 23171 25226 23177
rect 25168 23168 25180 23171
rect 25096 23140 25180 23168
rect 25096 23128 25102 23140
rect 25168 23137 25180 23140
rect 25214 23168 25226 23171
rect 26050 23168 26056 23180
rect 25214 23140 26056 23168
rect 25214 23137 25226 23140
rect 25168 23131 25226 23137
rect 26050 23128 26056 23140
rect 26108 23128 26114 23180
rect 33870 23128 33876 23180
rect 33928 23168 33934 23180
rect 34072 23177 34100 23208
rect 38838 23196 38844 23208
rect 38896 23196 38902 23248
rect 39316 23180 39344 23276
rect 39482 23264 39488 23316
rect 39540 23304 39546 23316
rect 40313 23307 40371 23313
rect 40313 23304 40325 23307
rect 39540 23276 40325 23304
rect 39540 23264 39546 23276
rect 40313 23273 40325 23276
rect 40359 23273 40371 23307
rect 40678 23304 40684 23316
rect 40639 23276 40684 23304
rect 40313 23267 40371 23273
rect 40678 23264 40684 23276
rect 40736 23264 40742 23316
rect 44266 23304 44272 23316
rect 42766 23276 44272 23304
rect 40037 23239 40095 23245
rect 40037 23205 40049 23239
rect 40083 23236 40095 23239
rect 41230 23236 41236 23248
rect 40083 23208 41236 23236
rect 40083 23205 40095 23208
rect 40037 23199 40095 23205
rect 41230 23196 41236 23208
rect 41288 23196 41294 23248
rect 41601 23239 41659 23245
rect 41601 23205 41613 23239
rect 41647 23236 41659 23239
rect 42766 23236 42794 23276
rect 44266 23264 44272 23276
rect 44324 23264 44330 23316
rect 44683 23307 44741 23313
rect 44683 23273 44695 23307
rect 44729 23304 44741 23307
rect 45462 23304 45468 23316
rect 44729 23276 45468 23304
rect 44729 23273 44741 23276
rect 44683 23267 44741 23273
rect 45462 23264 45468 23276
rect 45520 23264 45526 23316
rect 46106 23304 46112 23316
rect 46067 23276 46112 23304
rect 46106 23264 46112 23276
rect 46164 23264 46170 23316
rect 41647 23208 42794 23236
rect 41647 23205 41659 23208
rect 41601 23199 41659 23205
rect 34057 23171 34115 23177
rect 34057 23168 34069 23171
rect 33928 23140 34069 23168
rect 33928 23128 33934 23140
rect 34057 23137 34069 23140
rect 34103 23137 34115 23171
rect 34057 23131 34115 23137
rect 34146 23128 34152 23180
rect 34204 23168 34210 23180
rect 34241 23171 34299 23177
rect 34241 23168 34253 23171
rect 34204 23140 34253 23168
rect 34204 23128 34210 23140
rect 34241 23137 34253 23140
rect 34287 23137 34299 23171
rect 34241 23131 34299 23137
rect 35412 23171 35470 23177
rect 35412 23137 35424 23171
rect 35458 23168 35470 23171
rect 35986 23168 35992 23180
rect 35458 23140 35992 23168
rect 35458 23137 35470 23140
rect 35412 23131 35470 23137
rect 35986 23128 35992 23140
rect 36044 23128 36050 23180
rect 36541 23171 36599 23177
rect 36541 23137 36553 23171
rect 36587 23168 36599 23171
rect 36630 23168 36636 23180
rect 36587 23140 36636 23168
rect 36587 23137 36599 23140
rect 36541 23131 36599 23137
rect 36630 23128 36636 23140
rect 36688 23128 36694 23180
rect 37645 23171 37703 23177
rect 37645 23137 37657 23171
rect 37691 23168 37703 23171
rect 37734 23168 37740 23180
rect 37691 23140 37740 23168
rect 37691 23137 37703 23140
rect 37645 23131 37703 23137
rect 37734 23128 37740 23140
rect 37792 23128 37798 23180
rect 39298 23168 39304 23180
rect 39259 23140 39304 23168
rect 39298 23128 39304 23140
rect 39356 23128 39362 23180
rect 39390 23128 39396 23180
rect 39448 23168 39454 23180
rect 39853 23171 39911 23177
rect 39853 23168 39865 23171
rect 39448 23140 39865 23168
rect 39448 23128 39454 23140
rect 39853 23137 39865 23140
rect 39899 23137 39911 23171
rect 40862 23168 40868 23180
rect 40823 23140 40868 23168
rect 39853 23131 39911 23137
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23100 15807 23103
rect 16114 23100 16120 23112
rect 15795 23072 16120 23100
rect 15795 23069 15807 23072
rect 15749 23063 15807 23069
rect 16114 23060 16120 23072
rect 16172 23060 16178 23112
rect 18138 23100 18144 23112
rect 18099 23072 18144 23100
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 19751 23103 19809 23109
rect 19751 23100 19763 23103
rect 18288 23072 19763 23100
rect 18288 23060 18294 23072
rect 19751 23069 19763 23072
rect 19797 23069 19809 23103
rect 22462 23100 22468 23112
rect 22423 23072 22468 23100
rect 19751 23063 19809 23069
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 22738 23100 22744 23112
rect 22699 23072 22744 23100
rect 22738 23060 22744 23072
rect 22796 23100 22802 23112
rect 24394 23100 24400 23112
rect 22796 23072 24400 23100
rect 22796 23060 22802 23072
rect 24394 23060 24400 23072
rect 24452 23060 24458 23112
rect 24486 23060 24492 23112
rect 24544 23100 24550 23112
rect 26605 23103 26663 23109
rect 26605 23100 26617 23103
rect 24544 23072 26617 23100
rect 24544 23060 24550 23072
rect 26605 23069 26617 23072
rect 26651 23100 26663 23103
rect 27338 23100 27344 23112
rect 26651 23072 27344 23100
rect 26651 23069 26663 23072
rect 26605 23063 26663 23069
rect 27338 23060 27344 23072
rect 27396 23060 27402 23112
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23100 28411 23103
rect 28534 23100 28540 23112
rect 28399 23072 28540 23100
rect 28399 23069 28411 23072
rect 28353 23063 28411 23069
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 30006 23100 30012 23112
rect 29967 23072 30012 23100
rect 30006 23060 30012 23072
rect 30064 23060 30070 23112
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 32214 23100 32220 23112
rect 31067 23072 32220 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 32214 23060 32220 23072
rect 32272 23060 32278 23112
rect 33318 23060 33324 23112
rect 33376 23100 33382 23112
rect 37918 23100 37924 23112
rect 33376 23072 37924 23100
rect 33376 23060 33382 23072
rect 37918 23060 37924 23072
rect 37976 23060 37982 23112
rect 38930 23100 38936 23112
rect 38843 23072 38936 23100
rect 38930 23060 38936 23072
rect 38988 23100 38994 23112
rect 39408 23100 39436 23128
rect 38988 23072 39436 23100
rect 39868 23100 39896 23131
rect 40862 23128 40868 23140
rect 40920 23128 40926 23180
rect 40954 23128 40960 23180
rect 41012 23168 41018 23180
rect 41325 23171 41383 23177
rect 41325 23168 41337 23171
rect 41012 23140 41337 23168
rect 41012 23128 41018 23140
rect 41325 23137 41337 23140
rect 41371 23137 41383 23171
rect 41325 23131 41383 23137
rect 43416 23171 43474 23177
rect 43416 23137 43428 23171
rect 43462 23168 43474 23171
rect 43622 23168 43628 23180
rect 43462 23140 43628 23168
rect 43462 23137 43474 23140
rect 43416 23131 43474 23137
rect 43622 23128 43628 23140
rect 43680 23168 43686 23180
rect 43990 23168 43996 23180
rect 43680 23140 43996 23168
rect 43680 23128 43686 23140
rect 43990 23128 43996 23140
rect 44048 23128 44054 23180
rect 44634 23177 44640 23180
rect 44612 23171 44640 23177
rect 44612 23168 44624 23171
rect 44547 23140 44624 23168
rect 44612 23137 44624 23140
rect 44692 23168 44698 23180
rect 45002 23168 45008 23180
rect 44692 23140 45008 23168
rect 44612 23131 44640 23137
rect 44634 23128 44640 23131
rect 44692 23128 44698 23140
rect 45002 23128 45008 23140
rect 45060 23128 45066 23180
rect 40972 23100 41000 23128
rect 39868 23072 41000 23100
rect 38988 23060 38994 23072
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 23201 23035 23259 23041
rect 23201 23032 23213 23035
rect 21968 23004 23213 23032
rect 21968 22992 21974 23004
rect 23201 23001 23213 23004
rect 23247 23001 23259 23035
rect 24762 23032 24768 23044
rect 23201 22995 23259 23001
rect 23446 23004 24768 23032
rect 14323 22967 14381 22973
rect 14323 22933 14335 22967
rect 14369 22964 14381 22967
rect 15654 22964 15660 22976
rect 14369 22936 15660 22964
rect 14369 22933 14381 22936
rect 14323 22927 14381 22933
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 16666 22964 16672 22976
rect 16627 22936 16672 22964
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 20162 22964 20168 22976
rect 20123 22936 20168 22964
rect 20162 22924 20168 22936
rect 20220 22924 20226 22976
rect 21545 22967 21603 22973
rect 21545 22933 21557 22967
rect 21591 22964 21603 22967
rect 23446 22964 23474 23004
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 25406 22992 25412 23044
rect 25464 23032 25470 23044
rect 25593 23035 25651 23041
rect 25593 23032 25605 23035
rect 25464 23004 25605 23032
rect 25464 22992 25470 23004
rect 25593 23001 25605 23004
rect 25639 23001 25651 23035
rect 25593 22995 25651 23001
rect 38194 22992 38200 23044
rect 38252 23032 38258 23044
rect 40218 23032 40224 23044
rect 38252 23004 40224 23032
rect 38252 22992 38258 23004
rect 40218 22992 40224 23004
rect 40276 22992 40282 23044
rect 43162 22992 43168 23044
rect 43220 23032 43226 23044
rect 43898 23032 43904 23044
rect 43220 23004 43904 23032
rect 43220 22992 43226 23004
rect 43898 22992 43904 23004
rect 43956 22992 43962 23044
rect 23842 22964 23848 22976
rect 21591 22936 23474 22964
rect 23755 22936 23848 22964
rect 21591 22933 21603 22936
rect 21545 22927 21603 22933
rect 23842 22924 23848 22936
rect 23900 22964 23906 22976
rect 24075 22967 24133 22973
rect 24075 22964 24087 22967
rect 23900 22936 24087 22964
rect 23900 22924 23906 22936
rect 24075 22933 24087 22936
rect 24121 22933 24133 22967
rect 24075 22927 24133 22933
rect 25271 22967 25329 22973
rect 25271 22933 25283 22967
rect 25317 22964 25329 22967
rect 25498 22964 25504 22976
rect 25317 22936 25504 22964
rect 25317 22933 25329 22936
rect 25271 22927 25329 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 27706 22964 27712 22976
rect 27667 22936 27712 22964
rect 27706 22924 27712 22936
rect 27764 22964 27770 22976
rect 28258 22964 28264 22976
rect 27764 22936 28264 22964
rect 27764 22924 27770 22936
rect 28258 22924 28264 22936
rect 28316 22924 28322 22976
rect 28583 22967 28641 22973
rect 28583 22933 28595 22967
rect 28629 22964 28641 22967
rect 29178 22964 29184 22976
rect 28629 22936 29184 22964
rect 28629 22933 28641 22936
rect 28583 22927 28641 22933
rect 29178 22924 29184 22936
rect 29236 22924 29242 22976
rect 29362 22964 29368 22976
rect 29323 22936 29368 22964
rect 29362 22924 29368 22936
rect 29420 22924 29426 22976
rect 35250 22924 35256 22976
rect 35308 22964 35314 22976
rect 35483 22967 35541 22973
rect 35483 22964 35495 22967
rect 35308 22936 35495 22964
rect 35308 22924 35314 22936
rect 35483 22933 35495 22936
rect 35529 22933 35541 22967
rect 35483 22927 35541 22933
rect 37182 22924 37188 22976
rect 37240 22964 37246 22976
rect 37875 22967 37933 22973
rect 37875 22964 37887 22967
rect 37240 22936 37887 22964
rect 37240 22924 37246 22936
rect 37875 22933 37887 22936
rect 37921 22933 37933 22967
rect 37875 22927 37933 22933
rect 42610 22924 42616 22976
rect 42668 22964 42674 22976
rect 43487 22967 43545 22973
rect 43487 22964 43499 22967
rect 42668 22936 43499 22964
rect 42668 22924 42674 22936
rect 43487 22933 43499 22936
rect 43533 22933 43545 22967
rect 43487 22927 43545 22933
rect 1104 22874 48852 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 48852 22874
rect 1104 22800 48852 22822
rect 14274 22760 14280 22772
rect 14235 22732 14280 22760
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 15657 22763 15715 22769
rect 15657 22729 15669 22763
rect 15703 22760 15715 22763
rect 15838 22760 15844 22772
rect 15703 22732 15844 22760
rect 15703 22729 15715 22732
rect 15657 22723 15715 22729
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 17494 22760 17500 22772
rect 17455 22732 17500 22760
rect 17494 22720 17500 22732
rect 17552 22760 17558 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 17552 22732 17785 22760
rect 17552 22720 17558 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 17773 22723 17831 22729
rect 21913 22763 21971 22769
rect 21913 22729 21925 22763
rect 21959 22760 21971 22763
rect 22186 22760 22192 22772
rect 21959 22732 22192 22760
rect 21959 22729 21971 22732
rect 21913 22723 21971 22729
rect 22186 22720 22192 22732
rect 22244 22760 22250 22772
rect 23109 22763 23167 22769
rect 23109 22760 23121 22763
rect 22244 22732 23121 22760
rect 22244 22720 22250 22732
rect 23109 22729 23121 22732
rect 23155 22760 23167 22763
rect 23290 22760 23296 22772
rect 23155 22732 23296 22760
rect 23155 22729 23167 22732
rect 23109 22723 23167 22729
rect 23290 22720 23296 22732
rect 23348 22720 23354 22772
rect 25038 22720 25044 22772
rect 25096 22760 25102 22772
rect 25133 22763 25191 22769
rect 25133 22760 25145 22763
rect 25096 22732 25145 22760
rect 25096 22720 25102 22732
rect 25133 22729 25145 22732
rect 25179 22729 25191 22763
rect 26418 22760 26424 22772
rect 26379 22732 26424 22760
rect 25133 22723 25191 22729
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 29362 22720 29368 22772
rect 29420 22760 29426 22772
rect 30975 22763 31033 22769
rect 30975 22760 30987 22763
rect 29420 22732 30987 22760
rect 29420 22720 29426 22732
rect 30975 22729 30987 22732
rect 31021 22729 31033 22763
rect 31846 22760 31852 22772
rect 31807 22732 31852 22760
rect 30975 22723 31033 22729
rect 31846 22720 31852 22732
rect 31904 22720 31910 22772
rect 32214 22760 32220 22772
rect 32175 22732 32220 22760
rect 32214 22720 32220 22732
rect 32272 22720 32278 22772
rect 33870 22760 33876 22772
rect 33831 22732 33876 22760
rect 33870 22720 33876 22732
rect 33928 22720 33934 22772
rect 36630 22760 36636 22772
rect 34256 22732 35664 22760
rect 36543 22732 36636 22760
rect 20622 22692 20628 22704
rect 20583 22664 20628 22692
rect 20622 22652 20628 22664
rect 20680 22652 20686 22704
rect 21358 22652 21364 22704
rect 21416 22692 21422 22704
rect 21453 22695 21511 22701
rect 21453 22692 21465 22695
rect 21416 22664 21465 22692
rect 21416 22652 21422 22664
rect 21453 22661 21465 22664
rect 21499 22692 21511 22695
rect 23750 22692 23756 22704
rect 21499 22664 23756 22692
rect 21499 22661 21511 22664
rect 21453 22655 21511 22661
rect 23750 22652 23756 22664
rect 23808 22652 23814 22704
rect 24394 22652 24400 22704
rect 24452 22692 24458 22704
rect 25774 22692 25780 22704
rect 24452 22664 25780 22692
rect 24452 22652 24458 22664
rect 14875 22627 14933 22633
rect 14875 22593 14887 22627
rect 14921 22624 14933 22627
rect 16114 22624 16120 22636
rect 14921 22596 16120 22624
rect 14921 22593 14933 22596
rect 14875 22587 14933 22593
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 18417 22627 18475 22633
rect 18417 22624 18429 22627
rect 16531 22596 18429 22624
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 18417 22593 18429 22596
rect 18463 22624 18475 22627
rect 19150 22624 19156 22636
rect 18463 22596 19156 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 22370 22624 22376 22636
rect 22331 22596 22376 22624
rect 22370 22584 22376 22596
rect 22428 22624 22434 22636
rect 22922 22624 22928 22636
rect 22428 22596 22928 22624
rect 22428 22584 22434 22596
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23842 22624 23848 22636
rect 23803 22596 23848 22624
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 24854 22624 24860 22636
rect 24815 22596 24860 22624
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 25700 22633 25728 22664
rect 25774 22652 25780 22664
rect 25832 22652 25838 22704
rect 29917 22695 29975 22701
rect 29917 22661 29929 22695
rect 29963 22692 29975 22695
rect 30374 22692 30380 22704
rect 29963 22664 30380 22692
rect 29963 22661 29975 22664
rect 29917 22655 29975 22661
rect 30374 22652 30380 22664
rect 30432 22652 30438 22704
rect 25685 22627 25743 22633
rect 25685 22593 25697 22627
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26970 22624 26976 22636
rect 26384 22596 26976 22624
rect 26384 22584 26390 22596
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27154 22584 27160 22636
rect 27212 22624 27218 22636
rect 27249 22627 27307 22633
rect 27249 22624 27261 22627
rect 27212 22596 27261 22624
rect 27212 22584 27218 22596
rect 27249 22593 27261 22596
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 29178 22584 29184 22636
rect 29236 22624 29242 22636
rect 29365 22627 29423 22633
rect 29365 22624 29377 22627
rect 29236 22596 29377 22624
rect 29236 22584 29242 22596
rect 29365 22593 29377 22596
rect 29411 22624 29423 22627
rect 30653 22627 30711 22633
rect 30653 22624 30665 22627
rect 29411 22596 30665 22624
rect 29411 22593 29423 22596
rect 29365 22587 29423 22593
rect 30653 22593 30665 22596
rect 30699 22593 30711 22627
rect 31864 22624 31892 22720
rect 34256 22692 34284 22732
rect 35250 22692 35256 22704
rect 32370 22664 34284 22692
rect 34992 22664 35256 22692
rect 32370 22624 32398 22664
rect 32490 22624 32496 22636
rect 30653 22587 30711 22593
rect 30760 22596 31892 22624
rect 32324 22596 32398 22624
rect 32451 22596 32496 22624
rect 14642 22516 14648 22568
rect 14700 22556 14706 22568
rect 14788 22559 14846 22565
rect 14788 22556 14800 22559
rect 14700 22528 14800 22556
rect 14700 22516 14706 22528
rect 14788 22525 14800 22528
rect 14834 22556 14846 22559
rect 30377 22559 30435 22565
rect 14834 22528 15332 22556
rect 14834 22525 14846 22528
rect 14788 22519 14846 22525
rect 15304 22432 15332 22528
rect 30377 22525 30389 22559
rect 30423 22556 30435 22559
rect 30760 22556 30788 22596
rect 30423 22528 30788 22556
rect 30872 22559 30930 22565
rect 30423 22525 30435 22528
rect 30377 22519 30435 22525
rect 30872 22525 30884 22559
rect 30918 22525 30930 22559
rect 32324 22556 32352 22596
rect 32490 22584 32496 22596
rect 32548 22584 32554 22636
rect 32674 22584 32680 22636
rect 32732 22624 32738 22636
rect 34992 22633 35020 22664
rect 35250 22652 35256 22664
rect 35308 22652 35314 22704
rect 35342 22652 35348 22704
rect 35400 22692 35406 22704
rect 35529 22695 35587 22701
rect 35529 22692 35541 22695
rect 35400 22664 35541 22692
rect 35400 22652 35406 22664
rect 35529 22661 35541 22664
rect 35575 22661 35587 22695
rect 35636 22692 35664 22732
rect 36630 22720 36636 22732
rect 36688 22760 36694 22772
rect 38194 22760 38200 22772
rect 36688 22732 38200 22760
rect 36688 22720 36694 22732
rect 38194 22720 38200 22732
rect 38252 22720 38258 22772
rect 38930 22760 38936 22772
rect 38891 22732 38936 22760
rect 38930 22720 38936 22732
rect 38988 22720 38994 22772
rect 39945 22763 40003 22769
rect 39945 22729 39957 22763
rect 39991 22760 40003 22763
rect 40034 22760 40040 22772
rect 39991 22732 40040 22760
rect 39991 22729 40003 22732
rect 39945 22723 40003 22729
rect 37734 22692 37740 22704
rect 35636 22664 37740 22692
rect 35529 22655 35587 22661
rect 37734 22652 37740 22664
rect 37792 22692 37798 22704
rect 38105 22695 38163 22701
rect 38105 22692 38117 22695
rect 37792 22664 38117 22692
rect 37792 22652 37798 22664
rect 38105 22661 38117 22664
rect 38151 22661 38163 22695
rect 38105 22655 38163 22661
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 32732 22596 32781 22624
rect 32732 22584 32738 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32769 22587 32827 22593
rect 34977 22627 35035 22633
rect 34977 22593 34989 22627
rect 35023 22593 35035 22627
rect 37182 22624 37188 22636
rect 37143 22596 37188 22624
rect 34977 22587 35035 22593
rect 37182 22584 37188 22596
rect 37240 22584 37246 22636
rect 37274 22584 37280 22636
rect 37332 22624 37338 22636
rect 37461 22627 37519 22633
rect 37461 22624 37473 22627
rect 37332 22596 37473 22624
rect 37332 22584 37338 22596
rect 37461 22593 37473 22596
rect 37507 22593 37519 22627
rect 37461 22587 37519 22593
rect 30872 22519 30930 22525
rect 31312 22528 32352 22556
rect 39460 22559 39518 22565
rect 15654 22448 15660 22500
rect 15712 22488 15718 22500
rect 15841 22491 15899 22497
rect 15841 22488 15853 22491
rect 15712 22460 15853 22488
rect 15712 22448 15718 22460
rect 15841 22457 15853 22460
rect 15887 22457 15899 22491
rect 15841 22451 15899 22457
rect 15286 22420 15292 22432
rect 15247 22392 15292 22420
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 15856 22420 15884 22451
rect 15930 22448 15936 22500
rect 15988 22488 15994 22500
rect 15988 22460 16033 22488
rect 15988 22448 15994 22460
rect 17954 22448 17960 22500
rect 18012 22488 18018 22500
rect 18141 22491 18199 22497
rect 18141 22488 18153 22491
rect 18012 22460 18153 22488
rect 18012 22448 18018 22460
rect 18141 22457 18153 22460
rect 18187 22457 18199 22491
rect 18141 22451 18199 22457
rect 18233 22491 18291 22497
rect 18233 22457 18245 22491
rect 18279 22488 18291 22491
rect 18322 22488 18328 22500
rect 18279 22460 18328 22488
rect 18279 22457 18291 22460
rect 18233 22451 18291 22457
rect 16761 22423 16819 22429
rect 16761 22420 16773 22423
rect 15856 22392 16773 22420
rect 16761 22389 16773 22392
rect 16807 22389 16819 22423
rect 18156 22420 18184 22451
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 19610 22448 19616 22500
rect 19668 22448 19674 22500
rect 20070 22488 20076 22500
rect 20031 22460 20076 22488
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 20162 22448 20168 22500
rect 20220 22488 20226 22500
rect 22094 22488 22100 22500
rect 20220 22460 20265 22488
rect 22055 22460 22100 22488
rect 20220 22448 20226 22460
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 22186 22448 22192 22500
rect 22244 22488 22250 22500
rect 22244 22460 22289 22488
rect 22244 22448 22250 22460
rect 23474 22448 23480 22500
rect 23532 22488 23538 22500
rect 23937 22491 23995 22497
rect 23937 22488 23949 22491
rect 23532 22460 23949 22488
rect 23532 22448 23538 22460
rect 23937 22457 23949 22460
rect 23983 22488 23995 22491
rect 24302 22488 24308 22500
rect 23983 22460 24308 22488
rect 23983 22457 23995 22460
rect 23937 22451 23995 22457
rect 24302 22448 24308 22460
rect 24360 22448 24366 22500
rect 24486 22488 24492 22500
rect 24447 22460 24492 22488
rect 24486 22448 24492 22460
rect 24544 22448 24550 22500
rect 25406 22488 25412 22500
rect 25367 22460 25412 22488
rect 25406 22448 25412 22460
rect 25464 22448 25470 22500
rect 25501 22491 25559 22497
rect 25501 22457 25513 22491
rect 25547 22488 25559 22491
rect 25590 22488 25596 22500
rect 25547 22460 25596 22488
rect 25547 22457 25559 22460
rect 25501 22451 25559 22457
rect 25590 22448 25596 22460
rect 25648 22448 25654 22500
rect 27065 22491 27123 22497
rect 27065 22488 27077 22491
rect 26712 22460 27077 22488
rect 19061 22423 19119 22429
rect 19061 22420 19073 22423
rect 18156 22392 19073 22420
rect 16761 22383 16819 22389
rect 19061 22389 19073 22392
rect 19107 22389 19119 22423
rect 19628 22420 19656 22448
rect 19705 22423 19763 22429
rect 19705 22420 19717 22423
rect 19628 22392 19717 22420
rect 19061 22383 19119 22389
rect 19705 22389 19717 22392
rect 19751 22420 19763 22423
rect 20346 22420 20352 22432
rect 19751 22392 20352 22420
rect 19751 22389 19763 22392
rect 19705 22383 19763 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 25608 22420 25636 22448
rect 26712 22429 26740 22460
rect 27065 22457 27077 22460
rect 27111 22457 27123 22491
rect 27065 22451 27123 22457
rect 29089 22491 29147 22497
rect 29089 22457 29101 22491
rect 29135 22488 29147 22491
rect 29457 22491 29515 22497
rect 29457 22488 29469 22491
rect 29135 22460 29469 22488
rect 29135 22457 29147 22460
rect 29089 22451 29147 22457
rect 29457 22457 29469 22460
rect 29503 22488 29515 22491
rect 29638 22488 29644 22500
rect 29503 22460 29644 22488
rect 29503 22457 29515 22460
rect 29457 22451 29515 22457
rect 29638 22448 29644 22460
rect 29696 22488 29702 22500
rect 30392 22488 30420 22519
rect 29696 22460 30420 22488
rect 29696 22448 29702 22460
rect 30742 22448 30748 22500
rect 30800 22488 30806 22500
rect 30887 22488 30915 22519
rect 31312 22497 31340 22528
rect 39460 22525 39472 22559
rect 39506 22556 39518 22559
rect 39960 22556 39988 22723
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 43990 22760 43996 22772
rect 43951 22732 43996 22760
rect 43990 22720 43996 22732
rect 44048 22720 44054 22772
rect 42702 22652 42708 22704
rect 42760 22692 42766 22704
rect 42797 22695 42855 22701
rect 42797 22692 42809 22695
rect 42760 22664 42809 22692
rect 42760 22652 42766 22664
rect 42797 22661 42809 22664
rect 42843 22692 42855 22695
rect 43162 22692 43168 22704
rect 42843 22664 43168 22692
rect 42843 22661 42855 22664
rect 42797 22655 42855 22661
rect 43162 22652 43168 22664
rect 43220 22652 43226 22704
rect 43070 22624 43076 22636
rect 42983 22596 43076 22624
rect 43070 22584 43076 22596
rect 43128 22624 43134 22636
rect 46247 22627 46305 22633
rect 46247 22624 46259 22627
rect 43128 22596 46259 22624
rect 43128 22584 43134 22596
rect 46247 22593 46259 22596
rect 46293 22593 46305 22627
rect 46247 22587 46305 22593
rect 39506 22528 39988 22556
rect 39506 22525 39518 22528
rect 39460 22519 39518 22525
rect 40218 22516 40224 22568
rect 40276 22556 40282 22568
rect 41392 22559 41450 22565
rect 41392 22556 41404 22559
rect 40276 22528 41404 22556
rect 40276 22516 40282 22528
rect 41392 22525 41404 22528
rect 41438 22556 41450 22559
rect 41785 22559 41843 22565
rect 41785 22556 41797 22559
rect 41438 22528 41797 22556
rect 41438 22525 41450 22528
rect 41392 22519 41450 22525
rect 41785 22525 41797 22528
rect 41831 22525 41843 22559
rect 41785 22519 41843 22525
rect 44450 22516 44456 22568
rect 44508 22556 44514 22568
rect 44580 22559 44638 22565
rect 44580 22556 44592 22559
rect 44508 22528 44592 22556
rect 44508 22516 44514 22528
rect 44580 22525 44592 22528
rect 44626 22556 44638 22559
rect 45373 22559 45431 22565
rect 45373 22556 45385 22559
rect 44626 22528 45385 22556
rect 44626 22525 44638 22528
rect 44580 22519 44638 22525
rect 45373 22525 45385 22528
rect 45419 22525 45431 22559
rect 45373 22519 45431 22525
rect 45830 22516 45836 22568
rect 45888 22556 45894 22568
rect 46144 22559 46202 22565
rect 46144 22556 46156 22559
rect 45888 22528 46156 22556
rect 45888 22516 45894 22528
rect 46144 22525 46156 22528
rect 46190 22556 46202 22559
rect 46569 22559 46627 22565
rect 46569 22556 46581 22559
rect 46190 22528 46581 22556
rect 46190 22525 46202 22528
rect 46144 22519 46202 22525
rect 46569 22525 46581 22528
rect 46615 22525 46627 22559
rect 46569 22519 46627 22525
rect 31297 22491 31355 22497
rect 31297 22488 31309 22491
rect 30800 22460 31309 22488
rect 30800 22448 30806 22460
rect 31297 22457 31309 22460
rect 31343 22457 31355 22491
rect 31297 22451 31355 22457
rect 32585 22491 32643 22497
rect 32585 22457 32597 22491
rect 32631 22488 32643 22491
rect 34701 22491 34759 22497
rect 32631 22460 33134 22488
rect 32631 22457 32643 22460
rect 32585 22451 32643 22457
rect 33106 22432 33134 22460
rect 34701 22457 34713 22491
rect 34747 22488 34759 22491
rect 34790 22488 34796 22500
rect 34747 22460 34796 22488
rect 34747 22457 34759 22460
rect 34701 22451 34759 22457
rect 34790 22448 34796 22460
rect 34848 22488 34854 22500
rect 35069 22491 35127 22497
rect 35069 22488 35081 22491
rect 34848 22460 35081 22488
rect 34848 22448 34854 22460
rect 35069 22457 35081 22460
rect 35115 22488 35127 22491
rect 35802 22488 35808 22500
rect 35115 22460 35808 22488
rect 35115 22457 35127 22460
rect 35069 22451 35127 22457
rect 35802 22448 35808 22460
rect 35860 22448 35866 22500
rect 37001 22491 37059 22497
rect 37001 22457 37013 22491
rect 37047 22488 37059 22491
rect 37277 22491 37335 22497
rect 37277 22488 37289 22491
rect 37047 22460 37289 22488
rect 37047 22457 37059 22460
rect 37001 22451 37059 22457
rect 37277 22457 37289 22460
rect 37323 22488 37335 22491
rect 37826 22488 37832 22500
rect 37323 22460 37832 22488
rect 37323 22457 37335 22460
rect 37277 22451 37335 22457
rect 37826 22448 37832 22460
rect 37884 22448 37890 22500
rect 39666 22488 39672 22500
rect 37936 22460 39672 22488
rect 26697 22423 26755 22429
rect 26697 22420 26709 22423
rect 25608 22392 26709 22420
rect 26697 22389 26709 22392
rect 26743 22389 26755 22423
rect 28534 22420 28540 22432
rect 28495 22392 28540 22420
rect 26697 22383 26755 22389
rect 28534 22380 28540 22392
rect 28592 22380 28598 22432
rect 33042 22380 33048 22432
rect 33100 22420 33134 22432
rect 33413 22423 33471 22429
rect 33413 22420 33425 22423
rect 33100 22392 33425 22420
rect 33100 22380 33106 22392
rect 33413 22389 33425 22392
rect 33459 22389 33471 22423
rect 34146 22420 34152 22432
rect 34107 22392 34152 22420
rect 33413 22383 33471 22389
rect 34146 22380 34152 22392
rect 34204 22380 34210 22432
rect 35986 22420 35992 22432
rect 35947 22392 35992 22420
rect 35986 22380 35992 22392
rect 36044 22380 36050 22432
rect 37550 22380 37556 22432
rect 37608 22420 37614 22432
rect 37936 22420 37964 22460
rect 39666 22448 39672 22460
rect 39724 22488 39730 22500
rect 40862 22488 40868 22500
rect 39724 22460 40868 22488
rect 39724 22448 39730 22460
rect 40862 22448 40868 22460
rect 40920 22448 40926 22500
rect 43162 22448 43168 22500
rect 43220 22488 43226 22500
rect 43717 22491 43775 22497
rect 43220 22460 43265 22488
rect 43220 22448 43226 22460
rect 43717 22457 43729 22491
rect 43763 22488 43775 22491
rect 45186 22488 45192 22500
rect 43763 22460 45192 22488
rect 43763 22457 43775 22460
rect 43717 22451 43775 22457
rect 45186 22448 45192 22460
rect 45244 22448 45250 22500
rect 39298 22420 39304 22432
rect 37608 22392 37964 22420
rect 39259 22392 39304 22420
rect 37608 22380 37614 22392
rect 39298 22380 39304 22392
rect 39356 22380 39362 22432
rect 39531 22423 39589 22429
rect 39531 22389 39543 22423
rect 39577 22420 39589 22423
rect 40770 22420 40776 22432
rect 39577 22392 40776 22420
rect 39577 22389 39589 22392
rect 39531 22383 39589 22389
rect 40770 22380 40776 22392
rect 40828 22380 40834 22432
rect 41463 22423 41521 22429
rect 41463 22389 41475 22423
rect 41509 22420 41521 22423
rect 41598 22420 41604 22432
rect 41509 22392 41604 22420
rect 41509 22389 41521 22392
rect 41463 22383 41521 22389
rect 41598 22380 41604 22392
rect 41656 22380 41662 22432
rect 43438 22380 43444 22432
rect 43496 22420 43502 22432
rect 44683 22423 44741 22429
rect 44683 22420 44695 22423
rect 43496 22392 44695 22420
rect 43496 22380 43502 22392
rect 44683 22389 44695 22392
rect 44729 22389 44741 22423
rect 45002 22420 45008 22432
rect 44963 22392 45008 22420
rect 44683 22383 44741 22389
rect 45002 22380 45008 22392
rect 45060 22380 45066 22432
rect 1104 22330 48852 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 48852 22330
rect 1104 22256 48852 22278
rect 15838 22216 15844 22228
rect 15799 22188 15844 22216
rect 15838 22176 15844 22188
rect 15896 22176 15902 22228
rect 16114 22216 16120 22228
rect 16075 22188 16120 22216
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 18003 22219 18061 22225
rect 18003 22185 18015 22219
rect 18049 22216 18061 22219
rect 18138 22216 18144 22228
rect 18049 22188 18144 22216
rect 18049 22185 18061 22188
rect 18003 22179 18061 22185
rect 18138 22176 18144 22188
rect 18196 22216 18202 22228
rect 18325 22219 18383 22225
rect 18325 22216 18337 22219
rect 18196 22188 18337 22216
rect 18196 22176 18202 22188
rect 18325 22185 18337 22188
rect 18371 22185 18383 22219
rect 20162 22216 20168 22228
rect 18325 22179 18383 22185
rect 19444 22188 20168 22216
rect 19444 22160 19472 22188
rect 20162 22176 20168 22188
rect 20220 22176 20226 22228
rect 21683 22219 21741 22225
rect 21683 22185 21695 22219
rect 21729 22216 21741 22219
rect 22094 22216 22100 22228
rect 21729 22188 22100 22216
rect 21729 22185 21741 22188
rect 21683 22179 21741 22185
rect 22094 22176 22100 22188
rect 22152 22176 22158 22228
rect 22462 22216 22468 22228
rect 22423 22188 22468 22216
rect 22462 22176 22468 22188
rect 22520 22176 22526 22228
rect 23290 22176 23296 22228
rect 23348 22216 23354 22228
rect 23753 22219 23811 22225
rect 23753 22216 23765 22219
rect 23348 22188 23765 22216
rect 23348 22176 23354 22188
rect 23753 22185 23765 22188
rect 23799 22216 23811 22219
rect 23934 22216 23940 22228
rect 23799 22188 23940 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 25498 22176 25504 22228
rect 25556 22216 25562 22228
rect 25685 22219 25743 22225
rect 25685 22216 25697 22219
rect 25556 22188 25697 22216
rect 25556 22176 25562 22188
rect 25685 22185 25697 22188
rect 25731 22185 25743 22219
rect 26970 22216 26976 22228
rect 26931 22188 26976 22216
rect 25685 22179 25743 22185
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 27338 22216 27344 22228
rect 27299 22188 27344 22216
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 29549 22219 29607 22225
rect 29549 22185 29561 22219
rect 29595 22216 29607 22219
rect 32490 22216 32496 22228
rect 29595 22188 30604 22216
rect 32451 22188 32496 22216
rect 29595 22185 29607 22188
rect 29549 22179 29607 22185
rect 30576 22160 30604 22188
rect 32490 22176 32496 22188
rect 32548 22176 32554 22228
rect 33042 22216 33048 22228
rect 33003 22188 33048 22216
rect 33042 22176 33048 22188
rect 33100 22176 33106 22228
rect 34790 22216 34796 22228
rect 34751 22188 34796 22216
rect 34790 22176 34796 22188
rect 34848 22176 34854 22228
rect 35161 22219 35219 22225
rect 35161 22185 35173 22219
rect 35207 22216 35219 22219
rect 35250 22216 35256 22228
rect 35207 22188 35256 22216
rect 35207 22185 35219 22188
rect 35161 22179 35219 22185
rect 35250 22176 35256 22188
rect 35308 22176 35314 22228
rect 37182 22216 37188 22228
rect 37143 22188 37188 22216
rect 37182 22176 37188 22188
rect 37240 22176 37246 22228
rect 37642 22176 37648 22228
rect 37700 22216 37706 22228
rect 40954 22216 40960 22228
rect 37700 22188 38516 22216
rect 40915 22188 40960 22216
rect 37700 22176 37706 22188
rect 15427 22151 15485 22157
rect 15427 22117 15439 22151
rect 15473 22148 15485 22151
rect 16666 22148 16672 22160
rect 15473 22120 16672 22148
rect 15473 22117 15485 22120
rect 15427 22111 15485 22117
rect 16666 22108 16672 22120
rect 16724 22108 16730 22160
rect 19426 22148 19432 22160
rect 19387 22120 19432 22148
rect 19426 22108 19432 22120
rect 19484 22108 19490 22160
rect 19978 22148 19984 22160
rect 19939 22120 19984 22148
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 22741 22151 22799 22157
rect 22741 22117 22753 22151
rect 22787 22148 22799 22151
rect 23014 22148 23020 22160
rect 22787 22120 23020 22148
rect 22787 22117 22799 22120
rect 22741 22111 22799 22117
rect 23014 22108 23020 22120
rect 23072 22148 23078 22160
rect 24302 22148 24308 22160
rect 23072 22120 24308 22148
rect 23072 22108 23078 22120
rect 24302 22108 24308 22120
rect 24360 22108 24366 22160
rect 25406 22108 25412 22160
rect 25464 22148 25470 22160
rect 27663 22151 27721 22157
rect 27663 22148 27675 22151
rect 25464 22120 27675 22148
rect 25464 22108 25470 22120
rect 27663 22117 27675 22120
rect 27709 22117 27721 22151
rect 27663 22111 27721 22117
rect 28626 22108 28632 22160
rect 28684 22148 28690 22160
rect 28950 22151 29008 22157
rect 28950 22148 28962 22151
rect 28684 22120 28962 22148
rect 28684 22108 28690 22120
rect 28950 22117 28962 22120
rect 28996 22117 29008 22151
rect 30558 22148 30564 22160
rect 30471 22120 30564 22148
rect 28950 22111 29008 22117
rect 30558 22108 30564 22120
rect 30616 22108 30622 22160
rect 34235 22151 34293 22157
rect 34235 22117 34247 22151
rect 34281 22148 34293 22151
rect 34514 22148 34520 22160
rect 34281 22120 34520 22148
rect 34281 22117 34293 22120
rect 34235 22111 34293 22117
rect 34514 22108 34520 22120
rect 34572 22108 34578 22160
rect 35802 22148 35808 22160
rect 35763 22120 35808 22148
rect 35802 22108 35808 22120
rect 35860 22108 35866 22160
rect 36354 22148 36360 22160
rect 36315 22120 36360 22148
rect 36354 22108 36360 22120
rect 36412 22108 36418 22160
rect 37826 22108 37832 22160
rect 37884 22148 37890 22160
rect 38488 22157 38516 22188
rect 40954 22176 40960 22188
rect 41012 22176 41018 22228
rect 43070 22216 43076 22228
rect 43031 22188 43076 22216
rect 43070 22176 43076 22188
rect 43128 22176 43134 22228
rect 43346 22176 43352 22228
rect 43404 22216 43410 22228
rect 45646 22216 45652 22228
rect 43404 22188 45652 22216
rect 43404 22176 43410 22188
rect 45646 22176 45652 22188
rect 45704 22176 45710 22228
rect 37921 22151 37979 22157
rect 37921 22148 37933 22151
rect 37884 22120 37933 22148
rect 37884 22108 37890 22120
rect 37921 22117 37933 22120
rect 37967 22117 37979 22151
rect 37921 22111 37979 22117
rect 38473 22151 38531 22157
rect 38473 22117 38485 22151
rect 38519 22117 38531 22151
rect 41414 22148 41420 22160
rect 41375 22120 41420 22148
rect 38473 22111 38531 22117
rect 41414 22108 41420 22120
rect 41472 22108 41478 22160
rect 43438 22148 43444 22160
rect 43399 22120 43444 22148
rect 43438 22108 43444 22120
rect 43496 22108 43502 22160
rect 43530 22108 43536 22160
rect 43588 22148 43594 22160
rect 45370 22148 45376 22160
rect 43588 22120 43633 22148
rect 45331 22120 45376 22148
rect 43588 22108 43594 22120
rect 45370 22108 45376 22120
rect 45428 22108 45434 22160
rect 15194 22040 15200 22092
rect 15252 22080 15258 22092
rect 15324 22083 15382 22089
rect 15324 22080 15336 22083
rect 15252 22052 15336 22080
rect 15252 22040 15258 22052
rect 15324 22049 15336 22052
rect 15370 22049 15382 22083
rect 15324 22043 15382 22049
rect 16920 22083 16978 22089
rect 16920 22049 16932 22083
rect 16966 22080 16978 22083
rect 17218 22080 17224 22092
rect 16966 22052 17224 22080
rect 16966 22049 16978 22052
rect 16920 22043 16978 22049
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 17932 22083 17990 22089
rect 17932 22049 17944 22083
rect 17978 22080 17990 22083
rect 18138 22080 18144 22092
rect 17978 22052 18144 22080
rect 17978 22049 17990 22052
rect 17932 22043 17990 22049
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 20346 22040 20352 22092
rect 20404 22080 20410 22092
rect 21612 22083 21670 22089
rect 21612 22080 21624 22083
rect 20404 22052 21624 22080
rect 20404 22040 20410 22052
rect 21612 22049 21624 22052
rect 21658 22080 21670 22083
rect 22002 22080 22008 22092
rect 21658 22052 22008 22080
rect 21658 22049 21670 22052
rect 21612 22043 21670 22049
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 26602 22089 26608 22092
rect 26580 22083 26608 22089
rect 26580 22080 26592 22083
rect 26515 22052 26592 22080
rect 26580 22049 26592 22052
rect 26660 22080 26666 22092
rect 27246 22080 27252 22092
rect 26660 22052 27252 22080
rect 26580 22043 26608 22049
rect 26602 22040 26608 22043
rect 26660 22040 26666 22052
rect 27246 22040 27252 22052
rect 27304 22040 27310 22092
rect 27430 22040 27436 22092
rect 27488 22080 27494 22092
rect 27560 22083 27618 22089
rect 27560 22080 27572 22083
rect 27488 22052 27572 22080
rect 27488 22040 27494 22052
rect 27560 22049 27572 22052
rect 27606 22049 27618 22083
rect 27560 22043 27618 22049
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 29604 22052 29837 22080
rect 29604 22040 29610 22052
rect 29825 22049 29837 22052
rect 29871 22049 29883 22083
rect 29825 22043 29883 22049
rect 31113 22083 31171 22089
rect 31113 22049 31125 22083
rect 31159 22080 31171 22083
rect 32674 22080 32680 22092
rect 31159 22052 32680 22080
rect 31159 22049 31171 22052
rect 31113 22043 31171 22049
rect 32674 22040 32680 22052
rect 32732 22040 32738 22092
rect 39206 22040 39212 22092
rect 39264 22080 39270 22092
rect 39850 22080 39856 22092
rect 39264 22052 39856 22080
rect 39264 22040 39270 22052
rect 39850 22040 39856 22052
rect 39908 22080 39914 22092
rect 40256 22083 40314 22089
rect 40256 22080 40268 22083
rect 39908 22052 40268 22080
rect 39908 22040 39914 22052
rect 40256 22049 40268 22052
rect 40302 22049 40314 22083
rect 40256 22043 40314 22049
rect 46474 22040 46480 22092
rect 46532 22080 46538 22092
rect 46750 22080 46756 22092
rect 46532 22052 46756 22080
rect 46532 22040 46538 22052
rect 46750 22040 46756 22052
rect 46808 22040 46814 22092
rect 19334 22012 19340 22024
rect 19295 21984 19340 22012
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 22012 22707 22015
rect 22738 22012 22744 22024
rect 22695 21984 22744 22012
rect 22695 21981 22707 21984
rect 22649 21975 22707 21981
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 22922 22012 22928 22024
rect 22883 21984 22928 22012
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 24210 22012 24216 22024
rect 24171 21984 24216 22012
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 24394 21972 24400 22024
rect 24452 22012 24458 22024
rect 24489 22015 24547 22021
rect 24489 22012 24501 22015
rect 24452 21984 24501 22012
rect 24452 21972 24458 21984
rect 24489 21981 24501 21984
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 25409 22015 25467 22021
rect 25409 21981 25421 22015
rect 25455 22012 25467 22015
rect 25590 22012 25596 22024
rect 25455 21984 25596 22012
rect 25455 21981 25467 21984
rect 25409 21975 25467 21981
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 28350 21972 28356 22024
rect 28408 22012 28414 22024
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 28408 21984 28641 22012
rect 28408 21972 28414 21984
rect 28629 21981 28641 21984
rect 28675 21981 28687 22015
rect 30466 22012 30472 22024
rect 30427 21984 30472 22012
rect 28629 21975 28687 21981
rect 30466 21972 30472 21984
rect 30524 21972 30530 22024
rect 32122 22012 32128 22024
rect 32083 21984 32128 22012
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 33870 22012 33876 22024
rect 33831 21984 33876 22012
rect 33870 21972 33876 21984
rect 33928 21972 33934 22024
rect 35710 22012 35716 22024
rect 35671 21984 35716 22012
rect 35710 21972 35716 21984
rect 35768 21972 35774 22024
rect 37829 22015 37887 22021
rect 37829 21981 37841 22015
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 40359 22015 40417 22021
rect 40359 21981 40371 22015
rect 40405 22012 40417 22015
rect 41046 22012 41052 22024
rect 40405 21984 41052 22012
rect 40405 21981 40417 21984
rect 40359 21975 40417 21981
rect 16991 21947 17049 21953
rect 16991 21913 17003 21947
rect 17037 21944 17049 21947
rect 20070 21944 20076 21956
rect 17037 21916 20076 21944
rect 17037 21913 17049 21916
rect 16991 21907 17049 21913
rect 20070 21904 20076 21916
rect 20128 21944 20134 21956
rect 20257 21947 20315 21953
rect 20257 21944 20269 21947
rect 20128 21916 20269 21944
rect 20128 21904 20134 21916
rect 20257 21913 20269 21916
rect 20303 21913 20315 21947
rect 27982 21944 27988 21956
rect 20257 21907 20315 21913
rect 23446 21916 27988 21944
rect 21634 21836 21640 21888
rect 21692 21876 21698 21888
rect 23446 21876 23474 21916
rect 27982 21904 27988 21916
rect 28040 21904 28046 21956
rect 21692 21848 23474 21876
rect 21692 21836 21698 21848
rect 25314 21836 25320 21888
rect 25372 21876 25378 21888
rect 26651 21879 26709 21885
rect 26651 21876 26663 21879
rect 25372 21848 26663 21876
rect 25372 21836 25378 21848
rect 26651 21845 26663 21848
rect 26697 21845 26709 21879
rect 26651 21839 26709 21845
rect 30006 21836 30012 21888
rect 30064 21876 30070 21888
rect 31573 21879 31631 21885
rect 31573 21876 31585 21879
rect 30064 21848 31585 21876
rect 30064 21836 30070 21848
rect 31573 21845 31585 21848
rect 31619 21876 31631 21879
rect 31662 21876 31668 21888
rect 31619 21848 31668 21876
rect 31619 21845 31631 21848
rect 31573 21839 31631 21845
rect 31662 21836 31668 21848
rect 31720 21836 31726 21888
rect 36722 21876 36728 21888
rect 36683 21848 36728 21876
rect 36722 21836 36728 21848
rect 36780 21836 36786 21888
rect 37458 21876 37464 21888
rect 37419 21848 37464 21876
rect 37458 21836 37464 21848
rect 37516 21876 37522 21888
rect 37844 21876 37872 21975
rect 41046 21972 41052 21984
rect 41104 22012 41110 22024
rect 41325 22015 41383 22021
rect 41325 22012 41337 22015
rect 41104 21984 41337 22012
rect 41104 21972 41110 21984
rect 41325 21981 41337 21984
rect 41371 21981 41383 22015
rect 41325 21975 41383 21981
rect 41506 21972 41512 22024
rect 41564 22012 41570 22024
rect 41601 22015 41659 22021
rect 41601 22012 41613 22015
rect 41564 21984 41613 22012
rect 41564 21972 41570 21984
rect 41601 21981 41613 21984
rect 41647 21981 41659 22015
rect 45278 22012 45284 22024
rect 45239 21984 45284 22012
rect 41601 21975 41659 21981
rect 45278 21972 45284 21984
rect 45336 21972 45342 22024
rect 45462 22012 45468 22024
rect 45388 21984 45468 22012
rect 42978 21904 42984 21956
rect 43036 21944 43042 21956
rect 43993 21947 44051 21953
rect 43993 21944 44005 21947
rect 43036 21916 44005 21944
rect 43036 21904 43042 21916
rect 43993 21913 44005 21916
rect 44039 21944 44051 21947
rect 45388 21944 45416 21984
rect 45462 21972 45468 21984
rect 45520 22012 45526 22024
rect 45557 22015 45615 22021
rect 45557 22012 45569 22015
rect 45520 21984 45569 22012
rect 45520 21972 45526 21984
rect 45557 21981 45569 21984
rect 45603 21981 45615 22015
rect 45557 21975 45615 21981
rect 44039 21916 45416 21944
rect 44039 21913 44051 21916
rect 43993 21907 44051 21913
rect 44542 21876 44548 21888
rect 37516 21848 37872 21876
rect 44503 21848 44548 21876
rect 37516 21836 37522 21848
rect 44542 21836 44548 21848
rect 44600 21836 44606 21888
rect 45738 21836 45744 21888
rect 45796 21876 45802 21888
rect 46891 21879 46949 21885
rect 46891 21876 46903 21879
rect 45796 21848 46903 21876
rect 45796 21836 45802 21848
rect 46891 21845 46903 21848
rect 46937 21845 46949 21879
rect 46891 21839 46949 21845
rect 1104 21786 48852 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 48852 21786
rect 1104 21712 48852 21734
rect 17083 21675 17141 21681
rect 17083 21641 17095 21675
rect 17129 21672 17141 21675
rect 17954 21672 17960 21684
rect 17129 21644 17960 21672
rect 17129 21641 17141 21644
rect 17083 21635 17141 21641
rect 17954 21632 17960 21644
rect 18012 21632 18018 21684
rect 18969 21675 19027 21681
rect 18969 21641 18981 21675
rect 19015 21672 19027 21675
rect 19334 21672 19340 21684
rect 19015 21644 19340 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 19334 21632 19340 21644
rect 19392 21672 19398 21684
rect 19751 21675 19809 21681
rect 19751 21672 19763 21675
rect 19392 21644 19763 21672
rect 19392 21632 19398 21644
rect 19751 21641 19763 21644
rect 19797 21641 19809 21675
rect 19751 21635 19809 21641
rect 20165 21675 20223 21681
rect 20165 21641 20177 21675
rect 20211 21672 20223 21675
rect 20254 21672 20260 21684
rect 20211 21644 20260 21672
rect 20211 21641 20223 21644
rect 20165 21635 20223 21641
rect 16071 21607 16129 21613
rect 16071 21573 16083 21607
rect 16117 21604 16129 21607
rect 19058 21604 19064 21616
rect 16117 21576 19064 21604
rect 16117 21573 16129 21576
rect 16071 21567 16129 21573
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 16482 21536 16488 21548
rect 16443 21508 16488 21536
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 19426 21536 19432 21548
rect 19383 21508 19432 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20180 21536 20208 21635
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 21223 21675 21281 21681
rect 21223 21641 21235 21675
rect 21269 21672 21281 21675
rect 22462 21672 22468 21684
rect 21269 21644 22468 21672
rect 21269 21641 21281 21644
rect 21223 21635 21281 21641
rect 22462 21632 22468 21644
rect 22520 21632 22526 21684
rect 23014 21672 23020 21684
rect 22975 21644 23020 21672
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 24302 21632 24308 21684
rect 24360 21672 24366 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24360 21644 24777 21672
rect 24360 21632 24366 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 25225 21675 25283 21681
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 25590 21672 25596 21684
rect 25271 21644 25596 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 26602 21672 26608 21684
rect 26563 21644 26608 21672
rect 26602 21632 26608 21644
rect 26660 21632 26666 21684
rect 27430 21672 27436 21684
rect 27391 21644 27436 21672
rect 27430 21632 27436 21644
rect 27488 21632 27494 21684
rect 28626 21672 28632 21684
rect 28587 21644 28632 21672
rect 28626 21632 28632 21644
rect 28684 21672 28690 21684
rect 28997 21675 29055 21681
rect 28997 21672 29009 21675
rect 28684 21644 29009 21672
rect 28684 21632 28690 21644
rect 28997 21641 29009 21644
rect 29043 21641 29055 21675
rect 30558 21672 30564 21684
rect 30519 21644 30564 21672
rect 28997 21635 29055 21641
rect 24504 21576 25728 21604
rect 24504 21548 24532 21576
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 20180 21508 22569 21536
rect 16000 21471 16058 21477
rect 16000 21437 16012 21471
rect 16046 21468 16058 21471
rect 16500 21468 16528 21496
rect 16046 21440 16528 21468
rect 17012 21471 17070 21477
rect 16046 21437 16058 21440
rect 16000 21431 16058 21437
rect 17012 21437 17024 21471
rect 17058 21468 17070 21471
rect 19680 21471 19738 21477
rect 17058 21440 17540 21468
rect 17058 21437 17070 21440
rect 17012 21431 17070 21437
rect 17512 21409 17540 21440
rect 19680 21437 19692 21471
rect 19726 21468 19738 21471
rect 20180 21468 20208 21508
rect 19726 21440 20208 21468
rect 19726 21437 19738 21440
rect 19680 21431 19738 21437
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20588 21440 21005 21468
rect 20588 21428 20594 21440
rect 20993 21437 21005 21440
rect 21039 21468 21051 21471
rect 21120 21471 21178 21477
rect 21120 21468 21132 21471
rect 21039 21440 21132 21468
rect 21039 21437 21051 21440
rect 20993 21431 21051 21437
rect 21120 21437 21132 21440
rect 21166 21437 21178 21471
rect 21542 21468 21548 21480
rect 21120 21431 21178 21437
rect 21238 21440 21548 21468
rect 17497 21403 17555 21409
rect 17497 21369 17509 21403
rect 17543 21400 17555 21403
rect 21238 21400 21266 21440
rect 21542 21428 21548 21440
rect 21600 21428 21606 21480
rect 22147 21477 22175 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 24486 21536 24492 21548
rect 24447 21508 24492 21536
rect 22557 21499 22615 21505
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21536 25467 21539
rect 25498 21536 25504 21548
rect 25455 21508 25504 21536
rect 25455 21505 25467 21508
rect 25409 21499 25467 21505
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 25700 21545 25728 21576
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 22132 21471 22190 21477
rect 22132 21437 22144 21471
rect 22178 21437 22190 21471
rect 27614 21468 27620 21480
rect 22132 21431 22190 21437
rect 26706 21440 27620 21468
rect 17543 21372 21266 21400
rect 22235 21403 22293 21409
rect 17543 21369 17555 21372
rect 17497 21363 17555 21369
rect 22235 21369 22247 21403
rect 22281 21400 22293 21403
rect 22738 21400 22744 21412
rect 22281 21372 22744 21400
rect 22281 21369 22293 21372
rect 22235 21363 22293 21369
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 23477 21403 23535 21409
rect 23477 21369 23489 21403
rect 23523 21400 23535 21403
rect 23566 21400 23572 21412
rect 23523 21372 23572 21400
rect 23523 21369 23535 21372
rect 23477 21363 23535 21369
rect 23566 21360 23572 21372
rect 23624 21400 23630 21412
rect 23845 21403 23903 21409
rect 23845 21400 23857 21403
rect 23624 21372 23857 21400
rect 23624 21360 23630 21372
rect 23845 21369 23857 21372
rect 23891 21369 23903 21403
rect 23845 21363 23903 21369
rect 23934 21360 23940 21412
rect 23992 21400 23998 21412
rect 25501 21403 25559 21409
rect 23992 21372 24037 21400
rect 23992 21360 23998 21372
rect 25501 21369 25513 21403
rect 25547 21400 25559 21403
rect 25590 21400 25596 21412
rect 25547 21372 25596 21400
rect 25547 21369 25559 21372
rect 25501 21363 25559 21369
rect 25590 21360 25596 21372
rect 25648 21360 25654 21412
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 15194 21332 15200 21344
rect 13872 21304 15200 21332
rect 13872 21292 13878 21304
rect 15194 21292 15200 21304
rect 15252 21332 15258 21344
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 15252 21304 15301 21332
rect 15252 21292 15258 21304
rect 15289 21301 15301 21304
rect 15335 21301 15347 21335
rect 15289 21295 15347 21301
rect 16853 21335 16911 21341
rect 16853 21301 16865 21335
rect 16899 21332 16911 21335
rect 17218 21332 17224 21344
rect 16899 21304 17224 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18601 21335 18659 21341
rect 18601 21332 18613 21335
rect 18196 21304 18613 21332
rect 18196 21292 18202 21304
rect 18601 21301 18613 21304
rect 18647 21332 18659 21335
rect 20530 21332 20536 21344
rect 18647 21304 20536 21332
rect 18647 21301 18659 21304
rect 18601 21295 18659 21301
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 20993 21335 21051 21341
rect 20993 21301 21005 21335
rect 21039 21332 21051 21335
rect 21545 21335 21603 21341
rect 21545 21332 21557 21335
rect 21039 21304 21557 21332
rect 21039 21301 21051 21304
rect 20993 21295 21051 21301
rect 21545 21301 21557 21304
rect 21591 21332 21603 21335
rect 21634 21332 21640 21344
rect 21591 21304 21640 21332
rect 21591 21301 21603 21304
rect 21545 21295 21603 21301
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 22002 21332 22008 21344
rect 21915 21304 22008 21332
rect 22002 21292 22008 21304
rect 22060 21332 22066 21344
rect 23658 21332 23664 21344
rect 22060 21304 23664 21332
rect 22060 21292 22066 21304
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 26706 21332 26734 21440
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 28166 21468 28172 21480
rect 28127 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 27157 21403 27215 21409
rect 27157 21369 27169 21403
rect 27203 21400 27215 21403
rect 27706 21400 27712 21412
rect 27203 21372 27712 21400
rect 27203 21369 27215 21372
rect 27157 21363 27215 21369
rect 27706 21360 27712 21372
rect 27764 21400 27770 21412
rect 28184 21400 28212 21428
rect 28350 21400 28356 21412
rect 27764 21372 28212 21400
rect 28311 21372 28356 21400
rect 27764 21360 27770 21372
rect 28350 21360 28356 21372
rect 28408 21360 28414 21412
rect 29012 21400 29040 21635
rect 30558 21632 30564 21644
rect 30616 21632 30622 21684
rect 30742 21632 30748 21684
rect 30800 21672 30806 21684
rect 32490 21672 32496 21684
rect 30800 21644 32496 21672
rect 30800 21632 30806 21644
rect 32490 21632 32496 21644
rect 32548 21672 32554 21684
rect 32585 21675 32643 21681
rect 32585 21672 32597 21675
rect 32548 21644 32597 21672
rect 32548 21632 32554 21644
rect 32585 21641 32597 21644
rect 32631 21672 32643 21675
rect 34333 21675 34391 21681
rect 34333 21672 34345 21675
rect 32631 21644 34345 21672
rect 32631 21641 32643 21644
rect 32585 21635 32643 21641
rect 34333 21641 34345 21644
rect 34379 21672 34391 21675
rect 34514 21672 34520 21684
rect 34379 21644 34520 21672
rect 34379 21641 34391 21644
rect 34333 21635 34391 21641
rect 34514 21632 34520 21644
rect 34572 21632 34578 21684
rect 35710 21672 35716 21684
rect 35671 21644 35716 21672
rect 35710 21632 35716 21644
rect 35768 21632 35774 21684
rect 35802 21632 35808 21684
rect 35860 21672 35866 21684
rect 36081 21675 36139 21681
rect 36081 21672 36093 21675
rect 35860 21644 36093 21672
rect 35860 21632 35866 21644
rect 36081 21641 36093 21644
rect 36127 21672 36139 21675
rect 37826 21672 37832 21684
rect 36127 21644 37832 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 37826 21632 37832 21644
rect 37884 21632 37890 21684
rect 38102 21632 38108 21684
rect 38160 21672 38166 21684
rect 38381 21675 38439 21681
rect 38381 21672 38393 21675
rect 38160 21644 38393 21672
rect 38160 21632 38166 21644
rect 38381 21641 38393 21644
rect 38427 21641 38439 21675
rect 39850 21672 39856 21684
rect 39811 21644 39856 21672
rect 38381 21635 38439 21641
rect 30466 21564 30472 21616
rect 30524 21604 30530 21616
rect 30837 21607 30895 21613
rect 30837 21604 30849 21607
rect 30524 21576 30849 21604
rect 30524 21564 30530 21576
rect 30837 21573 30849 21576
rect 30883 21573 30895 21607
rect 30837 21567 30895 21573
rect 31202 21564 31208 21616
rect 31260 21604 31266 21616
rect 32766 21604 32772 21616
rect 31260 21576 32772 21604
rect 31260 21564 31266 21576
rect 32766 21564 32772 21576
rect 32824 21604 32830 21616
rect 32824 21576 33134 21604
rect 32824 21564 32830 21576
rect 31662 21536 31668 21548
rect 31623 21508 31668 21536
rect 31662 21496 31668 21508
rect 31720 21496 31726 21548
rect 29270 21468 29276 21480
rect 29231 21440 29276 21468
rect 29270 21428 29276 21440
rect 29328 21428 29334 21480
rect 33106 21468 33134 21576
rect 33870 21496 33876 21548
rect 33928 21536 33934 21548
rect 33965 21539 34023 21545
rect 33965 21536 33977 21539
rect 33928 21508 33977 21536
rect 33928 21496 33934 21508
rect 33965 21505 33977 21508
rect 34011 21536 34023 21539
rect 34609 21539 34667 21545
rect 34609 21536 34621 21539
rect 34011 21508 34621 21536
rect 34011 21505 34023 21508
rect 33965 21499 34023 21505
rect 34609 21505 34621 21508
rect 34655 21505 34667 21539
rect 34609 21499 34667 21505
rect 34977 21539 35035 21545
rect 34977 21505 34989 21539
rect 35023 21536 35035 21539
rect 35728 21536 35756 21632
rect 37550 21536 37556 21548
rect 35023 21508 35756 21536
rect 35820 21508 37556 21536
rect 35023 21505 35035 21508
rect 34977 21499 35035 21505
rect 33229 21471 33287 21477
rect 33229 21468 33241 21471
rect 33106 21440 33241 21468
rect 33229 21437 33241 21440
rect 33275 21437 33287 21471
rect 33229 21431 33287 21437
rect 29594 21403 29652 21409
rect 29594 21400 29606 21403
rect 29012 21372 29606 21400
rect 29594 21369 29606 21372
rect 29640 21400 29652 21403
rect 30742 21400 30748 21412
rect 29640 21372 30748 21400
rect 29640 21369 29652 21372
rect 29594 21363 29652 21369
rect 30742 21360 30748 21372
rect 30800 21360 30806 21412
rect 31754 21360 31760 21412
rect 31812 21400 31818 21412
rect 32306 21400 32312 21412
rect 31812 21372 31857 21400
rect 32267 21372 32312 21400
rect 31812 21360 31818 21372
rect 32306 21360 32312 21372
rect 32364 21400 32370 21412
rect 32674 21400 32680 21412
rect 32364 21372 32680 21400
rect 32364 21360 32370 21372
rect 32674 21360 32680 21372
rect 32732 21360 32738 21412
rect 33137 21403 33195 21409
rect 33137 21369 33149 21403
rect 33183 21400 33195 21403
rect 33244 21400 33272 21431
rect 33318 21428 33324 21480
rect 33376 21468 33382 21480
rect 33689 21471 33747 21477
rect 33689 21468 33701 21471
rect 33376 21440 33701 21468
rect 33376 21428 33382 21440
rect 33689 21437 33701 21440
rect 33735 21468 33747 21471
rect 34146 21468 34152 21480
rect 33735 21440 34152 21468
rect 33735 21437 33747 21440
rect 33689 21431 33747 21437
rect 34146 21428 34152 21440
rect 34204 21428 34210 21480
rect 35820 21400 35848 21508
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 36633 21471 36691 21477
rect 36633 21437 36645 21471
rect 36679 21468 36691 21471
rect 36722 21468 36728 21480
rect 36679 21440 36728 21468
rect 36679 21437 36691 21440
rect 36633 21431 36691 21437
rect 36722 21428 36728 21440
rect 36780 21428 36786 21480
rect 38396 21468 38424 21635
rect 39850 21632 39856 21644
rect 39908 21632 39914 21684
rect 41414 21672 41420 21684
rect 41327 21644 41420 21672
rect 41414 21632 41420 21644
rect 41472 21672 41478 21684
rect 41785 21675 41843 21681
rect 41785 21672 41797 21675
rect 41472 21644 41797 21672
rect 41472 21632 41478 21644
rect 41785 21641 41797 21644
rect 41831 21672 41843 21675
rect 42702 21672 42708 21684
rect 41831 21644 42708 21672
rect 41831 21641 41843 21644
rect 41785 21635 41843 21641
rect 42702 21632 42708 21644
rect 42760 21672 42766 21684
rect 42760 21644 42840 21672
rect 42760 21632 42766 21644
rect 42812 21604 42840 21644
rect 43438 21632 43444 21684
rect 43496 21672 43502 21684
rect 43717 21675 43775 21681
rect 43717 21672 43729 21675
rect 43496 21644 43729 21672
rect 43496 21632 43502 21644
rect 43717 21641 43729 21644
rect 43763 21641 43775 21675
rect 43717 21635 43775 21641
rect 45278 21632 45284 21684
rect 45336 21672 45342 21684
rect 45833 21675 45891 21681
rect 45833 21672 45845 21675
rect 45336 21644 45845 21672
rect 45336 21632 45342 21644
rect 45833 21641 45845 21644
rect 45879 21672 45891 21675
rect 47259 21675 47317 21681
rect 47259 21672 47271 21675
rect 45879 21644 47271 21672
rect 45879 21641 45891 21644
rect 45833 21635 45891 21641
rect 47259 21641 47271 21644
rect 47305 21641 47317 21675
rect 47259 21635 47317 21641
rect 42886 21604 42892 21616
rect 42799 21576 42892 21604
rect 42886 21564 42892 21576
rect 42944 21604 42950 21616
rect 42944 21576 43484 21604
rect 42944 21564 42950 21576
rect 40770 21496 40776 21548
rect 40828 21536 40834 21548
rect 42334 21536 42340 21548
rect 40828 21508 42340 21536
rect 40828 21496 40834 21508
rect 42334 21496 42340 21508
rect 42392 21496 42398 21548
rect 42978 21536 42984 21548
rect 42939 21508 42984 21536
rect 42978 21496 42984 21508
rect 43036 21496 43042 21548
rect 43456 21545 43484 21576
rect 45646 21564 45652 21616
rect 45704 21604 45710 21616
rect 46750 21604 46756 21616
rect 45704 21576 46756 21604
rect 45704 21564 45710 21576
rect 46750 21564 46756 21576
rect 46808 21604 46814 21616
rect 46937 21607 46995 21613
rect 46937 21604 46949 21607
rect 46808 21576 46949 21604
rect 46808 21564 46814 21576
rect 46937 21573 46949 21576
rect 46983 21573 46995 21607
rect 46937 21567 46995 21573
rect 43441 21539 43499 21545
rect 43441 21505 43453 21539
rect 43487 21536 43499 21539
rect 43530 21536 43536 21548
rect 43487 21508 43536 21536
rect 43487 21505 43499 21508
rect 43441 21499 43499 21505
rect 43530 21496 43536 21508
rect 43588 21496 43594 21548
rect 44542 21536 44548 21548
rect 44455 21508 44548 21536
rect 44542 21496 44548 21508
rect 44600 21536 44606 21548
rect 46247 21539 46305 21545
rect 46247 21536 46259 21539
rect 44600 21508 46259 21536
rect 44600 21496 44606 21508
rect 46247 21505 46259 21508
rect 46293 21505 46305 21539
rect 46247 21499 46305 21505
rect 38565 21471 38623 21477
rect 38565 21468 38577 21471
rect 38396 21440 38577 21468
rect 38565 21437 38577 21440
rect 38611 21437 38623 21471
rect 38565 21431 38623 21437
rect 39025 21471 39083 21477
rect 39025 21437 39037 21471
rect 39071 21437 39083 21471
rect 39025 21431 39083 21437
rect 39301 21471 39359 21477
rect 39301 21437 39313 21471
rect 39347 21468 39359 21471
rect 40494 21468 40500 21480
rect 39347 21440 40500 21468
rect 39347 21437 39359 21440
rect 39301 21431 39359 21437
rect 36954 21403 37012 21409
rect 36954 21400 36966 21403
rect 33183 21372 35848 21400
rect 36464 21372 36966 21400
rect 33183 21369 33195 21372
rect 33137 21363 33195 21369
rect 30190 21332 30196 21344
rect 23808 21304 26734 21332
rect 30151 21304 30196 21332
rect 23808 21292 23814 21304
rect 30190 21292 30196 21304
rect 30248 21292 30254 21344
rect 31481 21335 31539 21341
rect 31481 21301 31493 21335
rect 31527 21332 31539 21335
rect 31772 21332 31800 21360
rect 31527 21304 31800 21332
rect 31527 21301 31539 21304
rect 31481 21295 31539 21301
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 36464 21341 36492 21372
rect 36954 21369 36966 21372
rect 37000 21400 37012 21403
rect 38010 21400 38016 21412
rect 37000 21372 38016 21400
rect 37000 21369 37012 21372
rect 36954 21363 37012 21369
rect 38010 21360 38016 21372
rect 38068 21360 38074 21412
rect 39040 21400 39068 21431
rect 40494 21428 40500 21440
rect 40552 21428 40558 21480
rect 46160 21471 46218 21477
rect 46160 21437 46172 21471
rect 46206 21468 46218 21471
rect 46206 21440 46704 21468
rect 46206 21437 46218 21440
rect 46160 21431 46218 21437
rect 39758 21400 39764 21412
rect 38626 21372 39764 21400
rect 36449 21335 36507 21341
rect 36449 21332 36461 21335
rect 34572 21304 36461 21332
rect 34572 21292 34578 21304
rect 36449 21301 36461 21304
rect 36495 21301 36507 21335
rect 37550 21332 37556 21344
rect 37511 21304 37556 21332
rect 36449 21295 36507 21301
rect 37550 21292 37556 21304
rect 37608 21292 37614 21344
rect 38105 21335 38163 21341
rect 38105 21301 38117 21335
rect 38151 21332 38163 21335
rect 38378 21332 38384 21344
rect 38151 21304 38384 21332
rect 38151 21301 38163 21304
rect 38105 21295 38163 21301
rect 38378 21292 38384 21304
rect 38436 21332 38442 21344
rect 38626 21332 38654 21372
rect 39758 21360 39764 21372
rect 39816 21360 39822 21412
rect 40818 21403 40876 21409
rect 40818 21369 40830 21403
rect 40864 21369 40876 21403
rect 40818 21363 40876 21369
rect 42429 21403 42487 21409
rect 42429 21369 42441 21403
rect 42475 21369 42487 21403
rect 42429 21363 42487 21369
rect 44361 21403 44419 21409
rect 44361 21369 44373 21403
rect 44407 21400 44419 21403
rect 44634 21400 44640 21412
rect 44407 21372 44640 21400
rect 44407 21369 44419 21372
rect 44361 21363 44419 21369
rect 40310 21332 40316 21344
rect 38436 21304 38654 21332
rect 40271 21304 40316 21332
rect 38436 21292 38442 21304
rect 40310 21292 40316 21304
rect 40368 21332 40374 21344
rect 40833 21332 40861 21363
rect 40368 21304 40861 21332
rect 40368 21292 40374 21304
rect 41414 21292 41420 21344
rect 41472 21332 41478 21344
rect 42061 21335 42119 21341
rect 42061 21332 42073 21335
rect 41472 21304 42073 21332
rect 41472 21292 41478 21304
rect 42061 21301 42073 21304
rect 42107 21332 42119 21335
rect 42444 21332 42472 21363
rect 44634 21360 44640 21372
rect 44692 21360 44698 21412
rect 45186 21400 45192 21412
rect 45147 21372 45192 21400
rect 45186 21360 45192 21372
rect 45244 21360 45250 21412
rect 42107 21304 42472 21332
rect 44652 21332 44680 21360
rect 46676 21344 46704 21440
rect 46934 21428 46940 21480
rect 46992 21468 46998 21480
rect 47188 21471 47246 21477
rect 47188 21468 47200 21471
rect 46992 21440 47200 21468
rect 46992 21428 46998 21440
rect 47188 21437 47200 21440
rect 47234 21468 47246 21471
rect 47578 21468 47584 21480
rect 47234 21440 47584 21468
rect 47234 21437 47246 21440
rect 47188 21431 47246 21437
rect 47578 21428 47584 21440
rect 47636 21428 47642 21480
rect 45370 21332 45376 21344
rect 44652 21304 45376 21332
rect 42107 21301 42119 21304
rect 42061 21295 42119 21301
rect 45370 21292 45376 21304
rect 45428 21332 45434 21344
rect 45465 21335 45523 21341
rect 45465 21332 45477 21335
rect 45428 21304 45477 21332
rect 45428 21292 45434 21304
rect 45465 21301 45477 21304
rect 45511 21301 45523 21335
rect 46658 21332 46664 21344
rect 46619 21304 46664 21332
rect 45465 21295 45523 21301
rect 46658 21292 46664 21304
rect 46716 21292 46722 21344
rect 1104 21242 48852 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 48852 21242
rect 1104 21168 48852 21190
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 17083 21131 17141 21137
rect 17083 21128 17095 21131
rect 15344 21100 17095 21128
rect 15344 21088 15350 21100
rect 17083 21097 17095 21100
rect 17129 21097 17141 21131
rect 17083 21091 17141 21097
rect 17218 21088 17224 21140
rect 17276 21128 17282 21140
rect 19242 21128 19248 21140
rect 17276 21100 19248 21128
rect 17276 21088 17282 21100
rect 19242 21088 19248 21100
rect 19300 21128 19306 21140
rect 22738 21128 22744 21140
rect 19300 21100 20116 21128
rect 22699 21100 22744 21128
rect 19300 21088 19306 21100
rect 18141 21063 18199 21069
rect 18141 21029 18153 21063
rect 18187 21060 18199 21063
rect 18966 21060 18972 21072
rect 18187 21032 18972 21060
rect 18187 21029 18199 21032
rect 18141 21023 18199 21029
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 16991 20995 17049 21001
rect 16991 20961 17003 20995
rect 17037 20961 17049 20995
rect 16991 20955 17049 20961
rect 17006 20868 17034 20955
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 19556 20995 19614 21001
rect 19556 20992 19568 20995
rect 18932 20964 19568 20992
rect 18932 20952 18938 20964
rect 19556 20961 19568 20964
rect 19602 20992 19614 20995
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19602 20964 19993 20992
rect 19602 20961 19614 20964
rect 19556 20955 19614 20961
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 20088 20992 20116 21100
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 23566 21128 23572 21140
rect 23527 21100 23572 21128
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 24210 21128 24216 21140
rect 24171 21100 24216 21128
rect 24210 21088 24216 21100
rect 24268 21088 24274 21140
rect 27614 21128 27620 21140
rect 27575 21100 27620 21128
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 28350 21088 28356 21140
rect 28408 21128 28414 21140
rect 28905 21131 28963 21137
rect 28905 21128 28917 21131
rect 28408 21100 28917 21128
rect 28408 21088 28414 21100
rect 28905 21097 28917 21100
rect 28951 21097 28963 21131
rect 28905 21091 28963 21097
rect 31941 21131 31999 21137
rect 31941 21097 31953 21131
rect 31987 21128 31999 21131
rect 32122 21128 32128 21140
rect 31987 21100 32128 21128
rect 31987 21097 31999 21100
rect 31941 21091 31999 21097
rect 32122 21088 32128 21100
rect 32180 21128 32186 21140
rect 32217 21131 32275 21137
rect 32217 21128 32229 21131
rect 32180 21100 32229 21128
rect 32180 21088 32186 21100
rect 32217 21097 32229 21100
rect 32263 21097 32275 21131
rect 32217 21091 32275 21097
rect 32582 21088 32588 21140
rect 32640 21128 32646 21140
rect 37461 21131 37519 21137
rect 32640 21100 33134 21128
rect 32640 21088 32646 21100
rect 22419 21063 22477 21069
rect 22419 21029 22431 21063
rect 22465 21060 22477 21063
rect 24228 21060 24256 21088
rect 22465 21032 24256 21060
rect 28629 21063 28687 21069
rect 22465 21029 22477 21032
rect 22419 21023 22477 21029
rect 28629 21029 28641 21063
rect 28675 21060 28687 21063
rect 29270 21060 29276 21072
rect 28675 21032 29276 21060
rect 28675 21029 28687 21032
rect 28629 21023 28687 21029
rect 29270 21020 29276 21032
rect 29328 21020 29334 21072
rect 29825 21063 29883 21069
rect 29825 21029 29837 21063
rect 29871 21060 29883 21063
rect 30190 21060 30196 21072
rect 29871 21032 30196 21060
rect 29871 21029 29883 21032
rect 29825 21023 29883 21029
rect 30190 21020 30196 21032
rect 30248 21020 30254 21072
rect 30377 21063 30435 21069
rect 30377 21029 30389 21063
rect 30423 21060 30435 21063
rect 32306 21060 32312 21072
rect 30423 21032 32312 21060
rect 30423 21029 30435 21032
rect 30377 21023 30435 21029
rect 32306 21020 32312 21032
rect 32364 21020 32370 21072
rect 32600 21060 32628 21088
rect 32416 21032 32628 21060
rect 22332 20995 22390 21001
rect 22332 20992 22344 20995
rect 20088 20964 22344 20992
rect 19981 20955 20039 20961
rect 22332 20961 22344 20964
rect 22378 20992 22390 20995
rect 22646 20992 22652 21004
rect 22378 20964 22652 20992
rect 22378 20961 22390 20964
rect 22332 20955 22390 20961
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 25409 20995 25467 21001
rect 25409 20961 25421 20995
rect 25455 20992 25467 20995
rect 25866 20992 25872 21004
rect 25455 20964 25872 20992
rect 25455 20961 25467 20964
rect 25409 20955 25467 20961
rect 25866 20952 25872 20964
rect 25924 20992 25930 21004
rect 26548 20995 26606 21001
rect 26548 20992 26560 20995
rect 25924 20964 26560 20992
rect 25924 20952 25930 20964
rect 26548 20961 26560 20964
rect 26594 20961 26606 20995
rect 26548 20955 26606 20961
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 28074 20992 28080 21004
rect 27120 20964 28080 20992
rect 27120 20952 27126 20964
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 28166 20952 28172 21004
rect 28224 20992 28230 21004
rect 32416 21001 32444 21032
rect 28445 20995 28503 21001
rect 28445 20992 28457 20995
rect 28224 20964 28457 20992
rect 28224 20952 28230 20964
rect 28445 20961 28457 20964
rect 28491 20992 28503 20995
rect 32401 20995 32459 21001
rect 28491 20964 28994 20992
rect 28491 20961 28503 20964
rect 28445 20955 28503 20961
rect 17494 20884 17500 20936
rect 17552 20924 17558 20936
rect 18046 20924 18052 20936
rect 17552 20896 18052 20924
rect 17552 20884 17558 20896
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18690 20924 18696 20936
rect 18651 20896 18696 20924
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 21266 20924 21272 20936
rect 21227 20896 21272 20924
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 16942 20816 16948 20868
rect 17000 20828 17034 20868
rect 25593 20859 25651 20865
rect 17000 20816 17006 20828
rect 25593 20825 25605 20859
rect 25639 20856 25651 20859
rect 27706 20856 27712 20868
rect 25639 20828 27712 20856
rect 25639 20825 25651 20828
rect 25593 20819 25651 20825
rect 27706 20816 27712 20828
rect 27764 20816 27770 20868
rect 28966 20856 28994 20964
rect 32401 20961 32413 20995
rect 32447 20961 32459 20995
rect 32674 20992 32680 21004
rect 32635 20964 32680 20992
rect 32401 20955 32459 20961
rect 32674 20952 32680 20964
rect 32732 20952 32738 21004
rect 33106 20992 33134 21100
rect 37461 21097 37473 21131
rect 37507 21128 37519 21131
rect 37826 21128 37832 21140
rect 37507 21100 37832 21128
rect 37507 21097 37519 21100
rect 37461 21091 37519 21097
rect 37826 21088 37832 21100
rect 37884 21088 37890 21140
rect 40494 21128 40500 21140
rect 40455 21100 40500 21128
rect 40494 21088 40500 21100
rect 40552 21088 40558 21140
rect 41046 21128 41052 21140
rect 41007 21100 41052 21128
rect 41046 21088 41052 21100
rect 41104 21088 41110 21140
rect 42334 21128 42340 21140
rect 42295 21100 42340 21128
rect 42334 21088 42340 21100
rect 42392 21088 42398 21140
rect 44634 21088 44640 21140
rect 44692 21128 44698 21140
rect 44821 21131 44879 21137
rect 44821 21128 44833 21131
rect 44692 21100 44833 21128
rect 44692 21088 44698 21100
rect 44821 21097 44833 21100
rect 44867 21128 44879 21131
rect 44867 21100 45876 21128
rect 44867 21097 44879 21100
rect 44821 21091 44879 21097
rect 45848 21072 45876 21100
rect 35894 21020 35900 21072
rect 35952 21060 35958 21072
rect 35989 21063 36047 21069
rect 35989 21060 36001 21063
rect 35952 21032 36001 21060
rect 35952 21020 35958 21032
rect 35989 21029 36001 21032
rect 36035 21029 36047 21063
rect 35989 21023 36047 21029
rect 37550 21020 37556 21072
rect 37608 21060 37614 21072
rect 37921 21063 37979 21069
rect 37921 21060 37933 21063
rect 37608 21032 37933 21060
rect 37608 21020 37614 21032
rect 37921 21029 37933 21032
rect 37967 21029 37979 21063
rect 41414 21060 41420 21072
rect 41375 21032 41420 21060
rect 37921 21023 37979 21029
rect 41414 21020 41420 21032
rect 41472 21020 41478 21072
rect 43990 21020 43996 21072
rect 44048 21060 44054 21072
rect 44222 21063 44280 21069
rect 44222 21060 44234 21063
rect 44048 21032 44234 21060
rect 44048 21020 44054 21032
rect 44222 21029 44234 21032
rect 44268 21029 44280 21063
rect 44222 21023 44280 21029
rect 45370 21020 45376 21072
rect 45428 21060 45434 21072
rect 45554 21060 45560 21072
rect 45428 21032 45560 21060
rect 45428 21020 45434 21032
rect 45554 21020 45560 21032
rect 45612 21020 45618 21072
rect 45738 21060 45744 21072
rect 45699 21032 45744 21060
rect 45738 21020 45744 21032
rect 45796 21020 45802 21072
rect 45830 21020 45836 21072
rect 45888 21060 45894 21072
rect 45888 21032 45981 21060
rect 45888 21020 45894 21032
rect 34146 20992 34152 21004
rect 33106 20964 34152 20992
rect 34146 20952 34152 20964
rect 34204 20952 34210 21004
rect 34609 20995 34667 21001
rect 34609 20961 34621 20995
rect 34655 20992 34667 20995
rect 35250 20992 35256 21004
rect 34655 20964 35256 20992
rect 34655 20961 34667 20964
rect 34609 20955 34667 20961
rect 35250 20952 35256 20964
rect 35308 20952 35314 21004
rect 39022 20952 39028 21004
rect 39080 20992 39086 21004
rect 39301 20995 39359 21001
rect 39301 20992 39313 20995
rect 39080 20964 39313 20992
rect 39080 20952 39086 20964
rect 39301 20961 39313 20964
rect 39347 20961 39359 20995
rect 39758 20992 39764 21004
rect 39719 20964 39764 20992
rect 39301 20955 39359 20961
rect 39758 20952 39764 20964
rect 39816 20952 39822 21004
rect 42061 20995 42119 21001
rect 42061 20961 42073 20995
rect 42107 20992 42119 20995
rect 42107 20964 45600 20992
rect 42107 20961 42119 20964
rect 42061 20955 42119 20961
rect 45572 20936 45600 20964
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20924 29791 20927
rect 29822 20924 29828 20936
rect 29779 20896 29828 20924
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 34790 20924 34796 20936
rect 34703 20896 34796 20924
rect 34790 20884 34796 20896
rect 34848 20924 34854 20936
rect 35069 20927 35127 20933
rect 35069 20924 35081 20927
rect 34848 20896 35081 20924
rect 34848 20884 34854 20896
rect 35069 20893 35081 20896
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35897 20927 35955 20933
rect 35897 20893 35909 20927
rect 35943 20924 35955 20927
rect 36354 20924 36360 20936
rect 35943 20896 36360 20924
rect 35943 20893 35955 20896
rect 35897 20887 35955 20893
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 37274 20884 37280 20936
rect 37332 20924 37338 20936
rect 37829 20927 37887 20933
rect 37829 20924 37841 20927
rect 37332 20896 37841 20924
rect 37332 20884 37338 20896
rect 37829 20893 37841 20896
rect 37875 20924 37887 20927
rect 38102 20924 38108 20936
rect 37875 20896 38108 20924
rect 37875 20893 37887 20896
rect 37829 20887 37887 20893
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 38194 20884 38200 20936
rect 38252 20924 38258 20936
rect 40037 20927 40095 20933
rect 38252 20896 38297 20924
rect 38252 20884 38258 20896
rect 40037 20893 40049 20927
rect 40083 20924 40095 20927
rect 41322 20924 41328 20936
rect 40083 20896 40861 20924
rect 41283 20896 41328 20924
rect 40083 20893 40095 20896
rect 40037 20887 40095 20893
rect 30926 20856 30932 20868
rect 28966 20828 30932 20856
rect 30926 20816 30932 20828
rect 30984 20816 30990 20868
rect 36449 20859 36507 20865
rect 36449 20825 36461 20859
rect 36495 20856 36507 20859
rect 38212 20856 38240 20884
rect 36495 20828 38240 20856
rect 40833 20856 40861 20896
rect 41322 20884 41328 20896
rect 41380 20884 41386 20936
rect 43901 20927 43959 20933
rect 43901 20924 43913 20927
rect 41432 20896 43913 20924
rect 41432 20856 41460 20896
rect 43901 20893 43913 20896
rect 43947 20924 43959 20927
rect 44358 20924 44364 20936
rect 43947 20896 44364 20924
rect 43947 20893 43959 20896
rect 43901 20887 43959 20893
rect 44358 20884 44364 20896
rect 44416 20884 44422 20936
rect 45554 20884 45560 20936
rect 45612 20924 45618 20936
rect 46017 20927 46075 20933
rect 46017 20924 46029 20927
rect 45612 20896 46029 20924
rect 45612 20884 45618 20896
rect 46017 20893 46029 20896
rect 46063 20893 46075 20927
rect 46017 20887 46075 20893
rect 40833 20828 41460 20856
rect 36495 20825 36507 20828
rect 36449 20819 36507 20825
rect 41506 20816 41512 20868
rect 41564 20856 41570 20868
rect 41877 20859 41935 20865
rect 41877 20856 41889 20859
rect 41564 20828 41889 20856
rect 41564 20816 41570 20828
rect 41877 20825 41889 20828
rect 41923 20856 41935 20859
rect 42061 20859 42119 20865
rect 42061 20856 42073 20859
rect 41923 20828 42073 20856
rect 41923 20825 41935 20828
rect 41877 20819 41935 20825
rect 42061 20825 42073 20828
rect 42107 20825 42119 20859
rect 42061 20819 42119 20825
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 19659 20791 19717 20797
rect 19659 20788 19671 20791
rect 18840 20760 19671 20788
rect 18840 20748 18846 20760
rect 19659 20757 19671 20760
rect 19705 20757 19717 20791
rect 19659 20751 19717 20757
rect 26510 20748 26516 20800
rect 26568 20788 26574 20800
rect 26651 20791 26709 20797
rect 26651 20788 26663 20791
rect 26568 20760 26663 20788
rect 26568 20748 26574 20760
rect 26651 20757 26663 20760
rect 26697 20757 26709 20791
rect 31018 20788 31024 20800
rect 30979 20760 31024 20788
rect 26651 20751 26709 20757
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 33318 20788 33324 20800
rect 33279 20760 33324 20788
rect 33318 20748 33324 20760
rect 33376 20748 33382 20800
rect 38930 20788 38936 20800
rect 38891 20760 38936 20788
rect 38930 20748 38936 20760
rect 38988 20748 38994 20800
rect 44726 20748 44732 20800
rect 44784 20788 44790 20800
rect 46842 20788 46848 20800
rect 44784 20760 46848 20788
rect 44784 20748 44790 20760
rect 46842 20748 46848 20760
rect 46900 20748 46906 20800
rect 1104 20698 48852 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 48852 20698
rect 1104 20624 48852 20646
rect 17126 20544 17132 20596
rect 17184 20584 17190 20596
rect 17221 20587 17279 20593
rect 17221 20584 17233 20587
rect 17184 20556 17233 20584
rect 17184 20544 17190 20556
rect 17221 20553 17233 20556
rect 17267 20553 17279 20587
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 17221 20547 17279 20553
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 17770 20584 17776 20596
rect 17731 20556 17776 20584
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18966 20584 18972 20596
rect 18927 20556 18972 20584
rect 18966 20544 18972 20556
rect 19024 20584 19030 20596
rect 19245 20587 19303 20593
rect 19245 20584 19257 20587
rect 19024 20556 19257 20584
rect 19024 20544 19030 20556
rect 19245 20553 19257 20556
rect 19291 20553 19303 20587
rect 19245 20547 19303 20553
rect 21266 20544 21272 20596
rect 21324 20584 21330 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 21324 20556 21373 20584
rect 21324 20544 21330 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 22646 20584 22652 20596
rect 22607 20556 22652 20584
rect 21361 20547 21419 20553
rect 16853 20519 16911 20525
rect 16853 20485 16865 20519
rect 16899 20516 16911 20519
rect 16942 20516 16948 20528
rect 16899 20488 16948 20516
rect 16899 20485 16911 20488
rect 16853 20479 16911 20485
rect 16942 20476 16948 20488
rect 17000 20516 17006 20528
rect 18690 20516 18696 20528
rect 17000 20488 18696 20516
rect 17000 20476 17006 20488
rect 18690 20476 18696 20488
rect 18748 20476 18754 20528
rect 21376 20448 21404 20547
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 25866 20584 25872 20596
rect 25827 20556 25872 20584
rect 25866 20544 25872 20556
rect 25924 20584 25930 20596
rect 27065 20587 27123 20593
rect 27065 20584 27077 20587
rect 25924 20556 27077 20584
rect 25924 20544 25930 20556
rect 27065 20553 27077 20556
rect 27111 20553 27123 20587
rect 27065 20547 27123 20553
rect 27525 20587 27583 20593
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 28166 20584 28172 20596
rect 27571 20556 28172 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 30190 20544 30196 20596
rect 30248 20584 30254 20596
rect 30469 20587 30527 20593
rect 30469 20584 30481 20587
rect 30248 20556 30481 20584
rect 30248 20544 30254 20556
rect 30469 20553 30481 20556
rect 30515 20553 30527 20587
rect 30469 20547 30527 20553
rect 30742 20544 30748 20596
rect 30800 20584 30806 20596
rect 30837 20587 30895 20593
rect 30837 20584 30849 20587
rect 30800 20556 30849 20584
rect 30800 20544 30806 20556
rect 30837 20553 30849 20556
rect 30883 20553 30895 20587
rect 30837 20547 30895 20553
rect 31754 20544 31760 20596
rect 31812 20584 31818 20596
rect 31941 20587 31999 20593
rect 31941 20584 31953 20587
rect 31812 20556 31953 20584
rect 31812 20544 31818 20556
rect 31941 20553 31953 20556
rect 31987 20553 31999 20587
rect 31941 20547 31999 20553
rect 32309 20587 32367 20593
rect 32309 20553 32321 20587
rect 32355 20584 32367 20587
rect 32582 20584 32588 20596
rect 32355 20556 32588 20584
rect 32355 20553 32367 20556
rect 32309 20547 32367 20553
rect 32582 20544 32588 20556
rect 32640 20544 32646 20596
rect 32674 20544 32680 20596
rect 32732 20584 32738 20596
rect 32950 20584 32956 20596
rect 32732 20556 32777 20584
rect 32911 20556 32956 20584
rect 32732 20544 32738 20556
rect 32950 20544 32956 20556
rect 33008 20544 33014 20596
rect 34514 20544 34520 20596
rect 34572 20584 34578 20596
rect 34609 20587 34667 20593
rect 34609 20584 34621 20587
rect 34572 20556 34621 20584
rect 34572 20544 34578 20556
rect 34609 20553 34621 20556
rect 34655 20553 34667 20587
rect 34609 20547 34667 20553
rect 37550 20544 37556 20596
rect 37608 20584 37614 20596
rect 37737 20587 37795 20593
rect 37737 20584 37749 20587
rect 37608 20556 37749 20584
rect 37608 20544 37614 20556
rect 37737 20553 37749 20556
rect 37783 20553 37795 20587
rect 38102 20584 38108 20596
rect 38063 20556 38108 20584
rect 37737 20547 37795 20553
rect 38102 20544 38108 20556
rect 38160 20544 38166 20596
rect 38749 20587 38807 20593
rect 38749 20553 38761 20587
rect 38795 20584 38807 20587
rect 38838 20584 38844 20596
rect 38795 20556 38844 20584
rect 38795 20553 38807 20556
rect 38749 20547 38807 20553
rect 38838 20544 38844 20556
rect 38896 20544 38902 20596
rect 39022 20544 39028 20596
rect 39080 20584 39086 20596
rect 39853 20587 39911 20593
rect 39853 20584 39865 20587
rect 39080 20556 39865 20584
rect 39080 20544 39086 20556
rect 39853 20553 39865 20556
rect 39899 20553 39911 20587
rect 42886 20584 42892 20596
rect 42847 20556 42892 20584
rect 39853 20547 39911 20553
rect 42886 20544 42892 20556
rect 42944 20544 42950 20596
rect 44358 20584 44364 20596
rect 44319 20556 44364 20584
rect 44358 20544 44364 20556
rect 44416 20544 44422 20596
rect 44913 20587 44971 20593
rect 44913 20553 44925 20587
rect 44959 20584 44971 20587
rect 45738 20584 45744 20596
rect 44959 20556 45744 20584
rect 44959 20553 44971 20556
rect 44913 20547 44971 20553
rect 45738 20544 45744 20556
rect 45796 20544 45802 20596
rect 45830 20544 45836 20596
rect 45888 20584 45894 20596
rect 45888 20556 45933 20584
rect 45888 20544 45894 20556
rect 28074 20476 28080 20528
rect 28132 20516 28138 20528
rect 28721 20519 28779 20525
rect 28721 20516 28733 20519
rect 28132 20488 28733 20516
rect 28132 20476 28138 20488
rect 28721 20485 28733 20488
rect 28767 20516 28779 20519
rect 33042 20516 33048 20528
rect 28767 20488 33048 20516
rect 28767 20485 28779 20488
rect 28721 20479 28779 20485
rect 33042 20476 33048 20488
rect 33100 20476 33106 20528
rect 33318 20476 33324 20528
rect 33376 20516 33382 20528
rect 33781 20519 33839 20525
rect 33781 20516 33793 20519
rect 33376 20488 33793 20516
rect 33376 20476 33382 20488
rect 33781 20485 33793 20488
rect 33827 20516 33839 20519
rect 43990 20516 43996 20528
rect 33827 20488 35296 20516
rect 33827 20485 33839 20488
rect 33781 20479 33839 20485
rect 35268 20460 35296 20488
rect 40833 20488 43996 20516
rect 21637 20451 21695 20457
rect 21637 20448 21649 20451
rect 16995 20420 21036 20448
rect 21376 20420 21649 20448
rect 16995 20389 17023 20420
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 16980 20383 17038 20389
rect 16980 20380 16992 20383
rect 16531 20352 16992 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 16980 20349 16992 20352
rect 17026 20349 17038 20383
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 16980 20343 17038 20349
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20349 20039 20383
rect 19981 20343 20039 20349
rect 17770 20272 17776 20324
rect 17828 20312 17834 20324
rect 18370 20315 18428 20321
rect 18370 20312 18382 20315
rect 17828 20284 18382 20312
rect 17828 20272 17834 20284
rect 18370 20281 18382 20284
rect 18416 20281 18428 20315
rect 19889 20315 19947 20321
rect 19889 20312 19901 20315
rect 18370 20275 18428 20281
rect 19306 20284 19901 20312
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19306 20244 19334 20284
rect 19889 20281 19901 20284
rect 19935 20312 19947 20315
rect 19996 20312 20024 20343
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 20441 20383 20499 20389
rect 20441 20380 20453 20383
rect 20128 20352 20453 20380
rect 20128 20340 20134 20352
rect 20441 20349 20453 20352
rect 20487 20349 20499 20383
rect 20441 20343 20499 20349
rect 19935 20284 20024 20312
rect 20717 20315 20775 20321
rect 19935 20281 19947 20284
rect 19889 20275 19947 20281
rect 20717 20281 20729 20315
rect 20763 20312 20775 20315
rect 20898 20312 20904 20324
rect 20763 20284 20904 20312
rect 20763 20281 20775 20284
rect 20717 20275 20775 20281
rect 20898 20272 20904 20284
rect 20956 20272 20962 20324
rect 18288 20216 19334 20244
rect 21008 20244 21036 20420
rect 21637 20417 21649 20420
rect 21683 20417 21695 20451
rect 26878 20448 26884 20460
rect 21637 20411 21695 20417
rect 24136 20420 26884 20448
rect 24136 20389 24164 20420
rect 26878 20408 26884 20420
rect 26936 20408 26942 20460
rect 30098 20448 30104 20460
rect 29472 20420 30104 20448
rect 25130 20389 25136 20392
rect 23728 20383 23786 20389
rect 23728 20349 23740 20383
rect 23774 20380 23786 20383
rect 24121 20383 24179 20389
rect 24121 20380 24133 20383
rect 23774 20352 24133 20380
rect 23774 20349 23786 20352
rect 23728 20343 23786 20349
rect 24121 20349 24133 20352
rect 24167 20349 24179 20383
rect 25108 20383 25136 20389
rect 25108 20380 25120 20383
rect 25043 20352 25120 20380
rect 24121 20343 24179 20349
rect 25108 20349 25120 20352
rect 25188 20380 25194 20392
rect 25501 20383 25559 20389
rect 25501 20380 25513 20383
rect 25188 20352 25513 20380
rect 25108 20343 25136 20349
rect 25130 20340 25136 20343
rect 25188 20340 25194 20352
rect 25501 20349 25513 20352
rect 25547 20349 25559 20383
rect 26510 20380 26516 20392
rect 26471 20352 26516 20380
rect 25501 20343 25559 20349
rect 26510 20340 26516 20352
rect 26568 20340 26574 20392
rect 27706 20380 27712 20392
rect 27667 20352 27712 20380
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 29472 20389 29500 20420
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 31018 20448 31024 20460
rect 30979 20420 31024 20448
rect 31018 20408 31024 20420
rect 31076 20408 31082 20460
rect 33134 20448 33140 20460
rect 31128 20420 33140 20448
rect 29457 20383 29515 20389
rect 29457 20349 29469 20383
rect 29503 20349 29515 20383
rect 31128 20380 31156 20420
rect 33134 20408 33140 20420
rect 33192 20408 33198 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 34885 20451 34943 20457
rect 34885 20448 34897 20451
rect 34848 20420 34897 20448
rect 34848 20408 34854 20420
rect 34885 20417 34897 20420
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 35250 20408 35256 20460
rect 35308 20448 35314 20460
rect 36173 20451 36231 20457
rect 36173 20448 36185 20451
rect 35308 20420 36185 20448
rect 35308 20408 35314 20420
rect 36173 20417 36185 20420
rect 36219 20448 36231 20451
rect 36219 20420 36860 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 36832 20392 36860 20420
rect 29457 20343 29515 20349
rect 29748 20352 31156 20380
rect 32769 20383 32827 20389
rect 21085 20315 21143 20321
rect 21085 20281 21097 20315
rect 21131 20312 21143 20315
rect 21729 20315 21787 20321
rect 21729 20312 21741 20315
rect 21131 20284 21741 20312
rect 21131 20281 21143 20284
rect 21085 20275 21143 20281
rect 21729 20281 21741 20284
rect 21775 20312 21787 20315
rect 21818 20312 21824 20324
rect 21775 20284 21824 20312
rect 21775 20281 21787 20284
rect 21729 20275 21787 20281
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 22281 20315 22339 20321
rect 22281 20281 22293 20315
rect 22327 20312 22339 20315
rect 23474 20312 23480 20324
rect 22327 20284 23480 20312
rect 22327 20281 22339 20284
rect 22281 20275 22339 20281
rect 21542 20244 21548 20256
rect 21008 20216 21548 20244
rect 18288 20204 18294 20216
rect 21542 20204 21548 20216
rect 21600 20244 21606 20256
rect 22296 20244 22324 20275
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 26050 20312 26056 20324
rect 26011 20284 26056 20312
rect 26050 20272 26056 20284
rect 26108 20272 26114 20324
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 27617 20315 27675 20321
rect 27617 20312 27629 20315
rect 27304 20284 27629 20312
rect 27304 20272 27310 20284
rect 27617 20281 27629 20284
rect 27663 20281 27675 20315
rect 27617 20275 27675 20281
rect 28994 20272 29000 20324
rect 29052 20312 29058 20324
rect 29089 20315 29147 20321
rect 29089 20312 29101 20315
rect 29052 20284 29101 20312
rect 29052 20272 29058 20284
rect 29089 20281 29101 20284
rect 29135 20312 29147 20315
rect 29273 20315 29331 20321
rect 29273 20312 29285 20315
rect 29135 20284 29285 20312
rect 29135 20281 29147 20284
rect 29089 20275 29147 20281
rect 29273 20281 29285 20284
rect 29319 20312 29331 20315
rect 29748 20312 29776 20352
rect 32769 20349 32781 20383
rect 32815 20380 32827 20383
rect 33226 20380 33232 20392
rect 32815 20352 33232 20380
rect 32815 20349 32827 20352
rect 32769 20343 32827 20349
rect 33226 20340 33232 20352
rect 33284 20340 33290 20392
rect 33410 20340 33416 20392
rect 33468 20380 33474 20392
rect 36449 20383 36507 20389
rect 36449 20380 36461 20383
rect 33468 20352 36461 20380
rect 33468 20340 33474 20352
rect 36449 20349 36461 20352
rect 36495 20380 36507 20383
rect 36630 20380 36636 20392
rect 36495 20352 36636 20380
rect 36495 20349 36507 20352
rect 36449 20343 36507 20349
rect 36630 20340 36636 20352
rect 36688 20340 36694 20392
rect 36814 20340 36820 20392
rect 36872 20380 36878 20392
rect 37093 20383 37151 20389
rect 37093 20380 37105 20383
rect 36872 20352 37105 20380
rect 36872 20340 36878 20352
rect 37093 20349 37105 20352
rect 37139 20349 37151 20383
rect 38838 20380 38844 20392
rect 38799 20352 38844 20380
rect 37093 20343 37151 20349
rect 38838 20340 38844 20352
rect 38896 20340 38902 20392
rect 38930 20340 38936 20392
rect 38988 20380 38994 20392
rect 39301 20383 39359 20389
rect 39301 20380 39313 20383
rect 38988 20352 39313 20380
rect 38988 20340 38994 20352
rect 39301 20349 39313 20352
rect 39347 20349 39359 20383
rect 39301 20343 39359 20349
rect 39577 20383 39635 20389
rect 39577 20349 39589 20383
rect 39623 20380 39635 20383
rect 40494 20380 40500 20392
rect 39623 20352 40500 20380
rect 39623 20349 39635 20352
rect 39577 20343 39635 20349
rect 40494 20340 40500 20352
rect 40552 20340 40558 20392
rect 29319 20284 29776 20312
rect 29825 20315 29883 20321
rect 29319 20281 29331 20284
rect 29273 20275 29331 20281
rect 29825 20281 29837 20315
rect 29871 20312 29883 20315
rect 30190 20312 30196 20324
rect 29871 20284 30196 20312
rect 29871 20281 29883 20284
rect 29825 20275 29883 20281
rect 30190 20272 30196 20284
rect 30248 20272 30254 20324
rect 30742 20272 30748 20324
rect 30800 20312 30806 20324
rect 31342 20315 31400 20321
rect 31342 20312 31354 20315
rect 30800 20284 31354 20312
rect 30800 20272 30806 20284
rect 31342 20281 31354 20284
rect 31388 20281 31400 20315
rect 31342 20275 31400 20281
rect 34514 20272 34520 20324
rect 34572 20312 34578 20324
rect 35206 20315 35264 20321
rect 35206 20312 35218 20315
rect 34572 20284 35218 20312
rect 34572 20272 34578 20284
rect 35206 20281 35218 20284
rect 35252 20281 35264 20315
rect 40310 20312 40316 20324
rect 40223 20284 40316 20312
rect 35206 20275 35264 20281
rect 21600 20216 22324 20244
rect 21600 20204 21606 20216
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 23799 20247 23857 20253
rect 23799 20244 23811 20247
rect 22428 20216 23811 20244
rect 22428 20204 22434 20216
rect 23799 20213 23811 20216
rect 23845 20213 23857 20247
rect 23799 20207 23857 20213
rect 25038 20204 25044 20256
rect 25096 20244 25102 20256
rect 25179 20247 25237 20253
rect 25179 20244 25191 20247
rect 25096 20216 25191 20244
rect 25096 20204 25102 20216
rect 25179 20213 25191 20216
rect 25225 20213 25237 20247
rect 30098 20244 30104 20256
rect 30059 20216 30104 20244
rect 25179 20207 25237 20213
rect 30098 20204 30104 20216
rect 30156 20204 30162 20256
rect 34146 20244 34152 20256
rect 34107 20216 34152 20244
rect 34146 20204 34152 20216
rect 34204 20204 34210 20256
rect 35802 20244 35808 20256
rect 35763 20216 35808 20244
rect 35802 20204 35808 20216
rect 35860 20204 35866 20256
rect 36722 20244 36728 20256
rect 36683 20216 36728 20244
rect 36722 20204 36728 20216
rect 36780 20204 36786 20256
rect 38010 20204 38016 20256
rect 38068 20244 38074 20256
rect 40236 20253 40264 20284
rect 40310 20272 40316 20284
rect 40368 20312 40374 20324
rect 40833 20321 40861 20488
rect 43990 20476 43996 20488
rect 44048 20476 44054 20528
rect 45281 20519 45339 20525
rect 45281 20485 45293 20519
rect 45327 20516 45339 20519
rect 45370 20516 45376 20528
rect 45327 20488 45376 20516
rect 45327 20485 45339 20488
rect 45281 20479 45339 20485
rect 45370 20476 45376 20488
rect 45428 20516 45434 20528
rect 45557 20519 45615 20525
rect 45557 20516 45569 20519
rect 45428 20488 45569 20516
rect 45428 20476 45434 20488
rect 45557 20485 45569 20488
rect 45603 20516 45615 20519
rect 47026 20516 47032 20528
rect 45603 20488 47032 20516
rect 45603 20485 45615 20488
rect 45557 20479 45615 20485
rect 47026 20476 47032 20488
rect 47084 20476 47090 20528
rect 43162 20408 43168 20460
rect 43220 20448 43226 20460
rect 43717 20451 43775 20457
rect 43717 20448 43729 20451
rect 43220 20420 43729 20448
rect 43220 20408 43226 20420
rect 43717 20417 43729 20420
rect 43763 20448 43775 20451
rect 43763 20420 46888 20448
rect 43763 20417 43775 20420
rect 43717 20411 43775 20417
rect 45056 20383 45114 20389
rect 45056 20349 45068 20383
rect 45102 20380 45114 20383
rect 45281 20383 45339 20389
rect 45281 20380 45293 20383
rect 45102 20352 45293 20380
rect 45102 20349 45114 20352
rect 45056 20343 45114 20349
rect 45281 20349 45293 20352
rect 45327 20349 45339 20383
rect 45281 20343 45339 20349
rect 46860 20324 46888 20420
rect 40818 20315 40876 20321
rect 40818 20312 40830 20315
rect 40368 20284 40830 20312
rect 40368 20272 40374 20284
rect 40818 20281 40830 20284
rect 40864 20281 40876 20315
rect 40818 20275 40876 20281
rect 41322 20272 41328 20324
rect 41380 20312 41386 20324
rect 42061 20315 42119 20321
rect 42061 20312 42073 20315
rect 41380 20284 42073 20312
rect 41380 20272 41386 20284
rect 42061 20281 42073 20284
rect 42107 20281 42119 20315
rect 43070 20312 43076 20324
rect 43031 20284 43076 20312
rect 42061 20275 42119 20281
rect 43070 20272 43076 20284
rect 43128 20272 43134 20324
rect 43165 20315 43223 20321
rect 43165 20281 43177 20315
rect 43211 20281 43223 20315
rect 43165 20275 43223 20281
rect 45143 20315 45201 20321
rect 45143 20281 45155 20315
rect 45189 20312 45201 20315
rect 46198 20312 46204 20324
rect 45189 20284 46204 20312
rect 45189 20281 45201 20284
rect 45143 20275 45201 20281
rect 40221 20247 40279 20253
rect 40221 20244 40233 20247
rect 38068 20216 40233 20244
rect 38068 20204 38074 20216
rect 40221 20213 40233 20216
rect 40267 20213 40279 20247
rect 41414 20244 41420 20256
rect 41327 20216 41420 20244
rect 40221 20207 40279 20213
rect 41414 20204 41420 20216
rect 41472 20244 41478 20256
rect 41785 20247 41843 20253
rect 41785 20244 41797 20247
rect 41472 20216 41797 20244
rect 41472 20204 41478 20216
rect 41785 20213 41797 20216
rect 41831 20244 41843 20247
rect 41874 20244 41880 20256
rect 41831 20216 41880 20244
rect 41831 20213 41843 20216
rect 41785 20207 41843 20213
rect 41874 20204 41880 20216
rect 41932 20204 41938 20256
rect 42886 20204 42892 20256
rect 42944 20244 42950 20256
rect 43180 20244 43208 20275
rect 46198 20272 46204 20284
rect 46256 20272 46262 20324
rect 46293 20315 46351 20321
rect 46293 20281 46305 20315
rect 46339 20281 46351 20315
rect 46842 20312 46848 20324
rect 46803 20284 46848 20312
rect 46293 20275 46351 20281
rect 42944 20216 43208 20244
rect 42944 20204 42950 20216
rect 45738 20204 45744 20256
rect 45796 20244 45802 20256
rect 46308 20244 46336 20275
rect 46842 20272 46848 20284
rect 46900 20272 46906 20324
rect 45796 20216 46336 20244
rect 45796 20204 45802 20216
rect 1104 20154 48852 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 48852 20154
rect 1104 20080 48852 20102
rect 18046 20040 18052 20052
rect 18007 20012 18052 20040
rect 18046 20000 18052 20012
rect 18104 20040 18110 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18104 20012 18797 20040
rect 18104 20000 18110 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 18785 20003 18843 20009
rect 18943 20012 19533 20040
rect 18601 19975 18659 19981
rect 18601 19972 18613 19975
rect 16822 19944 18613 19972
rect 16822 19916 16850 19944
rect 18601 19941 18613 19944
rect 18647 19941 18659 19975
rect 18601 19935 18659 19941
rect 16822 19913 16856 19916
rect 16807 19907 16856 19913
rect 16807 19904 16819 19907
rect 16763 19876 16819 19904
rect 16807 19873 16819 19876
rect 16853 19873 16856 19907
rect 16807 19867 16856 19873
rect 16850 19864 16856 19867
rect 16908 19864 16914 19916
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17773 19907 17831 19913
rect 17773 19904 17785 19907
rect 17552 19876 17785 19904
rect 17552 19864 17558 19876
rect 17773 19873 17785 19876
rect 17819 19904 17831 19907
rect 18230 19904 18236 19916
rect 17819 19876 18236 19904
rect 17819 19873 17831 19876
rect 17773 19867 17831 19873
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18506 19904 18512 19916
rect 18371 19876 18512 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 18340 19836 18368 19867
rect 18506 19864 18512 19876
rect 18564 19904 18570 19916
rect 18943 19904 18971 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 21266 20040 21272 20052
rect 21227 20012 21272 20040
rect 19521 20003 19579 20009
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21818 20040 21824 20052
rect 21779 20012 21824 20040
rect 21818 20000 21824 20012
rect 21876 20000 21882 20052
rect 26145 20043 26203 20049
rect 26145 20009 26157 20043
rect 26191 20040 26203 20043
rect 26510 20040 26516 20052
rect 26191 20012 26516 20040
rect 26191 20009 26203 20012
rect 26145 20003 26203 20009
rect 26510 20000 26516 20012
rect 26568 20000 26574 20052
rect 27706 20040 27712 20052
rect 27667 20012 27712 20040
rect 27706 20000 27712 20012
rect 27764 20000 27770 20052
rect 29822 20040 29828 20052
rect 29783 20012 29828 20040
rect 29822 20000 29828 20012
rect 29880 20000 29886 20052
rect 32309 20043 32367 20049
rect 32309 20009 32321 20043
rect 32355 20040 32367 20043
rect 32398 20040 32404 20052
rect 32355 20012 32404 20040
rect 32355 20009 32367 20012
rect 32309 20003 32367 20009
rect 32398 20000 32404 20012
rect 32456 20000 32462 20052
rect 33321 20043 33379 20049
rect 33321 20009 33333 20043
rect 33367 20040 33379 20043
rect 33778 20040 33784 20052
rect 33367 20012 33784 20040
rect 33367 20009 33379 20012
rect 33321 20003 33379 20009
rect 33778 20000 33784 20012
rect 33836 20000 33842 20052
rect 34514 20000 34520 20052
rect 34572 20040 34578 20052
rect 34885 20043 34943 20049
rect 34885 20040 34897 20043
rect 34572 20012 34897 20040
rect 34572 20000 34578 20012
rect 34885 20009 34897 20012
rect 34931 20009 34943 20043
rect 34885 20003 34943 20009
rect 35802 20000 35808 20052
rect 35860 20040 35866 20052
rect 36081 20043 36139 20049
rect 36081 20040 36093 20043
rect 35860 20012 36093 20040
rect 35860 20000 35866 20012
rect 36081 20009 36093 20012
rect 36127 20009 36139 20043
rect 36081 20003 36139 20009
rect 36354 20000 36360 20052
rect 36412 20040 36418 20052
rect 36449 20043 36507 20049
rect 36449 20040 36461 20043
rect 36412 20012 36461 20040
rect 36412 20000 36418 20012
rect 36449 20009 36461 20012
rect 36495 20009 36507 20043
rect 36449 20003 36507 20009
rect 36771 20043 36829 20049
rect 36771 20009 36783 20043
rect 36817 20040 36829 20043
rect 37458 20040 37464 20052
rect 36817 20012 37464 20040
rect 36817 20009 36829 20012
rect 36771 20003 36829 20009
rect 37458 20000 37464 20012
rect 37516 20000 37522 20052
rect 38473 20043 38531 20049
rect 38473 20009 38485 20043
rect 38519 20040 38531 20043
rect 38930 20040 38936 20052
rect 38519 20012 38936 20040
rect 38519 20009 38531 20012
rect 38473 20003 38531 20009
rect 38930 20000 38936 20012
rect 38988 20000 38994 20052
rect 40494 20040 40500 20052
rect 40455 20012 40500 20040
rect 40494 20000 40500 20012
rect 40552 20000 40558 20052
rect 43070 20040 43076 20052
rect 42983 20012 43076 20040
rect 43070 20000 43076 20012
rect 43128 20040 43134 20052
rect 45051 20043 45109 20049
rect 45051 20040 45063 20043
rect 43128 20012 45063 20040
rect 43128 20000 43134 20012
rect 45051 20009 45063 20012
rect 45097 20009 45109 20043
rect 45738 20040 45744 20052
rect 45699 20012 45744 20040
rect 45051 20003 45109 20009
rect 45738 20000 45744 20012
rect 45796 20000 45802 20052
rect 46198 20000 46204 20052
rect 46256 20040 46262 20052
rect 46385 20043 46443 20049
rect 46385 20040 46397 20043
rect 46256 20012 46397 20040
rect 46256 20000 46262 20012
rect 46385 20009 46397 20012
rect 46431 20009 46443 20043
rect 46385 20003 46443 20009
rect 23290 19972 23296 19984
rect 23251 19944 23296 19972
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 26697 19975 26755 19981
rect 26697 19941 26709 19975
rect 26743 19972 26755 19975
rect 27246 19972 27252 19984
rect 26743 19944 27252 19972
rect 26743 19941 26755 19944
rect 26697 19935 26755 19941
rect 27246 19932 27252 19944
rect 27304 19932 27310 19984
rect 28994 19972 29000 19984
rect 28955 19944 29000 19972
rect 28994 19932 29000 19944
rect 29052 19932 29058 19984
rect 32674 19972 32680 19984
rect 30944 19944 32680 19972
rect 30944 19916 30972 19944
rect 32674 19932 32680 19944
rect 32732 19932 32738 19984
rect 33870 19972 33876 19984
rect 33152 19944 33876 19972
rect 19334 19904 19340 19916
rect 18564 19876 18971 19904
rect 19295 19876 19340 19904
rect 18564 19864 18570 19876
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 22370 19904 22376 19916
rect 19904 19876 22376 19904
rect 17727 19808 18368 19836
rect 18601 19839 18659 19845
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 19904 19836 19932 19876
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 24946 19904 24952 19916
rect 24907 19876 24952 19904
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 29181 19907 29239 19913
rect 29181 19873 29193 19907
rect 29227 19904 29239 19907
rect 29270 19904 29276 19916
rect 29227 19876 29276 19904
rect 29227 19873 29239 19876
rect 29181 19867 29239 19873
rect 29270 19864 29276 19876
rect 29328 19864 29334 19916
rect 30745 19907 30803 19913
rect 30745 19873 30757 19907
rect 30791 19904 30803 19907
rect 30834 19904 30840 19916
rect 30791 19876 30840 19904
rect 30791 19873 30803 19876
rect 30745 19867 30803 19873
rect 30834 19864 30840 19876
rect 30892 19864 30898 19916
rect 30926 19864 30932 19916
rect 30984 19904 30990 19916
rect 30984 19876 31077 19904
rect 30984 19864 30990 19876
rect 31938 19864 31944 19916
rect 31996 19904 32002 19916
rect 33152 19913 33180 19944
rect 33870 19932 33876 19944
rect 33928 19932 33934 19984
rect 38948 19972 38976 20000
rect 38948 19944 39804 19972
rect 32125 19907 32183 19913
rect 32125 19904 32137 19907
rect 31996 19876 32137 19904
rect 31996 19864 32002 19876
rect 32125 19873 32137 19876
rect 32171 19873 32183 19907
rect 32125 19867 32183 19873
rect 33137 19907 33195 19913
rect 33137 19873 33149 19907
rect 33183 19873 33195 19907
rect 34425 19907 34483 19913
rect 34425 19904 34437 19907
rect 33137 19867 33195 19873
rect 33244 19876 34437 19904
rect 20898 19836 20904 19848
rect 18647 19808 19932 19836
rect 20859 19808 20904 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 23201 19839 23259 19845
rect 23201 19836 23213 19839
rect 22940 19808 23213 19836
rect 22940 19777 22968 19808
rect 23201 19805 23213 19808
rect 23247 19805 23259 19839
rect 23474 19836 23480 19848
rect 23435 19808 23480 19836
rect 23201 19799 23259 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 25590 19836 25596 19848
rect 25551 19808 25596 19836
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 26605 19839 26663 19845
rect 26605 19805 26617 19839
rect 26651 19805 26663 19839
rect 26878 19836 26884 19848
rect 26839 19808 26884 19836
rect 26605 19799 26663 19805
rect 16899 19771 16957 19777
rect 16899 19737 16911 19771
rect 16945 19768 16957 19771
rect 22925 19771 22983 19777
rect 22925 19768 22937 19771
rect 16945 19740 22937 19768
rect 16945 19737 16957 19740
rect 16899 19731 16957 19737
rect 22925 19737 22937 19740
rect 22971 19737 22983 19771
rect 22925 19731 22983 19737
rect 25682 19728 25688 19780
rect 25740 19768 25746 19780
rect 26620 19768 26648 19799
rect 26878 19796 26884 19808
rect 26936 19796 26942 19848
rect 31018 19836 31024 19848
rect 30979 19808 31024 19836
rect 31018 19796 31024 19808
rect 31076 19796 31082 19848
rect 32950 19796 32956 19848
rect 33008 19836 33014 19848
rect 33244 19836 33272 19876
rect 34425 19873 34437 19876
rect 34471 19873 34483 19907
rect 35618 19904 35624 19916
rect 35579 19876 35624 19904
rect 34425 19867 34483 19873
rect 35618 19864 35624 19876
rect 35676 19864 35682 19916
rect 36170 19864 36176 19916
rect 36228 19904 36234 19916
rect 36668 19907 36726 19913
rect 36668 19904 36680 19907
rect 36228 19876 36680 19904
rect 36228 19864 36234 19876
rect 36668 19873 36680 19876
rect 36714 19873 36726 19907
rect 36668 19867 36726 19873
rect 38298 19907 38356 19913
rect 38298 19873 38310 19907
rect 38344 19873 38356 19907
rect 39298 19904 39304 19916
rect 39259 19876 39304 19904
rect 38298 19867 38356 19873
rect 33008 19808 33272 19836
rect 33008 19796 33014 19808
rect 27614 19768 27620 19780
rect 25740 19740 27620 19768
rect 25740 19728 25746 19740
rect 27614 19728 27620 19740
rect 27672 19728 27678 19780
rect 27706 19728 27712 19780
rect 27764 19768 27770 19780
rect 31110 19768 31116 19780
rect 27764 19740 31116 19768
rect 27764 19728 27770 19740
rect 31110 19728 31116 19740
rect 31168 19728 31174 19780
rect 35805 19771 35863 19777
rect 35805 19737 35817 19771
rect 35851 19768 35863 19771
rect 38304 19768 38332 19867
rect 39298 19864 39304 19876
rect 39356 19864 39362 19916
rect 39776 19913 39804 19944
rect 41598 19932 41604 19984
rect 41656 19972 41662 19984
rect 41785 19975 41843 19981
rect 41785 19972 41797 19975
rect 41656 19944 41797 19972
rect 41656 19932 41662 19944
rect 41785 19941 41797 19944
rect 41831 19941 41843 19975
rect 41785 19935 41843 19941
rect 41874 19932 41880 19984
rect 41932 19972 41938 19984
rect 42429 19975 42487 19981
rect 41932 19944 41977 19972
rect 41932 19932 41938 19944
rect 42429 19941 42441 19975
rect 42475 19972 42487 19975
rect 43533 19975 43591 19981
rect 42475 19944 42794 19972
rect 42475 19941 42487 19944
rect 42429 19935 42487 19941
rect 39761 19907 39819 19913
rect 39761 19873 39773 19907
rect 39807 19873 39819 19907
rect 39761 19867 39819 19873
rect 40034 19836 40040 19848
rect 39995 19808 40040 19836
rect 40034 19796 40040 19808
rect 40092 19796 40098 19848
rect 42766 19836 42794 19944
rect 43533 19941 43545 19975
rect 43579 19972 43591 19975
rect 43714 19972 43720 19984
rect 43579 19944 43720 19972
rect 43579 19941 43591 19944
rect 43533 19935 43591 19941
rect 43714 19932 43720 19944
rect 43772 19932 43778 19984
rect 44818 19864 44824 19916
rect 44876 19904 44882 19916
rect 44948 19907 45006 19913
rect 44948 19904 44960 19907
rect 44876 19876 44960 19904
rect 44876 19864 44882 19876
rect 44948 19873 44960 19876
rect 44994 19873 45006 19907
rect 45830 19904 45836 19916
rect 45791 19876 45836 19904
rect 44948 19867 45006 19873
rect 45830 19864 45836 19876
rect 45888 19864 45894 19916
rect 43438 19836 43444 19848
rect 42766 19808 43444 19836
rect 43438 19796 43444 19808
rect 43496 19796 43502 19848
rect 43622 19796 43628 19848
rect 43680 19836 43686 19848
rect 43717 19839 43775 19845
rect 43717 19836 43729 19839
rect 43680 19808 43729 19836
rect 43680 19796 43686 19808
rect 43717 19805 43729 19808
rect 43763 19805 43775 19839
rect 43717 19799 43775 19805
rect 38378 19768 38384 19780
rect 35851 19740 38384 19768
rect 35851 19737 35863 19740
rect 35805 19731 35863 19737
rect 38378 19728 38384 19740
rect 38436 19768 38442 19780
rect 39117 19771 39175 19777
rect 39117 19768 39129 19771
rect 38436 19740 39129 19768
rect 38436 19728 38442 19740
rect 39117 19737 39129 19740
rect 39163 19737 39175 19771
rect 39117 19731 39175 19737
rect 45278 19728 45284 19780
rect 45336 19768 45342 19780
rect 46063 19771 46121 19777
rect 46063 19768 46075 19771
rect 45336 19740 46075 19768
rect 45336 19728 45342 19740
rect 46063 19737 46075 19740
rect 46109 19737 46121 19771
rect 46063 19731 46121 19737
rect 20070 19700 20076 19712
rect 20031 19672 20076 19700
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 25406 19660 25412 19712
rect 25464 19700 25470 19712
rect 29273 19703 29331 19709
rect 29273 19700 29285 19703
rect 25464 19672 29285 19700
rect 25464 19660 25470 19672
rect 29273 19669 29285 19672
rect 29319 19669 29331 19703
rect 34606 19700 34612 19712
rect 34567 19672 34612 19700
rect 29273 19663 29331 19669
rect 34606 19660 34612 19672
rect 34664 19660 34670 19712
rect 35250 19700 35256 19712
rect 35211 19672 35256 19700
rect 35250 19660 35256 19672
rect 35308 19660 35314 19712
rect 41414 19700 41420 19712
rect 41375 19672 41420 19700
rect 41414 19660 41420 19672
rect 41472 19660 41478 19712
rect 1104 19610 48852 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 48852 19610
rect 1104 19536 48852 19558
rect 19334 19496 19340 19508
rect 19295 19468 19340 19496
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 20898 19456 20904 19508
rect 20956 19496 20962 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 20956 19468 22017 19496
rect 20956 19456 20962 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22281 19499 22339 19505
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 23382 19496 23388 19508
rect 22327 19468 23388 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 23382 19456 23388 19468
rect 23440 19456 23446 19508
rect 24946 19496 24952 19508
rect 24907 19468 24952 19496
rect 24946 19456 24952 19468
rect 25004 19456 25010 19508
rect 25682 19496 25688 19508
rect 25643 19468 25688 19496
rect 25682 19456 25688 19468
rect 25740 19456 25746 19508
rect 26050 19496 26056 19508
rect 26011 19468 26056 19496
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 27246 19496 27252 19508
rect 27207 19468 27252 19496
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 30561 19499 30619 19505
rect 30561 19465 30573 19499
rect 30607 19496 30619 19499
rect 30834 19496 30840 19508
rect 30607 19468 30840 19496
rect 30607 19465 30619 19468
rect 30561 19459 30619 19465
rect 30834 19456 30840 19468
rect 30892 19456 30898 19508
rect 30926 19456 30932 19508
rect 30984 19496 30990 19508
rect 30984 19468 31029 19496
rect 30984 19456 30990 19468
rect 31110 19456 31116 19508
rect 31168 19496 31174 19508
rect 33502 19496 33508 19508
rect 31168 19468 33508 19496
rect 31168 19456 31174 19468
rect 33502 19456 33508 19468
rect 33560 19456 33566 19508
rect 35618 19456 35624 19508
rect 35676 19496 35682 19508
rect 36081 19499 36139 19505
rect 36081 19496 36093 19499
rect 35676 19468 36093 19496
rect 35676 19456 35682 19468
rect 36081 19465 36093 19468
rect 36127 19465 36139 19499
rect 38378 19496 38384 19508
rect 38339 19468 38384 19496
rect 36081 19459 36139 19465
rect 38378 19456 38384 19468
rect 38436 19456 38442 19508
rect 38930 19496 38936 19508
rect 38891 19468 38936 19496
rect 38930 19456 38936 19468
rect 38988 19456 38994 19508
rect 39531 19499 39589 19505
rect 39531 19465 39543 19499
rect 39577 19496 39589 19499
rect 41322 19496 41328 19508
rect 39577 19468 41328 19496
rect 39577 19465 39589 19468
rect 39531 19459 39589 19465
rect 41322 19456 41328 19468
rect 41380 19456 41386 19508
rect 41874 19456 41880 19508
rect 41932 19496 41938 19508
rect 42337 19499 42395 19505
rect 42337 19496 42349 19499
rect 41932 19468 42349 19496
rect 41932 19456 41938 19468
rect 42337 19465 42349 19468
rect 42383 19465 42395 19499
rect 42337 19459 42395 19465
rect 44818 19456 44824 19508
rect 44876 19496 44882 19508
rect 45465 19499 45523 19505
rect 45465 19496 45477 19499
rect 44876 19468 45477 19496
rect 44876 19456 44882 19468
rect 45465 19465 45477 19468
rect 45511 19465 45523 19499
rect 45465 19459 45523 19465
rect 45830 19456 45836 19508
rect 45888 19496 45894 19508
rect 46293 19499 46351 19505
rect 46293 19496 46305 19499
rect 45888 19468 46305 19496
rect 45888 19456 45894 19468
rect 46293 19465 46305 19468
rect 46339 19465 46351 19499
rect 46293 19459 46351 19465
rect 16301 19431 16359 19437
rect 16301 19397 16313 19431
rect 16347 19428 16359 19431
rect 18046 19428 18052 19440
rect 16347 19400 18052 19428
rect 16347 19397 16359 19400
rect 16301 19391 16359 19397
rect 16408 19301 16436 19400
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 19352 19428 19380 19456
rect 25406 19428 25412 19440
rect 19352 19400 25412 19428
rect 25406 19388 25412 19400
rect 25464 19388 25470 19440
rect 26789 19431 26847 19437
rect 26789 19397 26801 19431
rect 26835 19428 26847 19431
rect 26878 19428 26884 19440
rect 26835 19400 26884 19428
rect 26835 19397 26847 19400
rect 26789 19391 26847 19397
rect 26878 19388 26884 19400
rect 26936 19388 26942 19440
rect 30852 19428 30880 19456
rect 36446 19428 36452 19440
rect 30852 19400 36452 19428
rect 36446 19388 36452 19400
rect 36504 19388 36510 19440
rect 36630 19388 36636 19440
rect 36688 19428 36694 19440
rect 39209 19431 39267 19437
rect 39209 19428 39221 19431
rect 36688 19400 39221 19428
rect 36688 19388 36694 19400
rect 39209 19397 39221 19400
rect 39255 19428 39267 19431
rect 39298 19428 39304 19440
rect 39255 19400 39304 19428
rect 39255 19397 39267 19400
rect 39209 19391 39267 19397
rect 39298 19388 39304 19400
rect 39356 19388 39362 19440
rect 20254 19360 20260 19372
rect 16960 19332 18552 19360
rect 20167 19332 20260 19360
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19261 16451 19295
rect 16393 19255 16451 19261
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 16960 19301 16988 19332
rect 18524 19304 18552 19332
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19360 20499 19363
rect 20714 19360 20720 19372
rect 20487 19332 20720 19360
rect 20487 19329 20499 19332
rect 20441 19323 20499 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 22646 19360 22652 19372
rect 21238 19332 22652 19360
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16540 19264 16957 19292
rect 16540 19252 16546 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19261 18383 19295
rect 18506 19292 18512 19304
rect 18467 19264 18512 19292
rect 18325 19255 18383 19261
rect 17126 19224 17132 19236
rect 17087 19196 17132 19224
rect 17126 19184 17132 19196
rect 17184 19184 17190 19236
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 18340 19224 18368 19255
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 19242 19292 19248 19304
rect 18616 19264 19248 19292
rect 18616 19224 18644 19264
rect 19242 19252 19248 19264
rect 19300 19292 19306 19304
rect 21238 19292 21266 19332
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 23750 19320 23756 19372
rect 23808 19360 23814 19372
rect 28261 19363 28319 19369
rect 28261 19360 28273 19363
rect 23808 19332 28273 19360
rect 23808 19320 23814 19332
rect 28261 19329 28273 19332
rect 28307 19329 28319 19363
rect 28261 19323 28319 19329
rect 34698 19320 34704 19372
rect 34756 19360 34762 19372
rect 34885 19363 34943 19369
rect 34885 19360 34897 19363
rect 34756 19332 34897 19360
rect 34756 19320 34762 19332
rect 34885 19329 34897 19332
rect 34931 19360 34943 19363
rect 35250 19360 35256 19372
rect 34931 19332 35256 19360
rect 34931 19329 34943 19332
rect 34885 19323 34943 19329
rect 35250 19320 35256 19332
rect 35308 19320 35314 19372
rect 37461 19363 37519 19369
rect 37461 19329 37473 19363
rect 37507 19360 37519 19363
rect 37642 19360 37648 19372
rect 37507 19332 37648 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 37642 19320 37648 19332
rect 37700 19320 37706 19372
rect 37918 19320 37924 19372
rect 37976 19360 37982 19372
rect 39853 19363 39911 19369
rect 39853 19360 39865 19363
rect 37976 19332 39865 19360
rect 37976 19320 37982 19332
rect 19300 19264 21266 19292
rect 22557 19295 22615 19301
rect 19300 19252 19306 19264
rect 22557 19261 22569 19295
rect 22603 19292 22615 19295
rect 23106 19292 23112 19304
rect 22603 19264 23112 19292
rect 22603 19261 22615 19264
rect 22557 19255 22615 19261
rect 23106 19252 23112 19264
rect 23164 19252 23170 19304
rect 23658 19292 23664 19304
rect 23619 19264 23664 19292
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 24019 19264 24593 19292
rect 17911 19196 18644 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 20254 19184 20260 19236
rect 20312 19224 20318 19236
rect 20622 19224 20628 19236
rect 20312 19196 20628 19224
rect 20312 19184 20318 19196
rect 20622 19184 20628 19196
rect 20680 19224 20686 19236
rect 20803 19227 20861 19233
rect 20803 19224 20815 19227
rect 20680 19196 20815 19224
rect 20680 19184 20686 19196
rect 20803 19193 20815 19196
rect 20849 19224 20861 19227
rect 21266 19224 21272 19236
rect 20849 19196 21272 19224
rect 20849 19193 20861 19196
rect 20803 19187 20861 19193
rect 21266 19184 21272 19196
rect 21324 19224 21330 19236
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 21324 19196 21649 19224
rect 21324 19184 21330 19196
rect 21637 19193 21649 19196
rect 21683 19224 21695 19227
rect 22281 19227 22339 19233
rect 22281 19224 22293 19227
rect 21683 19196 22293 19224
rect 21683 19193 21695 19196
rect 21637 19187 21695 19193
rect 22281 19193 22293 19196
rect 22327 19193 22339 19227
rect 22281 19187 22339 19193
rect 22465 19227 22523 19233
rect 22465 19193 22477 19227
rect 22511 19224 22523 19227
rect 23290 19224 23296 19236
rect 22511 19196 23296 19224
rect 22511 19193 22523 19196
rect 22465 19187 22523 19193
rect 23290 19184 23296 19196
rect 23348 19224 23354 19236
rect 24019 19224 24047 19264
rect 24581 19261 24593 19264
rect 24627 19261 24639 19295
rect 24581 19255 24639 19261
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19292 27767 19295
rect 27985 19295 28043 19301
rect 27985 19292 27997 19295
rect 27755 19264 27997 19292
rect 27755 19261 27767 19264
rect 27709 19255 27767 19261
rect 27985 19261 27997 19264
rect 28031 19292 28043 19295
rect 28629 19295 28687 19301
rect 28629 19292 28641 19295
rect 28031 19264 28641 19292
rect 28031 19261 28043 19264
rect 27985 19255 28043 19261
rect 28629 19261 28641 19264
rect 28675 19292 28687 19295
rect 29270 19292 29276 19304
rect 28675 19264 29276 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 29270 19252 29276 19264
rect 29328 19252 29334 19304
rect 29917 19295 29975 19301
rect 29917 19261 29929 19295
rect 29963 19292 29975 19295
rect 30098 19292 30104 19304
rect 29963 19264 30104 19292
rect 29963 19261 29975 19264
rect 29917 19255 29975 19261
rect 26234 19224 26240 19236
rect 23348 19196 24047 19224
rect 26195 19196 26240 19224
rect 23348 19184 23354 19196
rect 26234 19184 26240 19196
rect 26292 19184 26298 19236
rect 26329 19227 26387 19233
rect 26329 19193 26341 19227
rect 26375 19193 26387 19227
rect 27798 19224 27804 19236
rect 27759 19196 27804 19224
rect 26329 19187 26387 19193
rect 17494 19156 17500 19168
rect 17455 19128 17500 19156
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18138 19156 18144 19168
rect 18099 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 21358 19156 21364 19168
rect 21319 19128 21364 19156
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 22738 19156 22744 19168
rect 22699 19128 22744 19156
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 23106 19156 23112 19168
rect 23067 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 23934 19116 23940 19168
rect 23992 19156 23998 19168
rect 24029 19159 24087 19165
rect 24029 19156 24041 19159
rect 23992 19128 24041 19156
rect 23992 19116 23998 19128
rect 24029 19125 24041 19128
rect 24075 19125 24087 19159
rect 24029 19119 24087 19125
rect 26050 19116 26056 19168
rect 26108 19156 26114 19168
rect 26344 19156 26372 19187
rect 27798 19184 27804 19196
rect 27856 19184 27862 19236
rect 29089 19227 29147 19233
rect 29089 19193 29101 19227
rect 29135 19224 29147 19227
rect 29932 19224 29960 19255
rect 30098 19252 30104 19264
rect 30156 19292 30162 19304
rect 30742 19292 30748 19304
rect 30156 19264 30748 19292
rect 30156 19252 30162 19264
rect 30742 19252 30748 19264
rect 30800 19252 30806 19304
rect 31849 19295 31907 19301
rect 31849 19261 31861 19295
rect 31895 19292 31907 19295
rect 32398 19292 32404 19304
rect 31895 19264 32404 19292
rect 31895 19261 31907 19264
rect 31849 19255 31907 19261
rect 32398 19252 32404 19264
rect 32456 19252 32462 19304
rect 33045 19295 33103 19301
rect 33045 19261 33057 19295
rect 33091 19292 33103 19295
rect 33091 19264 33640 19292
rect 33091 19261 33103 19264
rect 33045 19255 33103 19261
rect 31665 19227 31723 19233
rect 31665 19224 31677 19227
rect 29135 19196 29960 19224
rect 31496 19196 31677 19224
rect 29135 19193 29147 19196
rect 29089 19187 29147 19193
rect 31496 19168 31524 19196
rect 31665 19193 31677 19196
rect 31711 19193 31723 19227
rect 32861 19227 32919 19233
rect 32861 19224 32873 19227
rect 31665 19187 31723 19193
rect 31956 19196 32873 19224
rect 31956 19168 31984 19196
rect 32861 19193 32873 19196
rect 32907 19193 32919 19227
rect 32861 19187 32919 19193
rect 33612 19168 33640 19264
rect 34514 19252 34520 19304
rect 34572 19292 34578 19304
rect 34572 19264 35249 19292
rect 34572 19252 34578 19264
rect 35221 19233 35249 19264
rect 36170 19252 36176 19304
rect 36228 19292 36234 19304
rect 39443 19301 39471 19332
rect 39853 19329 39865 19332
rect 39899 19329 39911 19363
rect 43254 19360 43260 19372
rect 39853 19323 39911 19329
rect 42766 19332 43260 19360
rect 36633 19295 36691 19301
rect 36633 19292 36645 19295
rect 36228 19264 36645 19292
rect 36228 19252 36234 19264
rect 36633 19261 36645 19264
rect 36679 19261 36691 19295
rect 36633 19255 36691 19261
rect 39428 19295 39486 19301
rect 39428 19261 39440 19295
rect 39474 19261 39486 19295
rect 39428 19255 39486 19261
rect 35206 19227 35264 19233
rect 35206 19193 35218 19227
rect 35252 19193 35264 19227
rect 36648 19224 36676 19255
rect 37458 19224 37464 19236
rect 36648 19196 37464 19224
rect 35206 19187 35264 19193
rect 37458 19184 37464 19196
rect 37516 19184 37522 19236
rect 37550 19184 37556 19236
rect 37608 19224 37614 19236
rect 38105 19227 38163 19233
rect 37608 19196 37653 19224
rect 37608 19184 37614 19196
rect 38105 19193 38117 19227
rect 38151 19224 38163 19227
rect 38194 19224 38200 19236
rect 38151 19196 38200 19224
rect 38151 19193 38163 19196
rect 38105 19187 38163 19193
rect 38194 19184 38200 19196
rect 38252 19184 38258 19236
rect 41414 19224 41420 19236
rect 41375 19196 41420 19224
rect 41414 19184 41420 19196
rect 41472 19184 41478 19236
rect 41509 19227 41567 19233
rect 41509 19193 41521 19227
rect 41555 19193 41567 19227
rect 41509 19187 41567 19193
rect 42061 19227 42119 19233
rect 42061 19193 42073 19227
rect 42107 19224 42119 19227
rect 42766 19224 42794 19332
rect 43254 19320 43260 19332
rect 43312 19360 43318 19372
rect 43622 19360 43628 19372
rect 43312 19332 43628 19360
rect 43312 19320 43318 19332
rect 43622 19320 43628 19332
rect 43680 19320 43686 19372
rect 42978 19224 42984 19236
rect 42107 19196 42794 19224
rect 42939 19196 42984 19224
rect 42107 19193 42119 19196
rect 42061 19187 42119 19193
rect 31478 19156 31484 19168
rect 26108 19128 26372 19156
rect 31439 19128 31484 19156
rect 26108 19116 26114 19128
rect 31478 19116 31484 19128
rect 31536 19116 31542 19168
rect 31938 19156 31944 19168
rect 31899 19128 31944 19156
rect 31938 19116 31944 19128
rect 31996 19116 32002 19168
rect 32398 19116 32404 19168
rect 32456 19156 32462 19168
rect 32493 19159 32551 19165
rect 32493 19156 32505 19159
rect 32456 19128 32505 19156
rect 32456 19116 32462 19128
rect 32493 19125 32505 19128
rect 32539 19125 32551 19159
rect 32493 19119 32551 19125
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 33229 19159 33287 19165
rect 33229 19156 33241 19159
rect 33192 19128 33241 19156
rect 33192 19116 33198 19128
rect 33229 19125 33241 19128
rect 33275 19156 33287 19159
rect 33410 19156 33416 19168
rect 33275 19128 33416 19156
rect 33275 19125 33287 19128
rect 33229 19119 33287 19125
rect 33410 19116 33416 19128
rect 33468 19116 33474 19168
rect 33594 19156 33600 19168
rect 33555 19128 33600 19156
rect 33594 19116 33600 19128
rect 33652 19116 33658 19168
rect 33870 19156 33876 19168
rect 33831 19128 33876 19156
rect 33870 19116 33876 19128
rect 33928 19116 33934 19168
rect 34514 19156 34520 19168
rect 34475 19128 34520 19156
rect 34514 19116 34520 19128
rect 34572 19116 34578 19168
rect 35618 19116 35624 19168
rect 35676 19156 35682 19168
rect 35805 19159 35863 19165
rect 35805 19156 35817 19159
rect 35676 19128 35817 19156
rect 35676 19116 35682 19128
rect 35805 19125 35817 19128
rect 35851 19125 35863 19159
rect 35805 19119 35863 19125
rect 37277 19159 37335 19165
rect 37277 19125 37289 19159
rect 37323 19156 37335 19159
rect 37568 19156 37596 19184
rect 37323 19128 37596 19156
rect 41233 19159 41291 19165
rect 37323 19125 37335 19128
rect 37277 19119 37335 19125
rect 41233 19125 41245 19159
rect 41279 19156 41291 19159
rect 41322 19156 41328 19168
rect 41279 19128 41328 19156
rect 41279 19125 41291 19128
rect 41233 19119 41291 19125
rect 41322 19116 41328 19128
rect 41380 19156 41386 19168
rect 41524 19156 41552 19187
rect 42978 19184 42984 19196
rect 43036 19184 43042 19236
rect 43073 19227 43131 19233
rect 43073 19193 43085 19227
rect 43119 19193 43131 19227
rect 43073 19187 43131 19193
rect 41380 19128 41552 19156
rect 41380 19116 41386 19128
rect 42610 19116 42616 19168
rect 42668 19156 42674 19168
rect 42705 19159 42763 19165
rect 42705 19156 42717 19159
rect 42668 19128 42717 19156
rect 42668 19116 42674 19128
rect 42705 19125 42717 19128
rect 42751 19156 42763 19159
rect 43088 19156 43116 19187
rect 43438 19184 43444 19236
rect 43496 19224 43502 19236
rect 44361 19227 44419 19233
rect 44361 19224 44373 19227
rect 43496 19196 44373 19224
rect 43496 19184 43502 19196
rect 44361 19193 44373 19196
rect 44407 19224 44419 19227
rect 45186 19224 45192 19236
rect 44407 19196 45192 19224
rect 44407 19193 44419 19196
rect 44361 19187 44419 19193
rect 45186 19184 45192 19196
rect 45244 19224 45250 19236
rect 46750 19224 46756 19236
rect 45244 19196 46756 19224
rect 45244 19184 45250 19196
rect 46750 19184 46756 19196
rect 46808 19184 46814 19236
rect 42751 19128 43116 19156
rect 42751 19125 42763 19128
rect 42705 19119 42763 19125
rect 43714 19116 43720 19168
rect 43772 19156 43778 19168
rect 43901 19159 43959 19165
rect 43901 19156 43913 19159
rect 43772 19128 43913 19156
rect 43772 19116 43778 19128
rect 43901 19125 43913 19128
rect 43947 19125 43959 19159
rect 45002 19156 45008 19168
rect 44963 19128 45008 19156
rect 43901 19119 43959 19125
rect 45002 19116 45008 19128
rect 45060 19116 45066 19168
rect 1104 19066 48852 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 48852 19066
rect 1104 18992 48852 19014
rect 16482 18952 16488 18964
rect 16443 18924 16488 18952
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 16850 18952 16856 18964
rect 16811 18924 16856 18952
rect 16850 18912 16856 18924
rect 16908 18952 16914 18964
rect 17402 18952 17408 18964
rect 16908 18924 17408 18952
rect 16908 18912 16914 18924
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 17770 18952 17776 18964
rect 17731 18924 17776 18952
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 18506 18912 18512 18964
rect 18564 18952 18570 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18564 18924 18613 18952
rect 18564 18912 18570 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 18601 18915 18659 18921
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 28994 18952 29000 18964
rect 28955 18924 29000 18952
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 32030 18952 32036 18964
rect 29104 18924 32036 18952
rect 21177 18887 21235 18893
rect 21177 18853 21189 18887
rect 21223 18884 21235 18887
rect 21358 18884 21364 18896
rect 21223 18856 21364 18884
rect 21223 18853 21235 18856
rect 21177 18847 21235 18853
rect 21358 18844 21364 18856
rect 21416 18844 21422 18896
rect 21542 18844 21548 18896
rect 21600 18884 21606 18896
rect 21729 18887 21787 18893
rect 21729 18884 21741 18887
rect 21600 18856 21741 18884
rect 21600 18844 21606 18856
rect 21729 18853 21741 18856
rect 21775 18853 21787 18887
rect 21729 18847 21787 18853
rect 23385 18887 23443 18893
rect 23385 18853 23397 18887
rect 23431 18884 23443 18887
rect 23676 18884 23704 18912
rect 23431 18856 23704 18884
rect 25593 18887 25651 18893
rect 23431 18853 23443 18856
rect 23385 18847 23443 18853
rect 25593 18853 25605 18887
rect 25639 18884 25651 18887
rect 26694 18884 26700 18896
rect 25639 18856 26700 18884
rect 25639 18853 25651 18856
rect 25593 18847 25651 18853
rect 26694 18844 26700 18856
rect 26752 18844 26758 18896
rect 27798 18844 27804 18896
rect 27856 18884 27862 18896
rect 27893 18887 27951 18893
rect 27893 18884 27905 18887
rect 27856 18856 27905 18884
rect 27856 18844 27862 18856
rect 27893 18853 27905 18856
rect 27939 18884 27951 18887
rect 29104 18884 29132 18924
rect 30576 18896 30604 18924
rect 32030 18912 32036 18924
rect 32088 18912 32094 18964
rect 32398 18912 32404 18964
rect 32456 18952 32462 18964
rect 34606 18952 34612 18964
rect 32456 18924 34612 18952
rect 32456 18912 32462 18924
rect 34606 18912 34612 18924
rect 34664 18912 34670 18964
rect 34790 18912 34796 18964
rect 34848 18952 34854 18964
rect 34977 18955 35035 18961
rect 34977 18952 34989 18955
rect 34848 18924 34989 18952
rect 34848 18912 34854 18924
rect 34977 18921 34989 18924
rect 35023 18921 35035 18955
rect 35342 18952 35348 18964
rect 35303 18924 35348 18952
rect 34977 18915 35035 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 37550 18912 37556 18964
rect 37608 18952 37614 18964
rect 38657 18955 38715 18961
rect 38657 18952 38669 18955
rect 37608 18924 38669 18952
rect 37608 18912 37614 18924
rect 38657 18921 38669 18924
rect 38703 18921 38715 18955
rect 38657 18915 38715 18921
rect 41598 18912 41604 18964
rect 41656 18952 41662 18964
rect 41969 18955 42027 18961
rect 41969 18952 41981 18955
rect 41656 18924 41981 18952
rect 41656 18912 41662 18924
rect 41969 18921 41981 18924
rect 42015 18921 42027 18955
rect 41969 18915 42027 18921
rect 42981 18955 43039 18961
rect 42981 18921 42993 18955
rect 43027 18952 43039 18955
rect 43162 18952 43168 18964
rect 43027 18924 43168 18952
rect 43027 18921 43039 18924
rect 42981 18915 43039 18921
rect 43162 18912 43168 18924
rect 43220 18912 43226 18964
rect 43947 18955 44005 18961
rect 43947 18921 43959 18955
rect 43993 18952 44005 18955
rect 43993 18924 46520 18952
rect 43993 18921 44005 18924
rect 43947 18915 44005 18921
rect 46492 18896 46520 18924
rect 27939 18856 29132 18884
rect 29181 18887 29239 18893
rect 27939 18853 27951 18856
rect 27893 18847 27951 18853
rect 29181 18853 29193 18887
rect 29227 18884 29239 18887
rect 29822 18884 29828 18896
rect 29227 18856 29828 18884
rect 29227 18853 29239 18856
rect 29181 18847 29239 18853
rect 29822 18844 29828 18856
rect 29880 18844 29886 18896
rect 30558 18884 30564 18896
rect 30471 18856 30564 18884
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 34698 18884 34704 18896
rect 30760 18856 32352 18884
rect 34659 18856 34704 18884
rect 30760 18828 30788 18856
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 17184 18788 17417 18816
rect 17184 18776 17190 18788
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19832 18819 19890 18825
rect 19832 18816 19844 18819
rect 19484 18788 19844 18816
rect 19484 18776 19490 18788
rect 19832 18785 19844 18788
rect 19878 18785 19890 18819
rect 19832 18779 19890 18785
rect 22738 18776 22744 18828
rect 22796 18816 22802 18828
rect 23106 18816 23112 18828
rect 22796 18788 23112 18816
rect 22796 18776 22802 18788
rect 23106 18776 23112 18788
rect 23164 18776 23170 18828
rect 25038 18816 25044 18828
rect 24999 18788 25044 18816
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 28169 18819 28227 18825
rect 28169 18785 28181 18819
rect 28215 18816 28227 18819
rect 28350 18816 28356 18828
rect 28215 18788 28356 18816
rect 28215 18785 28227 18788
rect 28169 18779 28227 18785
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 29270 18776 29276 18828
rect 29328 18816 29334 18828
rect 29365 18819 29423 18825
rect 29365 18816 29377 18819
rect 29328 18788 29377 18816
rect 29328 18776 29334 18788
rect 29365 18785 29377 18788
rect 29411 18785 29423 18819
rect 30742 18816 30748 18828
rect 30655 18788 30748 18816
rect 29365 18779 29423 18785
rect 30742 18776 30748 18788
rect 30800 18776 30806 18828
rect 31846 18776 31852 18828
rect 31904 18816 31910 18828
rect 32324 18825 32352 18856
rect 34698 18844 34704 18856
rect 34756 18844 34762 18896
rect 35618 18844 35624 18896
rect 35676 18884 35682 18896
rect 35713 18887 35771 18893
rect 35713 18884 35725 18887
rect 35676 18856 35725 18884
rect 35676 18844 35682 18856
rect 35713 18853 35725 18856
rect 35759 18853 35771 18887
rect 35713 18847 35771 18853
rect 37461 18887 37519 18893
rect 37461 18853 37473 18887
rect 37507 18884 37519 18887
rect 37642 18884 37648 18896
rect 37507 18856 37648 18884
rect 37507 18853 37519 18856
rect 37461 18847 37519 18853
rect 37642 18844 37648 18856
rect 37700 18844 37706 18896
rect 38010 18884 38016 18896
rect 37971 18856 38016 18884
rect 38010 18844 38016 18856
rect 38068 18844 38074 18896
rect 40954 18844 40960 18896
rect 41012 18884 41018 18896
rect 41094 18887 41152 18893
rect 41094 18884 41106 18887
rect 41012 18856 41106 18884
rect 41012 18844 41018 18856
rect 41094 18853 41106 18856
rect 41140 18884 41152 18887
rect 43622 18884 43628 18896
rect 41140 18856 43628 18884
rect 41140 18853 41152 18856
rect 41094 18847 41152 18853
rect 43622 18844 43628 18856
rect 43680 18844 43686 18896
rect 45005 18887 45063 18893
rect 45005 18853 45017 18887
rect 45051 18884 45063 18887
rect 45094 18884 45100 18896
rect 45051 18856 45100 18884
rect 45051 18853 45063 18856
rect 45005 18847 45063 18853
rect 45094 18844 45100 18856
rect 45152 18844 45158 18896
rect 45554 18884 45560 18896
rect 45515 18856 45560 18884
rect 45554 18844 45560 18856
rect 45612 18844 45618 18896
rect 46474 18884 46480 18896
rect 46387 18856 46480 18884
rect 46474 18844 46480 18856
rect 46532 18844 46538 18896
rect 46566 18844 46572 18896
rect 46624 18884 46630 18896
rect 46624 18856 46669 18884
rect 46624 18844 46630 18856
rect 32125 18819 32183 18825
rect 32125 18816 32137 18819
rect 31904 18788 32137 18816
rect 31904 18776 31910 18788
rect 32125 18785 32137 18788
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 32309 18819 32367 18825
rect 32309 18785 32321 18819
rect 32355 18816 32367 18819
rect 32766 18816 32772 18828
rect 32355 18788 32772 18816
rect 32355 18785 32367 18788
rect 32309 18779 32367 18785
rect 32766 18776 32772 18788
rect 32824 18776 32830 18828
rect 33502 18816 33508 18828
rect 33415 18788 33508 18816
rect 33502 18776 33508 18788
rect 33560 18816 33566 18828
rect 34241 18819 34299 18825
rect 34241 18816 34253 18819
rect 33560 18788 34253 18816
rect 33560 18776 33566 18788
rect 34241 18785 34253 18788
rect 34287 18816 34299 18819
rect 34330 18816 34336 18828
rect 34287 18788 34336 18816
rect 34287 18785 34299 18788
rect 34241 18779 34299 18785
rect 34330 18776 34336 18788
rect 34388 18776 34394 18828
rect 34517 18819 34575 18825
rect 34517 18785 34529 18819
rect 34563 18785 34575 18819
rect 34517 18779 34575 18785
rect 36265 18819 36323 18825
rect 36265 18785 36277 18819
rect 36311 18816 36323 18819
rect 38194 18816 38200 18828
rect 36311 18788 38200 18816
rect 36311 18785 36323 18788
rect 36265 18779 36323 18785
rect 19935 18751 19993 18757
rect 19935 18717 19947 18751
rect 19981 18748 19993 18751
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 19981 18720 21097 18748
rect 19981 18717 19993 18720
rect 19935 18711 19993 18717
rect 21085 18717 21097 18720
rect 21131 18748 21143 18751
rect 21542 18748 21548 18760
rect 21131 18720 21548 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 26602 18748 26608 18760
rect 26563 18720 26608 18748
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 27249 18751 27307 18757
rect 27249 18717 27261 18751
rect 27295 18748 27307 18751
rect 27614 18748 27620 18760
rect 27295 18720 27620 18748
rect 27295 18717 27307 18720
rect 27249 18711 27307 18717
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 30834 18708 30840 18760
rect 30892 18748 30898 18760
rect 31389 18751 31447 18757
rect 31389 18748 31401 18751
rect 30892 18720 31401 18748
rect 30892 18708 30898 18720
rect 31389 18717 31401 18720
rect 31435 18717 31447 18751
rect 31389 18711 31447 18717
rect 22557 18683 22615 18689
rect 22557 18649 22569 18683
rect 22603 18680 22615 18683
rect 22738 18680 22744 18692
rect 22603 18652 22744 18680
rect 22603 18649 22615 18652
rect 22557 18643 22615 18649
rect 22738 18640 22744 18652
rect 22796 18680 22802 18692
rect 28353 18683 28411 18689
rect 28353 18680 28365 18683
rect 22796 18652 28365 18680
rect 22796 18640 22802 18652
rect 28353 18649 28365 18652
rect 28399 18680 28411 18683
rect 31478 18680 31484 18692
rect 28399 18652 31484 18680
rect 28399 18649 28411 18652
rect 28353 18643 28411 18649
rect 31478 18640 31484 18652
rect 31536 18640 31542 18692
rect 34054 18640 34060 18692
rect 34112 18680 34118 18692
rect 34532 18680 34560 18779
rect 38194 18776 38200 18788
rect 38252 18816 38258 18828
rect 39552 18819 39610 18825
rect 39552 18816 39564 18819
rect 38252 18788 39564 18816
rect 38252 18776 38258 18788
rect 39552 18785 39564 18788
rect 39598 18816 39610 18819
rect 39942 18816 39948 18828
rect 39598 18788 39948 18816
rect 39598 18785 39610 18788
rect 39552 18779 39610 18785
rect 39942 18776 39948 18788
rect 40000 18776 40006 18828
rect 40034 18776 40040 18828
rect 40092 18816 40098 18828
rect 40773 18819 40831 18825
rect 40773 18816 40785 18819
rect 40092 18788 40785 18816
rect 40092 18776 40098 18788
rect 40773 18785 40785 18788
rect 40819 18816 40831 18819
rect 41690 18816 41696 18828
rect 40819 18788 41696 18816
rect 40819 18785 40831 18788
rect 40773 18779 40831 18785
rect 41690 18776 41696 18788
rect 41748 18776 41754 18828
rect 42794 18776 42800 18828
rect 42852 18816 42858 18828
rect 43844 18819 43902 18825
rect 43844 18816 43856 18819
rect 42852 18788 43856 18816
rect 42852 18776 42858 18788
rect 43844 18785 43856 18788
rect 43890 18785 43902 18819
rect 43844 18779 43902 18785
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 35621 18751 35679 18757
rect 35621 18748 35633 18751
rect 35400 18720 35633 18748
rect 35400 18708 35406 18720
rect 35621 18717 35633 18720
rect 35667 18717 35679 18751
rect 37734 18748 37740 18760
rect 37695 18720 37740 18748
rect 35621 18711 35679 18717
rect 37734 18708 37740 18720
rect 37792 18708 37798 18760
rect 43714 18748 43720 18760
rect 42029 18720 43720 18748
rect 41693 18683 41751 18689
rect 34112 18652 36676 18680
rect 34112 18640 34118 18652
rect 18322 18612 18328 18624
rect 18283 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 20533 18615 20591 18621
rect 20533 18581 20545 18615
rect 20579 18612 20591 18615
rect 20714 18612 20720 18624
rect 20579 18584 20720 18612
rect 20579 18581 20591 18584
rect 20533 18575 20591 18581
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 26234 18612 26240 18624
rect 26195 18584 26240 18612
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 27890 18572 27896 18624
rect 27948 18612 27954 18624
rect 29457 18615 29515 18621
rect 29457 18612 29469 18615
rect 27948 18584 29469 18612
rect 27948 18572 27954 18584
rect 29457 18581 29469 18584
rect 29503 18581 29515 18615
rect 29457 18575 29515 18581
rect 29546 18572 29552 18624
rect 29604 18612 29610 18624
rect 30837 18615 30895 18621
rect 30837 18612 30849 18615
rect 29604 18584 30849 18612
rect 29604 18572 29610 18584
rect 30837 18581 30849 18584
rect 30883 18581 30895 18615
rect 30837 18575 30895 18581
rect 32306 18572 32312 18624
rect 32364 18612 32370 18624
rect 36648 18621 36676 18652
rect 41693 18649 41705 18683
rect 41739 18680 41751 18683
rect 42029 18680 42057 18720
rect 43714 18708 43720 18720
rect 43772 18708 43778 18760
rect 44910 18748 44916 18760
rect 44871 18720 44916 18748
rect 44910 18708 44916 18720
rect 44968 18708 44974 18760
rect 46750 18748 46756 18760
rect 46711 18720 46756 18748
rect 46750 18708 46756 18720
rect 46808 18708 46814 18760
rect 41739 18652 42057 18680
rect 41739 18649 41751 18652
rect 41693 18643 41751 18649
rect 32401 18615 32459 18621
rect 32401 18612 32413 18615
rect 32364 18584 32413 18612
rect 32364 18572 32370 18584
rect 32401 18581 32413 18584
rect 32447 18581 32459 18615
rect 32401 18575 32459 18581
rect 36633 18615 36691 18621
rect 36633 18581 36645 18615
rect 36679 18612 36691 18615
rect 36814 18612 36820 18624
rect 36679 18584 36820 18612
rect 36679 18581 36691 18584
rect 36633 18575 36691 18581
rect 36814 18572 36820 18584
rect 36872 18572 36878 18624
rect 39623 18615 39681 18621
rect 39623 18581 39635 18615
rect 39669 18612 39681 18615
rect 39758 18612 39764 18624
rect 39669 18584 39764 18612
rect 39669 18581 39681 18584
rect 39623 18575 39681 18581
rect 39758 18572 39764 18584
rect 39816 18572 39822 18624
rect 40494 18612 40500 18624
rect 40455 18584 40500 18612
rect 40494 18572 40500 18584
rect 40552 18572 40558 18624
rect 43622 18612 43628 18624
rect 43583 18584 43628 18612
rect 43622 18572 43628 18584
rect 43680 18572 43686 18624
rect 1104 18522 48852 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 48852 18522
rect 1104 18448 48852 18470
rect 17126 18408 17132 18420
rect 17087 18380 17132 18408
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 17497 18411 17555 18417
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 17770 18408 17776 18420
rect 17543 18380 17776 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 21269 18411 21327 18417
rect 21269 18377 21281 18411
rect 21315 18408 21327 18411
rect 21358 18408 21364 18420
rect 21315 18380 21364 18408
rect 21315 18377 21327 18380
rect 21269 18371 21327 18377
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 21542 18408 21548 18420
rect 21503 18380 21548 18408
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 22738 18408 22744 18420
rect 22699 18380 22744 18408
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23106 18408 23112 18420
rect 23067 18380 23112 18408
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 24857 18411 24915 18417
rect 24857 18377 24869 18411
rect 24903 18408 24915 18411
rect 24946 18408 24952 18420
rect 24903 18380 24952 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 25130 18408 25136 18420
rect 25091 18380 25136 18408
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 25590 18408 25596 18420
rect 25551 18380 25596 18408
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 26694 18408 26700 18420
rect 26655 18380 26700 18408
rect 26694 18368 26700 18380
rect 26752 18368 26758 18420
rect 29089 18411 29147 18417
rect 29089 18377 29101 18411
rect 29135 18408 29147 18411
rect 29270 18408 29276 18420
rect 29135 18380 29276 18408
rect 29135 18377 29147 18380
rect 29089 18371 29147 18377
rect 29270 18368 29276 18380
rect 29328 18368 29334 18420
rect 30469 18411 30527 18417
rect 30469 18377 30481 18411
rect 30515 18408 30527 18411
rect 30742 18408 30748 18420
rect 30515 18380 30748 18408
rect 30515 18377 30527 18380
rect 30469 18371 30527 18377
rect 30742 18368 30748 18380
rect 30800 18368 30806 18420
rect 31846 18408 31852 18420
rect 31807 18380 31852 18408
rect 31846 18368 31852 18380
rect 31904 18368 31910 18420
rect 36265 18411 36323 18417
rect 36265 18377 36277 18411
rect 36311 18408 36323 18411
rect 36446 18408 36452 18420
rect 36311 18380 36452 18408
rect 36311 18377 36323 18380
rect 36265 18371 36323 18377
rect 36446 18368 36452 18380
rect 36504 18368 36510 18420
rect 37461 18411 37519 18417
rect 37461 18377 37473 18411
rect 37507 18408 37519 18411
rect 37734 18408 37740 18420
rect 37507 18380 37740 18408
rect 37507 18377 37519 18380
rect 37461 18371 37519 18377
rect 18690 18340 18696 18352
rect 18651 18312 18696 18340
rect 18690 18300 18696 18312
rect 18748 18300 18754 18352
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18272 18199 18275
rect 18506 18272 18512 18284
rect 18187 18244 18512 18272
rect 18187 18241 18199 18244
rect 18141 18235 18199 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 20714 18272 20720 18284
rect 20675 18244 20720 18272
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 23124 18272 23152 18368
rect 24581 18343 24639 18349
rect 24581 18309 24593 18343
rect 24627 18340 24639 18343
rect 25038 18340 25044 18352
rect 24627 18312 25044 18340
rect 24627 18309 24639 18312
rect 24581 18303 24639 18309
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 29178 18300 29184 18352
rect 29236 18340 29242 18352
rect 34790 18340 34796 18352
rect 29236 18312 34796 18340
rect 29236 18300 29242 18312
rect 34790 18300 34796 18312
rect 34848 18300 34854 18352
rect 27614 18272 27620 18284
rect 21376 18244 23152 18272
rect 27575 18244 27620 18272
rect 19978 18164 19984 18216
rect 20036 18204 20042 18216
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 20036 18176 20177 18204
rect 20036 18164 20042 18176
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18204 20683 18207
rect 21376 18204 21404 18244
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 29822 18272 29828 18284
rect 29735 18244 29828 18272
rect 29822 18232 29828 18244
rect 29880 18272 29886 18284
rect 31846 18272 31852 18284
rect 29880 18244 31852 18272
rect 29880 18232 29886 18244
rect 31846 18232 31852 18244
rect 31904 18232 31910 18284
rect 32493 18275 32551 18281
rect 32493 18241 32505 18275
rect 32539 18272 32551 18275
rect 32858 18272 32864 18284
rect 32539 18244 32864 18272
rect 32539 18241 32551 18244
rect 32493 18235 32551 18241
rect 32858 18232 32864 18244
rect 32916 18272 32922 18284
rect 33226 18272 33232 18284
rect 32916 18244 33232 18272
rect 32916 18232 32922 18244
rect 33226 18232 33232 18244
rect 33284 18232 33290 18284
rect 37093 18275 37151 18281
rect 33428 18244 35112 18272
rect 20671 18176 21404 18204
rect 21729 18207 21787 18213
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 21729 18173 21741 18207
rect 21775 18204 21787 18207
rect 21775 18176 22324 18204
rect 21775 18173 21787 18176
rect 21729 18167 21787 18173
rect 18233 18139 18291 18145
rect 18233 18105 18245 18139
rect 18279 18136 18291 18139
rect 18322 18136 18328 18148
rect 18279 18108 18328 18136
rect 18279 18105 18291 18108
rect 18233 18099 18291 18105
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18248 18068 18276 18099
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 19705 18139 19763 18145
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 20070 18136 20076 18148
rect 19751 18108 20076 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 20070 18096 20076 18108
rect 20128 18136 20134 18148
rect 20640 18136 20668 18167
rect 20128 18108 20668 18136
rect 20128 18096 20134 18108
rect 22296 18080 22324 18176
rect 22554 18164 22560 18216
rect 22612 18204 22618 18216
rect 23728 18207 23786 18213
rect 23728 18204 23740 18207
rect 22612 18176 23740 18204
rect 22612 18164 22618 18176
rect 23728 18173 23740 18176
rect 23774 18204 23786 18207
rect 24673 18207 24731 18213
rect 23774 18176 24256 18204
rect 23774 18173 23786 18176
rect 23728 18167 23786 18173
rect 24228 18080 24256 18176
rect 24673 18173 24685 18207
rect 24719 18204 24731 18207
rect 25130 18204 25136 18216
rect 24719 18176 25136 18204
rect 24719 18173 24731 18176
rect 24673 18167 24731 18173
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 28721 18207 28779 18213
rect 28721 18173 28733 18207
rect 28767 18204 28779 18207
rect 29273 18207 29331 18213
rect 29273 18204 29285 18207
rect 28767 18176 29285 18204
rect 28767 18173 28779 18176
rect 28721 18167 28779 18173
rect 29273 18173 29285 18176
rect 29319 18204 29331 18207
rect 29546 18204 29552 18216
rect 29319 18176 29552 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 29546 18164 29552 18176
rect 29604 18164 29610 18216
rect 30745 18207 30803 18213
rect 30745 18173 30757 18207
rect 30791 18204 30803 18207
rect 30834 18204 30840 18216
rect 30791 18176 30840 18204
rect 30791 18173 30803 18176
rect 30745 18167 30803 18173
rect 30834 18164 30840 18176
rect 30892 18164 30898 18216
rect 32125 18207 32183 18213
rect 32125 18173 32137 18207
rect 32171 18204 32183 18207
rect 32398 18204 32404 18216
rect 32171 18176 32404 18204
rect 32171 18173 32183 18176
rect 32125 18167 32183 18173
rect 32398 18164 32404 18176
rect 32456 18164 32462 18216
rect 32766 18204 32772 18216
rect 32679 18176 32772 18204
rect 32766 18164 32772 18176
rect 32824 18204 32830 18216
rect 33428 18204 33456 18244
rect 32824 18176 33456 18204
rect 33505 18207 33563 18213
rect 32824 18164 32830 18176
rect 33505 18173 33517 18207
rect 33551 18204 33563 18207
rect 33551 18176 34284 18204
rect 33551 18173 33563 18176
rect 33505 18167 33563 18173
rect 25774 18136 25780 18148
rect 25735 18108 25780 18136
rect 25774 18096 25780 18108
rect 25832 18096 25838 18148
rect 25869 18139 25927 18145
rect 25869 18105 25881 18139
rect 25915 18105 25927 18139
rect 25869 18099 25927 18105
rect 17911 18040 18276 18068
rect 19337 18071 19395 18077
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19426 18068 19432 18080
rect 19383 18040 19432 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19978 18068 19984 18080
rect 19939 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 21910 18068 21916 18080
rect 21871 18040 21916 18068
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22278 18068 22284 18080
rect 22239 18040 22284 18068
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 23799 18071 23857 18077
rect 23799 18037 23811 18071
rect 23845 18068 23857 18071
rect 23934 18068 23940 18080
rect 23845 18040 23940 18068
rect 23845 18037 23857 18040
rect 23799 18031 23857 18037
rect 23934 18028 23940 18040
rect 23992 18028 23998 18080
rect 24210 18068 24216 18080
rect 24171 18040 24216 18068
rect 24210 18028 24216 18040
rect 24268 18028 24274 18080
rect 25590 18028 25596 18080
rect 25648 18068 25654 18080
rect 25884 18068 25912 18099
rect 26234 18096 26240 18148
rect 26292 18136 26298 18148
rect 26421 18139 26479 18145
rect 26421 18136 26433 18139
rect 26292 18108 26433 18136
rect 26292 18096 26298 18108
rect 26421 18105 26433 18108
rect 26467 18136 26479 18139
rect 26786 18136 26792 18148
rect 26467 18108 26792 18136
rect 26467 18105 26479 18108
rect 26421 18099 26479 18105
rect 26786 18096 26792 18108
rect 26844 18096 26850 18148
rect 27338 18136 27344 18148
rect 27299 18108 27344 18136
rect 27338 18096 27344 18108
rect 27396 18096 27402 18148
rect 27433 18139 27491 18145
rect 27433 18105 27445 18139
rect 27479 18105 27491 18139
rect 27433 18099 27491 18105
rect 30561 18139 30619 18145
rect 30561 18105 30573 18139
rect 30607 18105 30619 18139
rect 31110 18136 31116 18148
rect 31071 18108 31116 18136
rect 30561 18099 30619 18105
rect 27065 18071 27123 18077
rect 27065 18068 27077 18071
rect 25648 18040 27077 18068
rect 25648 18028 25654 18040
rect 27065 18037 27077 18040
rect 27111 18068 27123 18071
rect 27448 18068 27476 18099
rect 28350 18068 28356 18080
rect 27111 18040 27476 18068
rect 28311 18040 28356 18068
rect 27111 18037 27123 18040
rect 27065 18031 27123 18037
rect 28350 18028 28356 18040
rect 28408 18028 28414 18080
rect 29362 18028 29368 18080
rect 29420 18068 29426 18080
rect 29457 18071 29515 18077
rect 29457 18068 29469 18071
rect 29420 18040 29469 18068
rect 29420 18028 29426 18040
rect 29457 18037 29469 18040
rect 29503 18037 29515 18071
rect 30576 18068 30604 18099
rect 31110 18096 31116 18108
rect 31168 18096 31174 18148
rect 31202 18096 31208 18148
rect 31260 18136 31266 18148
rect 31941 18139 31999 18145
rect 31941 18136 31953 18139
rect 31260 18108 31953 18136
rect 31260 18096 31266 18108
rect 31941 18105 31953 18108
rect 31987 18136 31999 18139
rect 33229 18139 33287 18145
rect 33229 18136 33241 18139
rect 31987 18108 33241 18136
rect 31987 18105 31999 18108
rect 31941 18099 31999 18105
rect 33229 18105 33241 18108
rect 33275 18136 33287 18139
rect 33318 18136 33324 18148
rect 33275 18108 33324 18136
rect 33275 18105 33287 18108
rect 33229 18099 33287 18105
rect 33318 18096 33324 18108
rect 33376 18096 33382 18148
rect 34256 18080 34284 18176
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 35084 18213 35112 18244
rect 37093 18241 37105 18275
rect 37139 18272 37151 18275
rect 37476 18272 37504 18371
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 38381 18411 38439 18417
rect 38381 18377 38393 18411
rect 38427 18408 38439 18411
rect 38930 18408 38936 18420
rect 38427 18380 38936 18408
rect 38427 18377 38439 18380
rect 38381 18371 38439 18377
rect 38930 18368 38936 18380
rect 38988 18368 38994 18420
rect 41322 18368 41328 18420
rect 41380 18408 41386 18420
rect 41417 18411 41475 18417
rect 41417 18408 41429 18411
rect 41380 18380 41429 18408
rect 41380 18368 41386 18380
rect 41417 18377 41429 18380
rect 41463 18377 41475 18411
rect 41690 18408 41696 18420
rect 41651 18380 41696 18408
rect 41417 18371 41475 18377
rect 41690 18368 41696 18380
rect 41748 18368 41754 18420
rect 42794 18368 42800 18420
rect 42852 18408 42858 18420
rect 43349 18411 43407 18417
rect 43349 18408 43361 18411
rect 42852 18380 43361 18408
rect 42852 18368 42858 18380
rect 43349 18377 43361 18380
rect 43395 18377 43407 18411
rect 43349 18371 43407 18377
rect 45002 18368 45008 18420
rect 45060 18408 45066 18420
rect 45833 18411 45891 18417
rect 45833 18408 45845 18411
rect 45060 18380 45845 18408
rect 45060 18368 45066 18380
rect 45833 18377 45845 18380
rect 45879 18408 45891 18411
rect 45879 18380 46244 18408
rect 45879 18377 45891 18380
rect 45833 18371 45891 18377
rect 38010 18300 38016 18352
rect 38068 18340 38074 18352
rect 39853 18343 39911 18349
rect 39853 18340 39865 18343
rect 38068 18312 39865 18340
rect 38068 18300 38074 18312
rect 39853 18309 39865 18312
rect 39899 18340 39911 18343
rect 40221 18343 40279 18349
rect 40221 18340 40233 18343
rect 39899 18312 40233 18340
rect 39899 18309 39911 18312
rect 39853 18303 39911 18309
rect 40221 18309 40233 18312
rect 40267 18309 40279 18343
rect 44910 18340 44916 18352
rect 40221 18303 40279 18309
rect 42766 18312 44916 18340
rect 37139 18244 37504 18272
rect 37139 18241 37151 18244
rect 37093 18235 37151 18241
rect 37550 18232 37556 18284
rect 37608 18272 37614 18284
rect 39206 18272 39212 18284
rect 37608 18244 39212 18272
rect 37608 18232 37614 18244
rect 39206 18232 39212 18244
rect 39264 18272 39270 18284
rect 42659 18275 42717 18281
rect 39264 18244 42057 18272
rect 39264 18232 39270 18244
rect 34885 18207 34943 18213
rect 34885 18204 34897 18207
rect 34848 18176 34897 18204
rect 34848 18164 34854 18176
rect 34885 18173 34897 18176
rect 34931 18173 34943 18207
rect 34885 18167 34943 18173
rect 35069 18207 35127 18213
rect 35069 18173 35081 18207
rect 35115 18204 35127 18207
rect 35802 18204 35808 18216
rect 35115 18176 35808 18204
rect 35115 18173 35127 18176
rect 35069 18167 35127 18173
rect 35802 18164 35808 18176
rect 35860 18164 35866 18216
rect 36446 18204 36452 18216
rect 36407 18176 36452 18204
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 36814 18204 36820 18216
rect 36775 18176 36820 18204
rect 36814 18164 36820 18176
rect 36872 18164 36878 18216
rect 36906 18164 36912 18216
rect 36964 18204 36970 18216
rect 38749 18207 38807 18213
rect 38749 18204 38761 18207
rect 36964 18176 38761 18204
rect 36964 18164 36970 18176
rect 38749 18173 38761 18176
rect 38795 18204 38807 18207
rect 38841 18207 38899 18213
rect 38841 18204 38853 18207
rect 38795 18176 38853 18204
rect 38795 18173 38807 18176
rect 38749 18167 38807 18173
rect 38841 18173 38853 18176
rect 38887 18173 38899 18207
rect 38841 18167 38899 18173
rect 38930 18164 38936 18216
rect 38988 18204 38994 18216
rect 39301 18207 39359 18213
rect 39301 18204 39313 18207
rect 38988 18176 39313 18204
rect 38988 18164 38994 18176
rect 39301 18173 39313 18176
rect 39347 18204 39359 18207
rect 39390 18204 39396 18216
rect 39347 18176 39396 18204
rect 39347 18173 39359 18176
rect 39301 18167 39359 18173
rect 39390 18164 39396 18176
rect 39448 18164 39454 18216
rect 39666 18164 39672 18216
rect 39724 18204 39730 18216
rect 40494 18204 40500 18216
rect 39724 18176 40500 18204
rect 39724 18164 39730 18176
rect 40494 18164 40500 18176
rect 40552 18164 40558 18216
rect 42029 18204 42057 18244
rect 42659 18241 42671 18275
rect 42705 18272 42717 18275
rect 42766 18272 42794 18312
rect 44910 18300 44916 18312
rect 44968 18340 44974 18352
rect 45189 18343 45247 18349
rect 45189 18340 45201 18343
rect 44968 18312 45201 18340
rect 44968 18300 44974 18312
rect 45189 18309 45201 18312
rect 45235 18309 45247 18343
rect 45189 18303 45247 18309
rect 42705 18244 42794 18272
rect 43073 18275 43131 18281
rect 42705 18241 42717 18244
rect 42659 18235 42717 18241
rect 43073 18241 43085 18275
rect 43119 18272 43131 18275
rect 43346 18272 43352 18284
rect 43119 18244 43352 18272
rect 43119 18241 43131 18244
rect 43073 18235 43131 18241
rect 42556 18207 42614 18213
rect 42556 18204 42568 18207
rect 42029 18176 42568 18204
rect 42556 18173 42568 18176
rect 42602 18204 42614 18207
rect 43088 18204 43116 18235
rect 43346 18232 43352 18244
rect 43404 18232 43410 18284
rect 43533 18275 43591 18281
rect 43533 18241 43545 18275
rect 43579 18272 43591 18275
rect 43806 18272 43812 18284
rect 43579 18244 43812 18272
rect 43579 18241 43591 18244
rect 43533 18235 43591 18241
rect 43806 18232 43812 18244
rect 43864 18232 43870 18284
rect 46216 18281 46244 18380
rect 46201 18275 46259 18281
rect 46201 18241 46213 18275
rect 46247 18241 46259 18275
rect 46842 18272 46848 18284
rect 46803 18244 46848 18272
rect 46201 18235 46259 18241
rect 46842 18232 46848 18244
rect 46900 18232 46906 18284
rect 42602 18176 43116 18204
rect 42602 18173 42614 18176
rect 42556 18167 42614 18173
rect 43438 18164 43444 18216
rect 43496 18204 43502 18216
rect 45922 18204 45928 18216
rect 43496 18176 45928 18204
rect 43496 18164 43502 18176
rect 45922 18164 45928 18176
rect 45980 18164 45986 18216
rect 35437 18139 35495 18145
rect 35437 18105 35449 18139
rect 35483 18136 35495 18139
rect 37642 18136 37648 18148
rect 35483 18108 37648 18136
rect 35483 18105 35495 18108
rect 35437 18099 35495 18105
rect 37642 18096 37648 18108
rect 37700 18096 37706 18148
rect 37829 18139 37887 18145
rect 37829 18105 37841 18139
rect 37875 18136 37887 18139
rect 38010 18136 38016 18148
rect 37875 18108 38016 18136
rect 37875 18105 37887 18108
rect 37829 18099 37887 18105
rect 38010 18096 38016 18108
rect 38068 18096 38074 18148
rect 39577 18139 39635 18145
rect 39577 18105 39589 18139
rect 39623 18136 39635 18139
rect 40678 18136 40684 18148
rect 39623 18108 40684 18136
rect 39623 18105 39635 18108
rect 39577 18099 39635 18105
rect 40678 18096 40684 18108
rect 40736 18096 40742 18148
rect 40859 18139 40917 18145
rect 40859 18105 40871 18139
rect 40905 18136 40917 18139
rect 40954 18136 40960 18148
rect 40905 18108 40960 18136
rect 40905 18105 40917 18108
rect 40859 18099 40917 18105
rect 40954 18096 40960 18108
rect 41012 18096 41018 18148
rect 43622 18096 43628 18148
rect 43680 18136 43686 18148
rect 43854 18139 43912 18145
rect 43854 18136 43866 18139
rect 43680 18108 43866 18136
rect 43680 18096 43686 18108
rect 43854 18105 43866 18108
rect 43900 18105 43912 18139
rect 43854 18099 43912 18105
rect 46293 18139 46351 18145
rect 46293 18105 46305 18139
rect 46339 18105 46351 18139
rect 46293 18099 46351 18105
rect 31478 18068 31484 18080
rect 30576 18040 31484 18068
rect 29457 18031 29515 18037
rect 31478 18028 31484 18040
rect 31536 18028 31542 18080
rect 33594 18068 33600 18080
rect 33555 18040 33600 18068
rect 33594 18028 33600 18040
rect 33652 18028 33658 18080
rect 34238 18068 34244 18080
rect 34199 18040 34244 18068
rect 34238 18028 34244 18040
rect 34296 18028 34302 18080
rect 34330 18028 34336 18080
rect 34388 18068 34394 18080
rect 34609 18071 34667 18077
rect 34609 18068 34621 18071
rect 34388 18040 34621 18068
rect 34388 18028 34394 18040
rect 34609 18037 34621 18040
rect 34655 18068 34667 18071
rect 35250 18068 35256 18080
rect 34655 18040 35256 18068
rect 34655 18037 34667 18040
rect 34609 18031 34667 18037
rect 35250 18028 35256 18040
rect 35308 18068 35314 18080
rect 38286 18068 38292 18080
rect 35308 18040 38292 18068
rect 35308 18028 35314 18040
rect 38286 18028 38292 18040
rect 38344 18028 38350 18080
rect 44453 18071 44511 18077
rect 44453 18037 44465 18071
rect 44499 18068 44511 18071
rect 44913 18071 44971 18077
rect 44913 18068 44925 18071
rect 44499 18040 44925 18068
rect 44499 18037 44511 18040
rect 44453 18031 44511 18037
rect 44913 18037 44925 18040
rect 44959 18068 44971 18071
rect 45094 18068 45100 18080
rect 44959 18040 45100 18068
rect 44959 18037 44971 18040
rect 44913 18031 44971 18037
rect 45094 18028 45100 18040
rect 45152 18068 45158 18080
rect 46198 18068 46204 18080
rect 45152 18040 46204 18068
rect 45152 18028 45158 18040
rect 46198 18028 46204 18040
rect 46256 18068 46262 18080
rect 46308 18068 46336 18099
rect 46566 18068 46572 18080
rect 46256 18040 46572 18068
rect 46256 18028 46262 18040
rect 46566 18028 46572 18040
rect 46624 18068 46630 18080
rect 47121 18071 47179 18077
rect 47121 18068 47133 18071
rect 46624 18040 47133 18068
rect 46624 18028 46630 18040
rect 47121 18037 47133 18040
rect 47167 18037 47179 18071
rect 47121 18031 47179 18037
rect 1104 17978 48852 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 48852 17978
rect 1104 17904 48852 17926
rect 20990 17864 20996 17876
rect 20951 17836 20996 17864
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 26329 17867 26387 17873
rect 26329 17833 26341 17867
rect 26375 17864 26387 17867
rect 26602 17864 26608 17876
rect 26375 17836 26608 17864
rect 26375 17833 26387 17836
rect 26329 17827 26387 17833
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 27338 17824 27344 17876
rect 27396 17864 27402 17876
rect 27525 17867 27583 17873
rect 27525 17864 27537 17867
rect 27396 17836 27537 17864
rect 27396 17824 27402 17836
rect 27525 17833 27537 17836
rect 27571 17833 27583 17867
rect 27525 17827 27583 17833
rect 28350 17824 28356 17876
rect 28408 17864 28414 17876
rect 32401 17867 32459 17873
rect 32401 17864 32413 17867
rect 28408 17836 32413 17864
rect 28408 17824 28414 17836
rect 32401 17833 32413 17836
rect 32447 17833 32459 17867
rect 33318 17864 33324 17876
rect 33279 17836 33324 17864
rect 32401 17827 32459 17833
rect 33318 17824 33324 17836
rect 33376 17824 33382 17876
rect 34054 17864 34060 17876
rect 34015 17836 34060 17864
rect 34054 17824 34060 17836
rect 34112 17824 34118 17876
rect 35618 17864 35624 17876
rect 35579 17836 35624 17864
rect 35618 17824 35624 17836
rect 35676 17824 35682 17876
rect 36173 17867 36231 17873
rect 36173 17833 36185 17867
rect 36219 17864 36231 17867
rect 36446 17864 36452 17876
rect 36219 17836 36452 17864
rect 36219 17833 36231 17836
rect 36173 17827 36231 17833
rect 36446 17824 36452 17836
rect 36504 17824 36510 17876
rect 39942 17864 39948 17876
rect 39903 17836 39948 17864
rect 39942 17824 39948 17836
rect 40000 17824 40006 17876
rect 40034 17824 40040 17876
rect 40092 17864 40098 17876
rect 43438 17864 43444 17876
rect 40092 17836 43444 17864
rect 40092 17824 40098 17836
rect 43438 17824 43444 17836
rect 43496 17824 43502 17876
rect 43530 17824 43536 17876
rect 43588 17864 43594 17876
rect 46198 17864 46204 17876
rect 43588 17836 45508 17864
rect 46159 17836 46204 17864
rect 43588 17824 43594 17836
rect 17307 17799 17365 17805
rect 17307 17765 17319 17799
rect 17353 17796 17365 17799
rect 17770 17796 17776 17808
rect 17353 17768 17776 17796
rect 17353 17765 17365 17768
rect 17307 17759 17365 17765
rect 17770 17756 17776 17768
rect 17828 17756 17834 17808
rect 26694 17796 26700 17808
rect 19812 17768 21220 17796
rect 26655 17768 26700 17796
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 16945 17731 17003 17737
rect 16945 17728 16957 17731
rect 16908 17700 16957 17728
rect 16908 17688 16914 17700
rect 16945 17697 16957 17700
rect 16991 17728 17003 17731
rect 18138 17728 18144 17740
rect 16991 17700 18144 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 19518 17728 19524 17740
rect 19479 17700 19524 17728
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 19812 17737 19840 17768
rect 21192 17740 21220 17768
rect 26694 17756 26700 17768
rect 26752 17756 26758 17808
rect 26786 17756 26792 17808
rect 26844 17796 26850 17808
rect 27249 17799 27307 17805
rect 27249 17796 27261 17799
rect 26844 17768 27261 17796
rect 26844 17756 26850 17768
rect 27249 17765 27261 17768
rect 27295 17765 27307 17799
rect 29178 17796 29184 17808
rect 29139 17768 29184 17796
rect 27249 17759 27307 17765
rect 29178 17756 29184 17768
rect 29236 17756 29242 17808
rect 30558 17796 30564 17808
rect 30519 17768 30564 17796
rect 30558 17756 30564 17768
rect 30616 17756 30622 17808
rect 31478 17756 31484 17808
rect 31536 17796 31542 17808
rect 32125 17799 32183 17805
rect 32125 17796 32137 17799
rect 31536 17768 32137 17796
rect 31536 17756 31542 17768
rect 32125 17765 32137 17768
rect 32171 17796 32183 17799
rect 32766 17796 32772 17808
rect 32171 17768 32772 17796
rect 32171 17765 32183 17768
rect 32125 17759 32183 17765
rect 32766 17756 32772 17768
rect 32824 17756 32830 17808
rect 36464 17796 36492 17824
rect 45480 17808 45508 17836
rect 46198 17824 46204 17836
rect 46256 17824 46262 17876
rect 46474 17864 46480 17876
rect 46435 17836 46480 17864
rect 46474 17824 46480 17836
rect 46532 17824 46538 17876
rect 38654 17796 38660 17808
rect 36464 17768 38660 17796
rect 38654 17756 38660 17768
rect 38712 17796 38718 17808
rect 39666 17796 39672 17808
rect 38712 17768 38976 17796
rect 39627 17768 39672 17796
rect 38712 17756 38718 17768
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 21085 17731 21143 17737
rect 21085 17697 21097 17731
rect 21131 17697 21143 17731
rect 21085 17691 21143 17697
rect 19886 17660 19892 17672
rect 19847 17632 19892 17660
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 21100 17660 21128 17691
rect 21174 17688 21180 17740
rect 21232 17728 21238 17740
rect 21453 17731 21511 17737
rect 21453 17728 21465 17731
rect 21232 17700 21465 17728
rect 21232 17688 21238 17700
rect 21453 17697 21465 17700
rect 21499 17728 21511 17731
rect 21910 17728 21916 17740
rect 21499 17700 21916 17728
rect 21499 17697 21511 17700
rect 21453 17691 21511 17697
rect 21910 17688 21916 17700
rect 21968 17688 21974 17740
rect 23382 17728 23388 17740
rect 23343 17700 23388 17728
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 24268 17700 24409 17728
rect 24268 17688 24274 17700
rect 24397 17697 24409 17700
rect 24443 17728 24455 17731
rect 25038 17728 25044 17740
rect 24443 17700 25044 17728
rect 24443 17697 24455 17700
rect 24397 17691 24455 17697
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 25409 17731 25467 17737
rect 25409 17697 25421 17731
rect 25455 17728 25467 17731
rect 25498 17728 25504 17740
rect 25455 17700 25504 17728
rect 25455 17697 25467 17700
rect 25409 17691 25467 17697
rect 25498 17688 25504 17700
rect 25556 17688 25562 17740
rect 28077 17731 28135 17737
rect 28077 17697 28089 17731
rect 28123 17728 28135 17731
rect 28258 17728 28264 17740
rect 28123 17700 28264 17728
rect 28123 17697 28135 17700
rect 28077 17691 28135 17697
rect 28258 17688 28264 17700
rect 28316 17688 28322 17740
rect 29270 17688 29276 17740
rect 29328 17728 29334 17740
rect 29365 17731 29423 17737
rect 29365 17728 29377 17731
rect 29328 17700 29377 17728
rect 29328 17688 29334 17700
rect 29365 17697 29377 17700
rect 29411 17697 29423 17731
rect 30650 17728 30656 17740
rect 30611 17700 30656 17728
rect 29365 17691 29423 17697
rect 30650 17688 30656 17700
rect 30708 17688 30714 17740
rect 30834 17728 30840 17740
rect 30795 17700 30840 17728
rect 30834 17688 30840 17700
rect 30892 17688 30898 17740
rect 32214 17688 32220 17740
rect 32272 17728 32278 17740
rect 32309 17731 32367 17737
rect 32309 17728 32321 17731
rect 32272 17700 32321 17728
rect 32272 17688 32278 17700
rect 32309 17697 32321 17700
rect 32355 17697 32367 17731
rect 34514 17728 34520 17740
rect 34475 17700 34520 17728
rect 32309 17691 32367 17697
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 35342 17688 35348 17740
rect 35400 17728 35406 17740
rect 35989 17731 36047 17737
rect 35989 17728 36001 17731
rect 35400 17700 36001 17728
rect 35400 17688 35406 17700
rect 35989 17697 36001 17700
rect 36035 17697 36047 17731
rect 35989 17691 36047 17697
rect 37642 17688 37648 17740
rect 37700 17728 37706 17740
rect 38948 17737 38976 17768
rect 39666 17756 39672 17768
rect 39724 17756 39730 17808
rect 40838 17799 40896 17805
rect 40838 17765 40850 17799
rect 40884 17796 40896 17799
rect 40954 17796 40960 17808
rect 40884 17768 40960 17796
rect 40884 17765 40896 17768
rect 40838 17759 40896 17765
rect 40954 17756 40960 17768
rect 41012 17756 41018 17808
rect 44910 17796 44916 17808
rect 44823 17768 44916 17796
rect 44910 17756 44916 17768
rect 44968 17796 44974 17808
rect 45094 17796 45100 17808
rect 44968 17768 45100 17796
rect 44968 17756 44974 17768
rect 45094 17756 45100 17768
rect 45152 17756 45158 17808
rect 45462 17796 45468 17808
rect 45423 17768 45468 17796
rect 45462 17756 45468 17768
rect 45520 17756 45526 17808
rect 37737 17731 37795 17737
rect 37737 17728 37749 17731
rect 37700 17700 37749 17728
rect 37700 17688 37706 17700
rect 37737 17697 37749 17700
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 38933 17731 38991 17737
rect 38933 17697 38945 17731
rect 38979 17697 38991 17731
rect 39390 17728 39396 17740
rect 39351 17700 39396 17728
rect 38933 17691 38991 17697
rect 39390 17688 39396 17700
rect 39448 17688 39454 17740
rect 43254 17728 43260 17740
rect 43215 17700 43260 17728
rect 43254 17688 43260 17700
rect 43312 17688 43318 17740
rect 22738 17660 22744 17672
rect 20404 17632 22744 17660
rect 20404 17620 20410 17632
rect 22738 17620 22744 17632
rect 22796 17620 22802 17672
rect 26602 17660 26608 17672
rect 26563 17632 26608 17660
rect 26602 17620 26608 17632
rect 26660 17620 26666 17672
rect 29641 17663 29699 17669
rect 29641 17660 29653 17663
rect 26706 17632 29653 17660
rect 22278 17552 22284 17604
rect 22336 17592 22342 17604
rect 26706 17592 26734 17632
rect 29641 17629 29653 17632
rect 29687 17629 29699 17663
rect 29641 17623 29699 17629
rect 34238 17620 34244 17672
rect 34296 17660 34302 17672
rect 35161 17663 35219 17669
rect 35161 17660 35173 17663
rect 34296 17632 35173 17660
rect 34296 17620 34302 17632
rect 35161 17629 35173 17632
rect 35207 17660 35219 17663
rect 35526 17660 35532 17672
rect 35207 17632 35532 17660
rect 35207 17629 35219 17632
rect 35161 17623 35219 17629
rect 35526 17620 35532 17632
rect 35584 17620 35590 17672
rect 40586 17660 40592 17672
rect 40547 17632 40592 17660
rect 40586 17620 40592 17632
rect 40644 17620 40650 17672
rect 44818 17660 44824 17672
rect 44779 17632 44824 17660
rect 44818 17620 44824 17632
rect 44876 17620 44882 17672
rect 31570 17592 31576 17604
rect 22336 17564 26734 17592
rect 31483 17564 31576 17592
rect 22336 17552 22342 17564
rect 31570 17552 31576 17564
rect 31628 17592 31634 17604
rect 32490 17592 32496 17604
rect 31628 17564 32496 17592
rect 31628 17552 31634 17564
rect 32490 17552 32496 17564
rect 32548 17552 32554 17604
rect 17865 17527 17923 17533
rect 17865 17493 17877 17527
rect 17911 17524 17923 17527
rect 18141 17527 18199 17533
rect 18141 17524 18153 17527
rect 17911 17496 18153 17524
rect 17911 17493 17923 17496
rect 17865 17487 17923 17493
rect 18141 17493 18153 17496
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18506 17524 18512 17536
rect 18467 17496 18512 17524
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 18874 17524 18880 17536
rect 18835 17496 18880 17524
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 23290 17524 23296 17536
rect 23251 17496 23296 17524
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 24578 17524 24584 17536
rect 24539 17496 24584 17524
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 25547 17527 25605 17533
rect 25547 17493 25559 17527
rect 25593 17524 25605 17527
rect 25682 17524 25688 17536
rect 25593 17496 25688 17524
rect 25593 17493 25605 17496
rect 25547 17487 25605 17493
rect 25682 17484 25688 17496
rect 25740 17484 25746 17536
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25832 17496 25881 17524
rect 25832 17484 25838 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 25869 17487 25927 17493
rect 28307 17527 28365 17533
rect 28307 17493 28319 17527
rect 28353 17524 28365 17527
rect 29454 17524 29460 17536
rect 28353 17496 29460 17524
rect 28353 17493 28365 17496
rect 28307 17487 28365 17493
rect 29454 17484 29460 17496
rect 29512 17484 29518 17536
rect 30098 17524 30104 17536
rect 30059 17496 30104 17524
rect 30098 17484 30104 17496
rect 30156 17484 30162 17536
rect 30926 17524 30932 17536
rect 30887 17496 30932 17524
rect 30926 17484 30932 17496
rect 30984 17484 30990 17536
rect 31941 17527 31999 17533
rect 31941 17493 31953 17527
rect 31987 17524 31999 17527
rect 32398 17524 32404 17536
rect 31987 17496 32404 17524
rect 31987 17493 31999 17496
rect 31941 17487 31999 17493
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 36538 17524 36544 17536
rect 36499 17496 36544 17524
rect 36538 17484 36544 17496
rect 36596 17484 36602 17536
rect 37918 17524 37924 17536
rect 37879 17496 37924 17524
rect 37918 17484 37924 17496
rect 37976 17484 37982 17536
rect 41509 17527 41567 17533
rect 41509 17493 41521 17527
rect 41555 17524 41567 17527
rect 43254 17524 43260 17536
rect 41555 17496 43260 17524
rect 41555 17493 41567 17496
rect 41509 17487 41567 17493
rect 43254 17484 43260 17496
rect 43312 17484 43318 17536
rect 43487 17527 43545 17533
rect 43487 17493 43499 17527
rect 43533 17524 43545 17527
rect 43622 17524 43628 17536
rect 43533 17496 43628 17524
rect 43533 17493 43545 17496
rect 43487 17487 43545 17493
rect 43622 17484 43628 17496
rect 43680 17484 43686 17536
rect 43806 17524 43812 17536
rect 43767 17496 43812 17524
rect 43806 17484 43812 17496
rect 43864 17484 43870 17536
rect 1104 17434 48852 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 48852 17434
rect 1104 17360 48852 17382
rect 16850 17320 16856 17332
rect 16811 17292 16856 17320
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 17083 17323 17141 17329
rect 17083 17289 17095 17323
rect 17129 17320 17141 17323
rect 18506 17320 18512 17332
rect 17129 17292 18512 17320
rect 17129 17289 17141 17292
rect 17083 17283 17141 17289
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 20346 17320 20352 17332
rect 18656 17292 20352 17320
rect 18656 17280 18662 17292
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 20622 17320 20628 17332
rect 20583 17292 20628 17320
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 22738 17320 22744 17332
rect 22699 17292 22744 17320
rect 22738 17280 22744 17292
rect 22796 17280 22802 17332
rect 23382 17320 23388 17332
rect 23343 17292 23388 17320
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23934 17320 23940 17332
rect 23895 17292 23940 17320
rect 23934 17280 23940 17292
rect 23992 17280 23998 17332
rect 25038 17320 25044 17332
rect 24999 17292 25044 17320
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 26513 17323 26571 17329
rect 26513 17289 26525 17323
rect 26559 17320 26571 17323
rect 26694 17320 26700 17332
rect 26559 17292 26700 17320
rect 26559 17289 26571 17292
rect 26513 17283 26571 17289
rect 26694 17280 26700 17292
rect 26752 17280 26758 17332
rect 28721 17323 28779 17329
rect 28721 17289 28733 17323
rect 28767 17320 28779 17323
rect 29270 17320 29276 17332
rect 28767 17292 29276 17320
rect 28767 17289 28779 17292
rect 28721 17283 28779 17289
rect 29270 17280 29276 17292
rect 29328 17280 29334 17332
rect 30650 17320 30656 17332
rect 30611 17292 30656 17320
rect 30650 17280 30656 17292
rect 30708 17280 30714 17332
rect 31113 17323 31171 17329
rect 31113 17289 31125 17323
rect 31159 17320 31171 17323
rect 31294 17320 31300 17332
rect 31159 17292 31300 17320
rect 31159 17289 31171 17292
rect 31113 17283 31171 17289
rect 31294 17280 31300 17292
rect 31352 17280 31358 17332
rect 31481 17323 31539 17329
rect 31481 17289 31493 17323
rect 31527 17320 31539 17323
rect 32214 17320 32220 17332
rect 31527 17292 32220 17320
rect 31527 17289 31539 17292
rect 31481 17283 31539 17289
rect 32214 17280 32220 17292
rect 32272 17280 32278 17332
rect 34514 17320 34520 17332
rect 34475 17292 34520 17320
rect 34514 17280 34520 17292
rect 34572 17280 34578 17332
rect 36906 17320 36912 17332
rect 34900 17292 36912 17320
rect 17497 17255 17555 17261
rect 17497 17221 17509 17255
rect 17543 17252 17555 17255
rect 17770 17252 17776 17264
rect 17543 17224 17776 17252
rect 17543 17221 17555 17224
rect 17497 17215 17555 17221
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 18690 17252 18696 17264
rect 18651 17224 18696 17252
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 25958 17252 25964 17264
rect 25608 17224 25964 17252
rect 18138 17184 18144 17196
rect 18051 17156 18144 17184
rect 18138 17144 18144 17156
rect 18196 17184 18202 17196
rect 18874 17184 18880 17196
rect 18196 17156 18880 17184
rect 18196 17144 18202 17156
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 20990 17184 20996 17196
rect 20855 17156 20996 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 20990 17144 20996 17156
rect 21048 17184 21054 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21048 17156 22017 17184
rect 21048 17144 21054 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 17012 17119 17070 17125
rect 17012 17085 17024 17119
rect 17058 17116 17070 17119
rect 19613 17119 19671 17125
rect 17058 17088 17908 17116
rect 17058 17085 17070 17088
rect 17012 17079 17070 17085
rect 17880 16989 17908 17088
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 20346 17116 20352 17128
rect 19659 17088 20352 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 22557 17119 22615 17125
rect 22557 17085 22569 17119
rect 22603 17116 22615 17119
rect 22603 17088 23152 17116
rect 22603 17085 22615 17088
rect 22557 17079 22615 17085
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 19245 17051 19303 17057
rect 18288 17020 18333 17048
rect 18288 17008 18294 17020
rect 19245 17017 19257 17051
rect 19291 17048 19303 17051
rect 19518 17048 19524 17060
rect 19291 17020 19524 17048
rect 19291 17017 19303 17020
rect 19245 17011 19303 17017
rect 19518 17008 19524 17020
rect 19576 17048 19582 17060
rect 20070 17048 20076 17060
rect 19576 17020 20076 17048
rect 19576 17008 19582 17020
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 20622 17008 20628 17060
rect 20680 17048 20686 17060
rect 21130 17051 21188 17057
rect 21130 17048 21142 17051
rect 20680 17020 21142 17048
rect 20680 17008 20686 17020
rect 21130 17017 21142 17020
rect 21176 17017 21188 17051
rect 21130 17011 21188 17017
rect 23124 16992 23152 17088
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 25608 17125 25636 17224
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 27706 17212 27712 17264
rect 27764 17252 27770 17264
rect 29730 17252 29736 17264
rect 27764 17224 29736 17252
rect 27764 17212 27770 17224
rect 29730 17212 29736 17224
rect 29788 17252 29794 17264
rect 29917 17255 29975 17261
rect 29917 17252 29929 17255
rect 29788 17224 29929 17252
rect 29788 17212 29794 17224
rect 29917 17221 29929 17224
rect 29963 17221 29975 17255
rect 30668 17252 30696 17280
rect 31662 17252 31668 17264
rect 30668 17224 31668 17252
rect 29917 17215 29975 17221
rect 31662 17212 31668 17224
rect 31720 17252 31726 17264
rect 31757 17255 31815 17261
rect 31757 17252 31769 17255
rect 31720 17224 31769 17252
rect 31720 17212 31726 17224
rect 31757 17221 31769 17224
rect 31803 17252 31815 17255
rect 32033 17255 32091 17261
rect 32033 17252 32045 17255
rect 31803 17224 32045 17252
rect 31803 17221 31815 17224
rect 31757 17215 31815 17221
rect 32033 17221 32045 17224
rect 32079 17221 32091 17255
rect 32033 17215 32091 17221
rect 33689 17255 33747 17261
rect 33689 17221 33701 17255
rect 33735 17252 33747 17255
rect 34146 17252 34152 17264
rect 33735 17224 34152 17252
rect 33735 17221 33747 17224
rect 33689 17215 33747 17221
rect 26602 17144 26608 17196
rect 26660 17184 26666 17196
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 26660 17156 27353 17184
rect 26660 17144 26666 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17184 28411 17187
rect 29178 17184 29184 17196
rect 28399 17156 29184 17184
rect 28399 17153 28411 17156
rect 28353 17147 28411 17153
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 29365 17187 29423 17193
rect 29365 17153 29377 17187
rect 29411 17184 29423 17187
rect 30098 17184 30104 17196
rect 29411 17156 30104 17184
rect 29411 17153 29423 17156
rect 29365 17147 29423 17153
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 32048 17184 32076 17215
rect 34146 17212 34152 17224
rect 34204 17252 34210 17264
rect 34900 17252 34928 17292
rect 36906 17280 36912 17292
rect 36964 17280 36970 17332
rect 37642 17280 37648 17332
rect 37700 17320 37706 17332
rect 37737 17323 37795 17329
rect 37737 17320 37749 17323
rect 37700 17292 37749 17320
rect 37700 17280 37706 17292
rect 37737 17289 37749 17292
rect 37783 17289 37795 17323
rect 38286 17320 38292 17332
rect 38247 17292 38292 17320
rect 37737 17283 37795 17289
rect 38286 17280 38292 17292
rect 38344 17280 38350 17332
rect 38654 17320 38660 17332
rect 38615 17292 38660 17320
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 39390 17280 39396 17332
rect 39448 17320 39454 17332
rect 39853 17323 39911 17329
rect 39853 17320 39865 17323
rect 39448 17292 39865 17320
rect 39448 17280 39454 17292
rect 39853 17289 39865 17292
rect 39899 17289 39911 17323
rect 42610 17320 42616 17332
rect 42571 17292 42616 17320
rect 39853 17283 39911 17289
rect 42610 17280 42616 17292
rect 42668 17280 42674 17332
rect 43254 17320 43260 17332
rect 43215 17292 43260 17320
rect 43254 17280 43260 17292
rect 43312 17280 43318 17332
rect 44818 17280 44824 17332
rect 44876 17320 44882 17332
rect 45143 17323 45201 17329
rect 45143 17320 45155 17323
rect 44876 17292 45155 17320
rect 44876 17280 44882 17292
rect 45143 17289 45155 17292
rect 45189 17289 45201 17323
rect 45143 17283 45201 17289
rect 34204 17224 34928 17252
rect 34204 17212 34210 17224
rect 35434 17212 35440 17264
rect 35492 17252 35498 17264
rect 36354 17252 36360 17264
rect 35492 17224 36360 17252
rect 35492 17212 35498 17224
rect 36354 17212 36360 17224
rect 36412 17212 36418 17264
rect 36538 17252 36544 17264
rect 36499 17224 36544 17252
rect 36538 17212 36544 17224
rect 36596 17212 36602 17264
rect 40586 17252 40592 17264
rect 39592 17224 40592 17252
rect 34057 17187 34115 17193
rect 34057 17184 34069 17187
rect 32048 17156 34069 17184
rect 34057 17153 34069 17156
rect 34103 17184 34115 17187
rect 34606 17184 34612 17196
rect 34103 17156 34612 17184
rect 34103 17153 34115 17156
rect 34057 17147 34115 17153
rect 34606 17144 34612 17156
rect 34664 17184 34670 17196
rect 39592 17193 39620 17224
rect 40586 17212 40592 17224
rect 40644 17212 40650 17264
rect 42981 17255 43039 17261
rect 42981 17221 42993 17255
rect 43027 17252 43039 17255
rect 43162 17252 43168 17264
rect 43027 17224 43168 17252
rect 43027 17221 43039 17224
rect 42981 17215 43039 17221
rect 43162 17212 43168 17224
rect 43220 17212 43226 17264
rect 34977 17187 35035 17193
rect 34977 17184 34989 17187
rect 34664 17156 34989 17184
rect 34664 17144 34670 17156
rect 34977 17153 34989 17156
rect 35023 17153 35035 17187
rect 35897 17187 35955 17193
rect 35897 17184 35909 17187
rect 34977 17147 35035 17153
rect 35065 17156 35909 17184
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23992 17088 24133 17116
rect 23992 17076 23998 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 25608 17119 25686 17125
rect 25608 17088 25640 17119
rect 24121 17079 24179 17085
rect 25628 17085 25640 17088
rect 25674 17085 25686 17119
rect 25628 17079 25686 17085
rect 30929 17119 30987 17125
rect 30929 17085 30941 17119
rect 30975 17116 30987 17119
rect 31570 17116 31576 17128
rect 30975 17088 31576 17116
rect 30975 17085 30987 17088
rect 30929 17079 30987 17085
rect 31570 17076 31576 17088
rect 31628 17076 31634 17128
rect 31941 17119 31999 17125
rect 31941 17085 31953 17119
rect 31987 17116 31999 17119
rect 32030 17116 32036 17128
rect 31987 17088 32036 17116
rect 31987 17085 31999 17088
rect 31941 17079 31999 17085
rect 24765 17051 24823 17057
rect 24765 17017 24777 17051
rect 24811 17048 24823 17051
rect 24946 17048 24952 17060
rect 24811 17020 24952 17048
rect 24811 17017 24823 17020
rect 24765 17011 24823 17017
rect 24946 17008 24952 17020
rect 25004 17048 25010 17060
rect 26142 17048 26148 17060
rect 25004 17020 26148 17048
rect 25004 17008 25010 17020
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 27054 17051 27112 17057
rect 27054 17048 27066 17051
rect 26896 17020 27066 17048
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18414 16980 18420 16992
rect 17911 16952 18420 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19797 16983 19855 16989
rect 19797 16980 19809 16983
rect 19392 16952 19809 16980
rect 19392 16940 19398 16952
rect 19797 16949 19809 16952
rect 19843 16949 19855 16983
rect 19797 16943 19855 16949
rect 21542 16940 21548 16992
rect 21600 16980 21606 16992
rect 21729 16983 21787 16989
rect 21729 16980 21741 16983
rect 21600 16952 21741 16980
rect 21600 16940 21606 16952
rect 21729 16949 21741 16952
rect 21775 16949 21787 16983
rect 23106 16980 23112 16992
rect 23067 16952 23112 16980
rect 21729 16943 21787 16949
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 25498 16980 25504 16992
rect 25459 16952 25504 16980
rect 25498 16940 25504 16952
rect 25556 16940 25562 16992
rect 25731 16983 25789 16989
rect 25731 16949 25743 16983
rect 25777 16980 25789 16983
rect 25866 16980 25872 16992
rect 25777 16952 25872 16980
rect 25777 16949 25789 16952
rect 25731 16943 25789 16949
rect 25866 16940 25872 16952
rect 25924 16940 25930 16992
rect 25958 16940 25964 16992
rect 26016 16980 26022 16992
rect 26053 16983 26111 16989
rect 26053 16980 26065 16983
rect 26016 16952 26065 16980
rect 26016 16940 26022 16952
rect 26053 16949 26065 16952
rect 26099 16949 26111 16983
rect 26786 16980 26792 16992
rect 26747 16952 26792 16980
rect 26053 16943 26111 16949
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 26896 16980 26924 17020
rect 27054 17017 27066 17020
rect 27100 17017 27112 17051
rect 27054 17011 27112 17017
rect 27150 17051 27208 17057
rect 27150 17017 27162 17051
rect 27196 17048 27208 17051
rect 27246 17048 27252 17060
rect 27196 17020 27252 17048
rect 27196 17017 27208 17020
rect 27150 17011 27208 17017
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 29457 17051 29515 17057
rect 29457 17048 29469 17051
rect 29012 17020 29469 17048
rect 29012 16992 29040 17020
rect 29457 17017 29469 17020
rect 29503 17017 29515 17051
rect 29457 17011 29515 17017
rect 30377 17051 30435 17057
rect 30377 17017 30389 17051
rect 30423 17048 30435 17051
rect 30834 17048 30840 17060
rect 30423 17020 30840 17048
rect 30423 17017 30435 17020
rect 30377 17011 30435 17017
rect 30834 17008 30840 17020
rect 30892 17048 30898 17060
rect 31956 17048 31984 17079
rect 32030 17076 32036 17088
rect 32088 17076 32094 17128
rect 32217 17119 32275 17125
rect 32217 17085 32229 17119
rect 32263 17116 32275 17119
rect 32398 17116 32404 17128
rect 32263 17088 32404 17116
rect 32263 17085 32275 17088
rect 32217 17079 32275 17085
rect 32398 17076 32404 17088
rect 32456 17076 32462 17128
rect 33505 17119 33563 17125
rect 33505 17116 33517 17119
rect 33428 17088 33517 17116
rect 30892 17020 31984 17048
rect 30892 17008 30898 17020
rect 33428 16992 33456 17088
rect 33505 17085 33517 17088
rect 33551 17085 33563 17119
rect 33505 17079 33563 17085
rect 34330 17076 34336 17128
rect 34388 17116 34394 17128
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 34388 17088 34897 17116
rect 34388 17076 34394 17088
rect 34885 17085 34897 17088
rect 34931 17116 34943 17119
rect 35065 17116 35093 17156
rect 35897 17153 35909 17156
rect 35943 17153 35955 17187
rect 35897 17147 35955 17153
rect 39577 17187 39635 17193
rect 39577 17153 39589 17187
rect 39623 17153 39635 17187
rect 39577 17147 39635 17153
rect 40678 17144 40684 17196
rect 40736 17184 40742 17196
rect 41690 17184 41696 17196
rect 40736 17156 41696 17184
rect 40736 17144 40742 17156
rect 41690 17144 41696 17156
rect 41748 17144 41754 17196
rect 43180 17184 43208 17212
rect 43809 17187 43867 17193
rect 43809 17184 43821 17187
rect 43180 17156 43821 17184
rect 43809 17153 43821 17156
rect 43855 17153 43867 17187
rect 43809 17147 43867 17153
rect 44821 17187 44879 17193
rect 44821 17153 44833 17187
rect 44867 17184 44879 17187
rect 44910 17184 44916 17196
rect 44867 17156 44916 17184
rect 44867 17153 44879 17156
rect 44821 17147 44879 17153
rect 44910 17144 44916 17156
rect 44968 17144 44974 17196
rect 34931 17088 35093 17116
rect 35161 17119 35219 17125
rect 34931 17085 34943 17088
rect 34885 17079 34943 17085
rect 35161 17085 35173 17119
rect 35207 17116 35219 17119
rect 35526 17116 35532 17128
rect 35207 17088 35532 17116
rect 35207 17085 35219 17088
rect 35161 17079 35219 17085
rect 35526 17076 35532 17088
rect 35584 17076 35590 17128
rect 36354 17076 36360 17128
rect 36412 17116 36418 17128
rect 36449 17119 36507 17125
rect 36449 17116 36461 17119
rect 36412 17088 36461 17116
rect 36412 17076 36418 17088
rect 36449 17085 36461 17088
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 36725 17119 36783 17125
rect 36725 17085 36737 17119
rect 36771 17085 36783 17119
rect 36725 17079 36783 17085
rect 35544 17048 35572 17076
rect 36740 17048 36768 17079
rect 38286 17076 38292 17128
rect 38344 17116 38350 17128
rect 38841 17119 38899 17125
rect 38841 17116 38853 17119
rect 38344 17088 38853 17116
rect 38344 17076 38350 17088
rect 38841 17085 38853 17088
rect 38887 17085 38899 17119
rect 39390 17116 39396 17128
rect 39351 17088 39396 17116
rect 38841 17079 38899 17085
rect 39390 17076 39396 17088
rect 39448 17076 39454 17128
rect 40532 17119 40590 17125
rect 40532 17116 40544 17119
rect 40236 17088 40544 17116
rect 35544 17020 36768 17048
rect 40236 16992 40264 17088
rect 40532 17085 40544 17088
rect 40578 17085 40590 17119
rect 40532 17079 40590 17085
rect 45072 17119 45130 17125
rect 45072 17085 45084 17119
rect 45118 17116 45130 17119
rect 45186 17116 45192 17128
rect 45118 17088 45192 17116
rect 45118 17085 45130 17088
rect 45072 17079 45130 17085
rect 45186 17076 45192 17088
rect 45244 17116 45250 17128
rect 45465 17119 45523 17125
rect 45465 17116 45477 17119
rect 45244 17088 45477 17116
rect 45244 17076 45250 17088
rect 45465 17085 45477 17088
rect 45511 17085 45523 17119
rect 45465 17079 45523 17085
rect 46144 17119 46202 17125
rect 46144 17085 46156 17119
rect 46190 17085 46202 17119
rect 46144 17079 46202 17085
rect 42014 17051 42072 17057
rect 42014 17048 42026 17051
rect 41524 17020 42026 17048
rect 27706 16980 27712 16992
rect 26896 16952 27712 16980
rect 27706 16940 27712 16952
rect 27764 16940 27770 16992
rect 28994 16980 29000 16992
rect 28955 16952 29000 16980
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 32401 16983 32459 16989
rect 32401 16949 32413 16983
rect 32447 16980 32459 16983
rect 32490 16980 32496 16992
rect 32447 16952 32496 16980
rect 32447 16949 32459 16952
rect 32401 16943 32459 16949
rect 32490 16940 32496 16952
rect 32548 16940 32554 16992
rect 32766 16940 32772 16992
rect 32824 16980 32830 16992
rect 32953 16983 33011 16989
rect 32953 16980 32965 16983
rect 32824 16952 32965 16980
rect 32824 16940 32830 16952
rect 32953 16949 32965 16952
rect 32999 16949 33011 16983
rect 33410 16980 33416 16992
rect 33371 16952 33416 16980
rect 32953 16943 33011 16949
rect 33410 16940 33416 16952
rect 33468 16940 33474 16992
rect 34790 16940 34796 16992
rect 34848 16980 34854 16992
rect 35342 16980 35348 16992
rect 34848 16952 35348 16980
rect 34848 16940 34854 16952
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 36354 16940 36360 16992
rect 36412 16980 36418 16992
rect 36909 16983 36967 16989
rect 36909 16980 36921 16983
rect 36412 16952 36921 16980
rect 36412 16940 36418 16952
rect 36909 16949 36921 16952
rect 36955 16949 36967 16983
rect 40218 16980 40224 16992
rect 40179 16952 40224 16980
rect 36909 16943 36967 16949
rect 40218 16940 40224 16952
rect 40276 16940 40282 16992
rect 40310 16940 40316 16992
rect 40368 16980 40374 16992
rect 40635 16983 40693 16989
rect 40635 16980 40647 16983
rect 40368 16952 40647 16980
rect 40368 16940 40374 16952
rect 40635 16949 40647 16952
rect 40681 16949 40693 16983
rect 40954 16980 40960 16992
rect 40915 16952 40960 16980
rect 40635 16943 40693 16949
rect 40954 16940 40960 16952
rect 41012 16980 41018 16992
rect 41524 16989 41552 17020
rect 42014 17017 42026 17020
rect 42060 17017 42072 17051
rect 43530 17048 43536 17060
rect 43491 17020 43536 17048
rect 42014 17011 42072 17017
rect 43530 17008 43536 17020
rect 43588 17008 43594 17060
rect 43625 17051 43683 17057
rect 43625 17017 43637 17051
rect 43671 17017 43683 17051
rect 43625 17011 43683 17017
rect 41509 16983 41567 16989
rect 41509 16980 41521 16983
rect 41012 16952 41521 16980
rect 41012 16940 41018 16952
rect 41509 16949 41521 16952
rect 41555 16949 41567 16983
rect 41509 16943 41567 16949
rect 43254 16940 43260 16992
rect 43312 16980 43318 16992
rect 43640 16980 43668 17011
rect 44634 17008 44640 17060
rect 44692 17048 44698 17060
rect 46159 17048 46187 17079
rect 46569 17051 46627 17057
rect 46569 17048 46581 17051
rect 44692 17020 46581 17048
rect 44692 17008 44698 17020
rect 46569 17017 46581 17020
rect 46615 17017 46627 17051
rect 46569 17011 46627 17017
rect 43312 16952 43668 16980
rect 46247 16983 46305 16989
rect 43312 16940 43318 16952
rect 46247 16949 46259 16983
rect 46293 16980 46305 16983
rect 46382 16980 46388 16992
rect 46293 16952 46388 16980
rect 46293 16949 46305 16952
rect 46247 16943 46305 16949
rect 46382 16940 46388 16952
rect 46440 16940 46446 16992
rect 1104 16890 48852 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 48852 16890
rect 1104 16816 48852 16838
rect 16807 16779 16865 16785
rect 16807 16745 16819 16779
rect 16853 16776 16865 16779
rect 18138 16776 18144 16788
rect 16853 16748 18144 16776
rect 16853 16745 16865 16748
rect 16807 16739 16865 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 19334 16776 19340 16788
rect 18831 16748 19340 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 18598 16708 18604 16720
rect 17972 16680 18604 16708
rect 16736 16643 16794 16649
rect 16736 16609 16748 16643
rect 16782 16640 16794 16643
rect 16942 16640 16948 16652
rect 16782 16612 16948 16640
rect 16782 16609 16794 16612
rect 16736 16603 16794 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17494 16600 17500 16652
rect 17552 16640 17558 16652
rect 17972 16649 18000 16680
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17552 16612 17969 16640
rect 17552 16600 17558 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 18141 16643 18199 16649
rect 18141 16609 18153 16643
rect 18187 16640 18199 16643
rect 18506 16640 18512 16652
rect 18187 16612 18512 16640
rect 18187 16609 18199 16612
rect 18141 16603 18199 16609
rect 18506 16600 18512 16612
rect 18564 16640 18570 16652
rect 18800 16640 18828 16739
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 21174 16776 21180 16788
rect 21135 16748 21180 16776
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 23063 16779 23121 16785
rect 23063 16745 23075 16779
rect 23109 16776 23121 16779
rect 23382 16776 23388 16788
rect 23109 16748 23388 16776
rect 23109 16745 23121 16748
rect 23063 16739 23121 16745
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 26329 16779 26387 16785
rect 26329 16745 26341 16779
rect 26375 16776 26387 16779
rect 26602 16776 26608 16788
rect 26375 16748 26608 16776
rect 26375 16745 26387 16748
rect 26329 16739 26387 16745
rect 26602 16736 26608 16748
rect 26660 16776 26666 16788
rect 27706 16776 27712 16788
rect 26660 16748 27476 16776
rect 27667 16748 27712 16776
rect 26660 16736 26666 16748
rect 19153 16711 19211 16717
rect 19153 16677 19165 16711
rect 19199 16708 19211 16711
rect 19199 16680 19748 16708
rect 19199 16677 19211 16680
rect 19153 16671 19211 16677
rect 19720 16652 19748 16680
rect 19242 16640 19248 16652
rect 18564 16612 18828 16640
rect 19203 16612 19248 16640
rect 18564 16600 18570 16612
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19760 16612 19809 16640
rect 19760 16600 19766 16612
rect 19797 16609 19809 16612
rect 19843 16640 19855 16643
rect 21192 16640 21220 16736
rect 21542 16708 21548 16720
rect 21503 16680 21548 16708
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 24949 16711 25007 16717
rect 24949 16677 24961 16711
rect 24995 16708 25007 16711
rect 26786 16708 26792 16720
rect 24995 16680 26792 16708
rect 24995 16677 25007 16680
rect 24949 16671 25007 16677
rect 26786 16668 26792 16680
rect 26844 16668 26850 16720
rect 26878 16668 26884 16720
rect 26936 16708 26942 16720
rect 27448 16717 27476 16748
rect 27706 16736 27712 16748
rect 27764 16736 27770 16788
rect 34330 16776 34336 16788
rect 34291 16748 34336 16776
rect 34330 16736 34336 16748
rect 34388 16736 34394 16788
rect 35342 16736 35348 16788
rect 35400 16776 35406 16788
rect 36817 16779 36875 16785
rect 36817 16776 36829 16779
rect 35400 16748 36829 16776
rect 35400 16736 35406 16748
rect 36817 16745 36829 16748
rect 36863 16745 36875 16779
rect 36817 16739 36875 16745
rect 36906 16736 36912 16788
rect 36964 16776 36970 16788
rect 37277 16779 37335 16785
rect 37277 16776 37289 16779
rect 36964 16748 37289 16776
rect 36964 16736 36970 16748
rect 37277 16745 37289 16748
rect 37323 16776 37335 16779
rect 37918 16776 37924 16788
rect 37323 16748 37924 16776
rect 37323 16745 37335 16748
rect 37277 16739 37335 16745
rect 37918 16736 37924 16748
rect 37976 16736 37982 16788
rect 39117 16779 39175 16785
rect 39117 16745 39129 16779
rect 39163 16776 39175 16779
rect 39390 16776 39396 16788
rect 39163 16748 39396 16776
rect 39163 16745 39175 16748
rect 39117 16739 39175 16745
rect 39390 16736 39396 16748
rect 39448 16736 39454 16788
rect 40586 16736 40592 16788
rect 40644 16776 40650 16788
rect 40957 16779 41015 16785
rect 40957 16776 40969 16779
rect 40644 16748 40969 16776
rect 40644 16736 40650 16748
rect 40957 16745 40969 16748
rect 41003 16745 41015 16779
rect 41690 16776 41696 16788
rect 41651 16748 41696 16776
rect 40957 16739 41015 16745
rect 41690 16736 41696 16748
rect 41748 16736 41754 16788
rect 43530 16736 43536 16788
rect 43588 16776 43594 16788
rect 44177 16779 44235 16785
rect 44177 16776 44189 16779
rect 43588 16748 44189 16776
rect 43588 16736 43594 16748
rect 44177 16745 44189 16748
rect 44223 16745 44235 16779
rect 44177 16739 44235 16745
rect 44818 16736 44824 16788
rect 44876 16776 44882 16788
rect 45097 16779 45155 16785
rect 45097 16776 45109 16779
rect 44876 16748 45109 16776
rect 44876 16736 44882 16748
rect 45097 16745 45109 16748
rect 45143 16745 45155 16779
rect 45097 16739 45155 16745
rect 27433 16711 27491 16717
rect 26936 16680 26981 16708
rect 26936 16668 26942 16680
rect 27433 16677 27445 16711
rect 27479 16677 27491 16711
rect 27433 16671 27491 16677
rect 29086 16668 29092 16720
rect 29144 16708 29150 16720
rect 29318 16711 29376 16717
rect 29318 16708 29330 16711
rect 29144 16680 29330 16708
rect 29144 16668 29150 16680
rect 29318 16677 29330 16680
rect 29364 16677 29376 16711
rect 29318 16671 29376 16677
rect 35897 16711 35955 16717
rect 35897 16677 35909 16711
rect 35943 16708 35955 16711
rect 36538 16708 36544 16720
rect 35943 16680 36544 16708
rect 35943 16677 35955 16680
rect 35897 16671 35955 16677
rect 36538 16668 36544 16680
rect 36596 16668 36602 16720
rect 38010 16668 38016 16720
rect 38068 16708 38074 16720
rect 38150 16711 38208 16717
rect 38150 16708 38162 16711
rect 38068 16680 38162 16708
rect 38068 16668 38074 16680
rect 38150 16677 38162 16680
rect 38196 16677 38208 16711
rect 39408 16708 39436 16736
rect 40313 16711 40371 16717
rect 39408 16680 40080 16708
rect 38150 16671 38208 16677
rect 22922 16640 22928 16652
rect 19843 16612 21220 16640
rect 22883 16612 22928 16640
rect 19843 16609 19855 16612
rect 19797 16603 19855 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 24578 16640 24584 16652
rect 24539 16612 24584 16640
rect 24578 16600 24584 16612
rect 24636 16600 24642 16652
rect 31021 16643 31079 16649
rect 31021 16609 31033 16643
rect 31067 16640 31079 16643
rect 31110 16640 31116 16652
rect 31067 16612 31116 16640
rect 31067 16609 31079 16612
rect 31021 16603 31079 16609
rect 31110 16600 31116 16612
rect 31168 16600 31174 16652
rect 32214 16600 32220 16652
rect 32272 16640 32278 16652
rect 32401 16643 32459 16649
rect 32401 16640 32413 16643
rect 32272 16612 32413 16640
rect 32272 16600 32278 16612
rect 32401 16609 32413 16612
rect 32447 16609 32459 16643
rect 32401 16603 32459 16609
rect 32677 16643 32735 16649
rect 32677 16609 32689 16643
rect 32723 16640 32735 16643
rect 33502 16640 33508 16652
rect 32723 16612 33508 16640
rect 32723 16609 32735 16612
rect 32677 16603 32735 16609
rect 33502 16600 33508 16612
rect 33560 16600 33566 16652
rect 34146 16640 34152 16652
rect 34107 16612 34152 16640
rect 34146 16600 34152 16612
rect 34204 16600 34210 16652
rect 35802 16640 35808 16652
rect 35763 16612 35808 16640
rect 35802 16600 35808 16612
rect 35860 16600 35866 16652
rect 39574 16640 39580 16652
rect 39535 16612 39580 16640
rect 39574 16600 39580 16612
rect 39632 16600 39638 16652
rect 40052 16649 40080 16680
rect 40313 16677 40325 16711
rect 40359 16708 40371 16711
rect 43806 16708 43812 16720
rect 40359 16680 43812 16708
rect 40359 16677 40371 16680
rect 40313 16671 40371 16677
rect 43806 16668 43812 16680
rect 43864 16668 43870 16720
rect 47302 16708 47308 16720
rect 43916 16680 47308 16708
rect 43916 16652 43944 16680
rect 47302 16668 47308 16680
rect 47360 16668 47366 16720
rect 40037 16643 40095 16649
rect 40037 16609 40049 16643
rect 40083 16609 40095 16643
rect 41138 16640 41144 16652
rect 41196 16649 41202 16652
rect 41196 16643 41234 16649
rect 40037 16603 40095 16609
rect 40420 16612 41144 16640
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 19978 16572 19984 16584
rect 19939 16544 19984 16572
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 21726 16572 21732 16584
rect 21687 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 26789 16575 26847 16581
rect 26789 16541 26801 16575
rect 26835 16572 26847 16575
rect 27062 16572 27068 16584
rect 26835 16544 27068 16572
rect 26835 16541 26847 16544
rect 26789 16535 26847 16541
rect 27062 16532 27068 16544
rect 27120 16532 27126 16584
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28997 16575 29055 16581
rect 28997 16572 29009 16575
rect 28408 16544 29009 16572
rect 28408 16532 28414 16544
rect 28997 16541 29009 16544
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 31662 16532 31668 16584
rect 31720 16572 31726 16584
rect 32493 16575 32551 16581
rect 32493 16572 32505 16575
rect 31720 16544 32505 16572
rect 31720 16532 31726 16544
rect 32493 16541 32505 16544
rect 32539 16541 32551 16575
rect 32493 16535 32551 16541
rect 33137 16575 33195 16581
rect 33137 16541 33149 16575
rect 33183 16572 33195 16575
rect 33410 16572 33416 16584
rect 33183 16544 33416 16572
rect 33183 16541 33195 16544
rect 33137 16535 33195 16541
rect 33410 16532 33416 16544
rect 33468 16572 33474 16584
rect 33686 16572 33692 16584
rect 33468 16544 33692 16572
rect 33468 16532 33474 16544
rect 33686 16532 33692 16544
rect 33744 16532 33750 16584
rect 37826 16572 37832 16584
rect 37787 16544 37832 16572
rect 37826 16532 37832 16544
rect 37884 16532 37890 16584
rect 20346 16504 20352 16516
rect 20259 16476 20352 16504
rect 20346 16464 20352 16476
rect 20404 16504 20410 16516
rect 27890 16504 27896 16516
rect 20404 16476 21220 16504
rect 20404 16464 20410 16476
rect 21192 16436 21220 16476
rect 23446 16476 27896 16504
rect 23446 16436 23474 16476
rect 27890 16464 27896 16476
rect 27948 16464 27954 16516
rect 38749 16507 38807 16513
rect 38749 16473 38761 16507
rect 38795 16504 38807 16507
rect 40420 16504 40448 16612
rect 41138 16600 41144 16612
rect 41222 16609 41234 16643
rect 41196 16603 41234 16609
rect 42220 16643 42278 16649
rect 42220 16609 42232 16643
rect 42266 16640 42278 16643
rect 42426 16640 42432 16652
rect 42266 16612 42432 16640
rect 42266 16609 42278 16612
rect 42220 16603 42278 16609
rect 41196 16600 41202 16603
rect 42426 16600 42432 16612
rect 42484 16600 42490 16652
rect 43438 16649 43444 16652
rect 43416 16643 43444 16649
rect 43416 16640 43428 16643
rect 43351 16612 43428 16640
rect 43416 16609 43428 16612
rect 43496 16640 43502 16652
rect 43898 16640 43904 16652
rect 43496 16612 43904 16640
rect 43416 16603 43444 16609
rect 43438 16600 43444 16603
rect 43496 16600 43502 16612
rect 43898 16600 43904 16612
rect 43956 16600 43962 16652
rect 44634 16640 44640 16652
rect 44595 16612 44640 16640
rect 44634 16600 44640 16612
rect 44692 16600 44698 16652
rect 45554 16600 45560 16652
rect 45612 16640 45618 16652
rect 45741 16643 45799 16649
rect 45741 16640 45753 16643
rect 45612 16612 45753 16640
rect 45612 16600 45618 16612
rect 45741 16609 45753 16612
rect 45787 16609 45799 16643
rect 47210 16640 47216 16652
rect 47171 16612 47216 16640
rect 45741 16603 45799 16609
rect 47210 16600 47216 16612
rect 47268 16600 47274 16652
rect 42334 16532 42340 16584
rect 42392 16572 42398 16584
rect 42392 16544 46203 16572
rect 42392 16532 42398 16544
rect 38795 16476 40448 16504
rect 38795 16473 38807 16476
rect 38749 16467 38807 16473
rect 40586 16464 40592 16516
rect 40644 16504 40650 16516
rect 40681 16507 40739 16513
rect 40681 16504 40693 16507
rect 40644 16476 40693 16504
rect 40644 16464 40650 16476
rect 40681 16473 40693 16476
rect 40727 16504 40739 16507
rect 41279 16507 41337 16513
rect 41279 16504 41291 16507
rect 40727 16476 41291 16504
rect 40727 16473 40739 16476
rect 40681 16467 40739 16473
rect 41279 16473 41291 16476
rect 41325 16473 41337 16507
rect 41279 16467 41337 16473
rect 43901 16507 43959 16513
rect 43901 16473 43913 16507
rect 43947 16504 43959 16507
rect 44266 16504 44272 16516
rect 43947 16476 44272 16504
rect 43947 16473 43959 16476
rect 43901 16467 43959 16473
rect 44266 16464 44272 16476
rect 44324 16464 44330 16516
rect 44821 16507 44879 16513
rect 44821 16473 44833 16507
rect 44867 16504 44879 16507
rect 45554 16504 45560 16516
rect 44867 16476 45560 16504
rect 44867 16473 44879 16476
rect 44821 16467 44879 16473
rect 45554 16464 45560 16476
rect 45612 16464 45618 16516
rect 46175 16504 46203 16544
rect 47397 16507 47455 16513
rect 47397 16504 47409 16507
rect 46175 16476 47409 16504
rect 47397 16473 47409 16476
rect 47443 16473 47455 16507
rect 47397 16467 47455 16473
rect 25222 16436 25228 16448
rect 21192 16408 23474 16436
rect 25183 16408 25228 16436
rect 25222 16396 25228 16408
rect 25280 16396 25286 16448
rect 28258 16436 28264 16448
rect 28219 16408 28264 16436
rect 28258 16396 28264 16408
rect 28316 16396 28322 16448
rect 29917 16439 29975 16445
rect 29917 16405 29929 16439
rect 29963 16436 29975 16439
rect 30374 16436 30380 16448
rect 29963 16408 30380 16436
rect 29963 16405 29975 16408
rect 29917 16399 29975 16405
rect 30374 16396 30380 16408
rect 30432 16396 30438 16448
rect 31202 16436 31208 16448
rect 31163 16408 31208 16436
rect 31202 16396 31208 16408
rect 31260 16396 31266 16448
rect 31570 16436 31576 16448
rect 31531 16408 31576 16436
rect 31570 16396 31576 16408
rect 31628 16396 31634 16448
rect 31941 16439 31999 16445
rect 31941 16405 31953 16439
rect 31987 16436 31999 16439
rect 32030 16436 32036 16448
rect 31987 16408 32036 16436
rect 31987 16405 31999 16408
rect 31941 16399 31999 16405
rect 32030 16396 32036 16408
rect 32088 16436 32094 16448
rect 34514 16436 34520 16448
rect 32088 16408 34520 16436
rect 32088 16396 32094 16408
rect 34514 16396 34520 16408
rect 34572 16396 34578 16448
rect 34977 16439 35035 16445
rect 34977 16405 34989 16439
rect 35023 16436 35035 16439
rect 35526 16436 35532 16448
rect 35023 16408 35532 16436
rect 35023 16405 35035 16408
rect 34977 16399 35035 16405
rect 35526 16396 35532 16408
rect 35584 16436 35590 16448
rect 36449 16439 36507 16445
rect 36449 16436 36461 16439
rect 35584 16408 36461 16436
rect 35584 16396 35590 16408
rect 36449 16405 36461 16408
rect 36495 16405 36507 16439
rect 36449 16399 36507 16405
rect 42150 16396 42156 16448
rect 42208 16436 42214 16448
rect 42291 16439 42349 16445
rect 42291 16436 42303 16439
rect 42208 16408 42303 16436
rect 42208 16396 42214 16408
rect 42291 16405 42303 16408
rect 42337 16405 42349 16439
rect 42291 16399 42349 16405
rect 43487 16439 43545 16445
rect 43487 16405 43499 16439
rect 43533 16436 43545 16439
rect 43714 16436 43720 16448
rect 43533 16408 43720 16436
rect 43533 16405 43545 16408
rect 43487 16399 43545 16405
rect 43714 16396 43720 16408
rect 43772 16396 43778 16448
rect 46109 16439 46167 16445
rect 46109 16405 46121 16439
rect 46155 16436 46167 16439
rect 46290 16436 46296 16448
rect 46155 16408 46296 16436
rect 46155 16405 46167 16408
rect 46109 16399 46167 16405
rect 46290 16396 46296 16408
rect 46348 16396 46354 16448
rect 1104 16346 48852 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 48852 16346
rect 1104 16272 48852 16294
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 19242 16232 19248 16244
rect 17911 16204 19248 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18340 16037 18368 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19702 16232 19708 16244
rect 19663 16204 19708 16232
rect 19702 16192 19708 16204
rect 19760 16192 19766 16244
rect 20349 16235 20407 16241
rect 20349 16201 20361 16235
rect 20395 16232 20407 16235
rect 20622 16232 20628 16244
rect 20395 16204 20628 16232
rect 20395 16201 20407 16204
rect 20349 16195 20407 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 22005 16235 22063 16241
rect 22005 16232 22017 16235
rect 21600 16204 22017 16232
rect 21600 16192 21606 16204
rect 22005 16201 22017 16204
rect 22051 16201 22063 16235
rect 22005 16195 22063 16201
rect 24213 16235 24271 16241
rect 24213 16201 24225 16235
rect 24259 16232 24271 16235
rect 24578 16232 24584 16244
rect 24259 16204 24584 16232
rect 24259 16201 24271 16204
rect 24213 16195 24271 16201
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 25593 16235 25651 16241
rect 25593 16201 25605 16235
rect 25639 16232 25651 16235
rect 25958 16232 25964 16244
rect 25639 16204 25964 16232
rect 25639 16201 25651 16204
rect 25593 16195 25651 16201
rect 25958 16192 25964 16204
rect 26016 16192 26022 16244
rect 26142 16232 26148 16244
rect 26103 16204 26148 16232
rect 26142 16192 26148 16204
rect 26200 16232 26206 16244
rect 26878 16232 26884 16244
rect 26200 16204 26884 16232
rect 26200 16192 26206 16204
rect 26878 16192 26884 16204
rect 26936 16192 26942 16244
rect 30374 16232 30380 16244
rect 30335 16204 30380 16232
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30837 16235 30895 16241
rect 30837 16201 30849 16235
rect 30883 16232 30895 16235
rect 31110 16232 31116 16244
rect 30883 16204 31116 16232
rect 30883 16201 30895 16204
rect 30837 16195 30895 16201
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 31662 16232 31668 16244
rect 31623 16204 31668 16232
rect 31662 16192 31668 16204
rect 31720 16192 31726 16244
rect 34146 16192 34152 16244
rect 34204 16232 34210 16244
rect 34333 16235 34391 16241
rect 34333 16232 34345 16235
rect 34204 16204 34345 16232
rect 34204 16192 34210 16204
rect 34333 16201 34345 16204
rect 34379 16232 34391 16235
rect 35529 16235 35587 16241
rect 35529 16232 35541 16235
rect 34379 16204 35541 16232
rect 34379 16201 34391 16204
rect 34333 16195 34391 16201
rect 35529 16201 35541 16204
rect 35575 16232 35587 16235
rect 35802 16232 35808 16244
rect 35575 16204 35808 16232
rect 35575 16201 35587 16204
rect 35529 16195 35587 16201
rect 35802 16192 35808 16204
rect 35860 16192 35866 16244
rect 35897 16235 35955 16241
rect 35897 16201 35909 16235
rect 35943 16232 35955 16235
rect 36354 16232 36360 16244
rect 35943 16204 36360 16232
rect 35943 16201 35955 16204
rect 35897 16195 35955 16201
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 22462 16164 22468 16176
rect 21140 16136 22468 16164
rect 21140 16124 21146 16136
rect 22462 16124 22468 16136
rect 22520 16164 22526 16176
rect 22922 16164 22928 16176
rect 22520 16136 22928 16164
rect 22520 16124 22526 16136
rect 22922 16124 22928 16136
rect 22980 16164 22986 16176
rect 23293 16167 23351 16173
rect 23293 16164 23305 16167
rect 22980 16136 23305 16164
rect 22980 16124 22986 16136
rect 23293 16133 23305 16136
rect 23339 16133 23351 16167
rect 27709 16167 27767 16173
rect 27709 16164 27721 16167
rect 23293 16127 23351 16133
rect 26804 16136 27721 16164
rect 18598 16096 18604 16108
rect 18559 16068 18604 16096
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20438 16096 20444 16108
rect 20036 16068 20444 16096
rect 20036 16056 20042 16068
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 21729 16099 21787 16105
rect 21729 16096 21741 16099
rect 21508 16068 21741 16096
rect 21508 16056 21514 16068
rect 21729 16065 21741 16068
rect 21775 16096 21787 16099
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 21775 16068 23673 16096
rect 21775 16065 21787 16068
rect 21729 16059 21787 16065
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 25222 16096 25228 16108
rect 24719 16068 25228 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 26804 16105 26832 16136
rect 27709 16133 27721 16136
rect 27755 16133 27767 16167
rect 27709 16127 27767 16133
rect 33413 16167 33471 16173
rect 33413 16133 33425 16167
rect 33459 16164 33471 16167
rect 33597 16167 33655 16173
rect 33597 16164 33609 16167
rect 33459 16136 33609 16164
rect 33459 16133 33471 16136
rect 33413 16127 33471 16133
rect 33597 16133 33609 16136
rect 33643 16164 33655 16167
rect 34238 16164 34244 16176
rect 33643 16136 34244 16164
rect 33643 16133 33655 16136
rect 33597 16127 33655 16133
rect 34238 16124 34244 16136
rect 34296 16124 34302 16176
rect 35161 16167 35219 16173
rect 35161 16133 35173 16167
rect 35207 16164 35219 16167
rect 35250 16164 35256 16176
rect 35207 16136 35256 16164
rect 35207 16133 35219 16136
rect 35161 16127 35219 16133
rect 35250 16124 35256 16136
rect 35308 16124 35314 16176
rect 26789 16099 26847 16105
rect 26789 16096 26801 16099
rect 25740 16068 26801 16096
rect 25740 16056 25746 16068
rect 26789 16065 26801 16068
rect 26835 16065 26847 16099
rect 27062 16096 27068 16108
rect 27023 16068 27068 16096
rect 26789 16059 26847 16065
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 29454 16096 29460 16108
rect 29415 16068 29460 16096
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 29730 16096 29736 16108
rect 29691 16068 29736 16096
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 30098 16056 30104 16108
rect 30156 16096 30162 16108
rect 31067 16099 31125 16105
rect 31067 16096 31079 16099
rect 30156 16068 31079 16096
rect 30156 16056 30162 16068
rect 31067 16065 31079 16068
rect 31113 16065 31125 16099
rect 31067 16059 31125 16065
rect 32861 16099 32919 16105
rect 32861 16065 32873 16099
rect 32907 16096 32919 16099
rect 33318 16096 33324 16108
rect 32907 16068 33324 16096
rect 32907 16065 32919 16068
rect 32861 16059 32919 16065
rect 33318 16056 33324 16068
rect 33376 16096 33382 16108
rect 33870 16096 33876 16108
rect 33376 16068 33876 16096
rect 33376 16056 33382 16068
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18506 16028 18512 16040
rect 18467 16000 18512 16028
rect 18325 15991 18383 15997
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 22462 16028 22468 16040
rect 22423 16000 22468 16028
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 23290 15988 23296 16040
rect 23348 16028 23354 16040
rect 23348 16000 26648 16028
rect 23348 15988 23354 16000
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 20762 15963 20820 15969
rect 20762 15960 20774 15963
rect 20680 15932 20774 15960
rect 20680 15920 20686 15932
rect 20762 15929 20774 15932
rect 20808 15960 20820 15963
rect 24489 15963 24547 15969
rect 24489 15960 24501 15963
rect 20808 15932 24501 15960
rect 20808 15929 20820 15932
rect 20762 15923 20820 15929
rect 24489 15929 24501 15932
rect 24535 15960 24547 15963
rect 24994 15963 25052 15969
rect 24994 15960 25006 15963
rect 24535 15932 25006 15960
rect 24535 15929 24547 15932
rect 24489 15923 24547 15929
rect 24994 15929 25006 15932
rect 25040 15960 25052 15963
rect 26142 15960 26148 15972
rect 25040 15932 26148 15960
rect 25040 15929 25052 15932
rect 24994 15923 25052 15929
rect 26142 15920 26148 15932
rect 26200 15920 26206 15972
rect 26620 15969 26648 16000
rect 30374 15988 30380 16040
rect 30432 16028 30438 16040
rect 30964 16031 31022 16037
rect 30964 16028 30976 16031
rect 30432 16000 30976 16028
rect 30432 15988 30438 16000
rect 30964 15997 30976 16000
rect 31010 15997 31022 16031
rect 32122 16028 32128 16040
rect 32083 16000 32128 16028
rect 30964 15991 31022 15997
rect 32122 15988 32128 16000
rect 32180 15988 32186 16040
rect 32217 16031 32275 16037
rect 32217 15997 32229 16031
rect 32263 15997 32275 16031
rect 32217 15991 32275 15997
rect 26605 15963 26663 15969
rect 26605 15929 26617 15963
rect 26651 15960 26663 15963
rect 26881 15963 26939 15969
rect 26881 15960 26893 15963
rect 26651 15932 26893 15960
rect 26651 15929 26663 15932
rect 26605 15923 26663 15929
rect 26881 15929 26893 15932
rect 26927 15929 26939 15963
rect 29549 15963 29607 15969
rect 29549 15960 29561 15963
rect 26881 15923 26939 15929
rect 28644 15932 29561 15960
rect 28644 15904 28672 15932
rect 29549 15929 29561 15932
rect 29595 15960 29607 15963
rect 32232 15960 32260 15991
rect 32398 15988 32404 16040
rect 32456 16028 32462 16040
rect 33781 16031 33839 16037
rect 32456 16000 32501 16028
rect 32456 15988 32462 16000
rect 33781 15997 33793 16031
rect 33827 16028 33839 16031
rect 34698 16028 34704 16040
rect 33827 16000 34704 16028
rect 33827 15997 33839 16000
rect 33781 15991 33839 15997
rect 34698 15988 34704 16000
rect 34756 15988 34762 16040
rect 34977 16031 35035 16037
rect 34977 15997 34989 16031
rect 35023 16028 35035 16031
rect 35342 16028 35348 16040
rect 35023 16000 35348 16028
rect 35023 15997 35035 16000
rect 34977 15991 35035 15997
rect 35342 15988 35348 16000
rect 35400 16028 35406 16040
rect 35912 16028 35940 16195
rect 36354 16192 36360 16204
rect 36412 16192 36418 16244
rect 38841 16235 38899 16241
rect 38841 16201 38853 16235
rect 38887 16232 38899 16235
rect 40218 16232 40224 16244
rect 38887 16204 40224 16232
rect 38887 16201 38899 16204
rect 38841 16195 38899 16201
rect 40218 16192 40224 16204
rect 40276 16192 40282 16244
rect 41969 16235 42027 16241
rect 41969 16201 41981 16235
rect 42015 16232 42027 16235
rect 42426 16232 42432 16244
rect 42015 16204 42432 16232
rect 42015 16201 42027 16204
rect 41969 16195 42027 16201
rect 42426 16192 42432 16204
rect 42484 16232 42490 16244
rect 43438 16232 43444 16244
rect 42484 16204 42794 16232
rect 43399 16204 43444 16232
rect 42484 16192 42490 16204
rect 39301 16167 39359 16173
rect 39301 16133 39313 16167
rect 39347 16164 39359 16167
rect 39390 16164 39396 16176
rect 39347 16136 39396 16164
rect 39347 16133 39359 16136
rect 39301 16127 39359 16133
rect 39390 16124 39396 16136
rect 39448 16124 39454 16176
rect 39574 16164 39580 16176
rect 39535 16136 39580 16164
rect 39574 16124 39580 16136
rect 39632 16124 39638 16176
rect 42766 16164 42794 16204
rect 43438 16192 43444 16204
rect 43496 16192 43502 16244
rect 44634 16232 44640 16244
rect 44595 16204 44640 16232
rect 44634 16192 44640 16204
rect 44692 16192 44698 16244
rect 45554 16232 45560 16244
rect 45515 16204 45560 16232
rect 45554 16192 45560 16204
rect 45612 16192 45618 16244
rect 47210 16164 47216 16176
rect 42766 16136 47216 16164
rect 47210 16124 47216 16136
rect 47268 16124 47274 16176
rect 40586 16096 40592 16108
rect 40547 16068 40592 16096
rect 40586 16056 40592 16068
rect 40644 16056 40650 16108
rect 40770 16056 40776 16108
rect 40828 16096 40834 16108
rect 40865 16099 40923 16105
rect 40865 16096 40877 16099
rect 40828 16068 40877 16096
rect 40828 16056 40834 16068
rect 40865 16065 40877 16068
rect 40911 16065 40923 16099
rect 40865 16059 40923 16065
rect 35400 16000 35940 16028
rect 36357 16031 36415 16037
rect 35400 15988 35406 16000
rect 36357 15997 36369 16031
rect 36403 15997 36415 16031
rect 36906 16028 36912 16040
rect 36867 16000 36912 16028
rect 36357 15991 36415 15997
rect 29595 15932 30420 15960
rect 29595 15929 29607 15932
rect 29549 15923 29607 15929
rect 30392 15904 30420 15932
rect 32048 15932 32260 15960
rect 33229 15963 33287 15969
rect 32048 15904 32076 15932
rect 33229 15929 33241 15963
rect 33275 15960 33287 15963
rect 33502 15960 33508 15972
rect 33275 15932 33508 15960
rect 33275 15929 33287 15932
rect 33229 15923 33287 15929
rect 33502 15920 33508 15932
rect 33560 15920 33566 15972
rect 36173 15963 36231 15969
rect 36173 15960 36185 15963
rect 33980 15932 36185 15960
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 16942 15892 16948 15904
rect 16807 15864 16948 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 21358 15892 21364 15904
rect 21319 15864 21364 15892
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 22646 15892 22652 15904
rect 22607 15864 22652 15892
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 28626 15892 28632 15904
rect 28587 15864 28632 15892
rect 28626 15852 28632 15864
rect 28684 15852 28690 15904
rect 29086 15892 29092 15904
rect 29047 15864 29092 15892
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 30374 15852 30380 15904
rect 30432 15852 30438 15904
rect 32030 15892 32036 15904
rect 31991 15864 32036 15892
rect 32030 15852 32036 15864
rect 32088 15852 32094 15904
rect 32214 15852 32220 15904
rect 32272 15892 32278 15904
rect 33413 15895 33471 15901
rect 33413 15892 33425 15895
rect 32272 15864 33425 15892
rect 32272 15852 32278 15864
rect 33413 15861 33425 15864
rect 33459 15861 33471 15895
rect 33413 15855 33471 15861
rect 33778 15852 33784 15904
rect 33836 15892 33842 15904
rect 33980 15901 34008 15932
rect 36173 15929 36185 15932
rect 36219 15960 36231 15963
rect 36372 15960 36400 15991
rect 36906 15988 36912 16000
rect 36964 15988 36970 16040
rect 37918 16028 37924 16040
rect 37879 16000 37924 16028
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 41601 16031 41659 16037
rect 41601 15997 41613 16031
rect 41647 16028 41659 16031
rect 42150 16028 42156 16040
rect 41647 16000 42156 16028
rect 41647 15997 41659 16000
rect 41601 15991 41659 15997
rect 42150 15988 42156 16000
rect 42208 15988 42214 16040
rect 44266 16028 44272 16040
rect 44227 16000 44272 16028
rect 44266 15988 44272 16000
rect 44324 15988 44330 16040
rect 45925 16031 45983 16037
rect 45925 15997 45937 16031
rect 45971 16028 45983 16031
rect 46382 16028 46388 16040
rect 45971 16000 46388 16028
rect 45971 15997 45983 16000
rect 45925 15991 45983 15997
rect 46382 15988 46388 16000
rect 46440 15988 46446 16040
rect 36219 15932 36400 15960
rect 37093 15963 37151 15969
rect 36219 15929 36231 15932
rect 36173 15923 36231 15929
rect 37093 15929 37105 15963
rect 37139 15960 37151 15963
rect 37826 15960 37832 15972
rect 37139 15932 37832 15960
rect 37139 15929 37151 15932
rect 37093 15923 37151 15929
rect 37826 15920 37832 15932
rect 37884 15920 37890 15972
rect 38242 15963 38300 15969
rect 38242 15960 38254 15963
rect 38028 15932 38254 15960
rect 38028 15904 38056 15932
rect 38242 15929 38254 15932
rect 38288 15929 38300 15963
rect 38242 15923 38300 15929
rect 40218 15920 40224 15972
rect 40276 15960 40282 15972
rect 40313 15963 40371 15969
rect 40313 15960 40325 15963
rect 40276 15932 40325 15960
rect 40276 15920 40282 15932
rect 40313 15929 40325 15932
rect 40359 15960 40371 15963
rect 40681 15963 40739 15969
rect 40681 15960 40693 15963
rect 40359 15932 40693 15960
rect 40359 15929 40371 15932
rect 40313 15923 40371 15929
rect 40681 15929 40693 15932
rect 40727 15960 40739 15963
rect 42061 15963 42119 15969
rect 42061 15960 42073 15963
rect 40727 15932 42073 15960
rect 40727 15929 40739 15932
rect 40681 15923 40739 15929
rect 42061 15929 42073 15932
rect 42107 15929 42119 15963
rect 42061 15923 42119 15929
rect 43530 15920 43536 15972
rect 43588 15960 43594 15972
rect 43625 15963 43683 15969
rect 43625 15960 43637 15963
rect 43588 15932 43637 15960
rect 43588 15920 43594 15932
rect 43625 15929 43637 15932
rect 43671 15929 43683 15963
rect 46106 15960 46112 15972
rect 46067 15932 46112 15960
rect 43625 15923 43683 15929
rect 46106 15920 46112 15932
rect 46164 15920 46170 15972
rect 33965 15895 34023 15901
rect 33965 15892 33977 15895
rect 33836 15864 33977 15892
rect 33836 15852 33842 15864
rect 33965 15861 33977 15864
rect 34011 15861 34023 15895
rect 34698 15892 34704 15904
rect 34659 15864 34704 15892
rect 33965 15855 34023 15861
rect 34698 15852 34704 15864
rect 34756 15852 34762 15904
rect 37461 15895 37519 15901
rect 37461 15861 37473 15895
rect 37507 15892 37519 15895
rect 37737 15895 37795 15901
rect 37737 15892 37749 15895
rect 37507 15864 37749 15892
rect 37507 15861 37519 15864
rect 37461 15855 37519 15861
rect 37737 15861 37749 15864
rect 37783 15892 37795 15895
rect 38010 15892 38016 15904
rect 37783 15864 38016 15892
rect 37783 15861 37795 15864
rect 37737 15855 37795 15861
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 1104 15802 48852 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 48852 15802
rect 1104 15728 48852 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 26418 15688 26424 15700
rect 20548 15660 21772 15688
rect 17773 15623 17831 15629
rect 17773 15589 17785 15623
rect 17819 15620 17831 15623
rect 19705 15623 19763 15629
rect 17819 15592 18460 15620
rect 17819 15589 17831 15592
rect 17773 15583 17831 15589
rect 18138 15552 18144 15564
rect 18099 15524 18144 15552
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 18432 15561 18460 15592
rect 19705 15589 19717 15623
rect 19751 15620 19763 15623
rect 20548 15620 20576 15660
rect 21744 15632 21772 15660
rect 23446 15660 26424 15688
rect 19751 15592 20576 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 18417 15555 18475 15561
rect 18417 15521 18429 15555
rect 18463 15552 18475 15555
rect 18506 15552 18512 15564
rect 18463 15524 18512 15552
rect 18463 15521 18475 15524
rect 18417 15515 18475 15521
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 19847 15561 19875 15592
rect 20714 15580 20720 15632
rect 20772 15620 20778 15632
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 20772 15592 21189 15620
rect 20772 15580 20778 15592
rect 21177 15589 21189 15592
rect 21223 15620 21235 15623
rect 21358 15620 21364 15632
rect 21223 15592 21364 15620
rect 21223 15589 21235 15592
rect 21177 15583 21235 15589
rect 21358 15580 21364 15592
rect 21416 15580 21422 15632
rect 21726 15620 21732 15632
rect 21687 15592 21732 15620
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 19832 15555 19890 15561
rect 19832 15552 19844 15555
rect 19810 15524 19844 15552
rect 19832 15521 19844 15524
rect 19878 15521 19890 15555
rect 19832 15515 19890 15521
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 22741 15555 22799 15561
rect 22741 15552 22753 15555
rect 22704 15524 22753 15552
rect 22704 15512 22710 15524
rect 22741 15521 22753 15524
rect 22787 15521 22799 15555
rect 22741 15515 22799 15521
rect 23446 15496 23474 15660
rect 26418 15648 26424 15660
rect 26476 15688 26482 15700
rect 26476 15660 26740 15688
rect 26476 15648 26482 15660
rect 24949 15623 25007 15629
rect 24949 15589 24961 15623
rect 24995 15620 25007 15623
rect 25222 15620 25228 15632
rect 24995 15592 25228 15620
rect 24995 15589 25007 15592
rect 24949 15583 25007 15589
rect 25222 15580 25228 15592
rect 25280 15580 25286 15632
rect 25866 15580 25872 15632
rect 25924 15620 25930 15632
rect 26712 15629 26740 15660
rect 28350 15648 28356 15700
rect 28408 15688 28414 15700
rect 28905 15691 28963 15697
rect 28905 15688 28917 15691
rect 28408 15660 28917 15688
rect 28408 15648 28414 15660
rect 28905 15657 28917 15660
rect 28951 15657 28963 15691
rect 28905 15651 28963 15657
rect 29454 15648 29460 15700
rect 29512 15688 29518 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 29512 15660 29837 15688
rect 29512 15648 29518 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 29825 15651 29883 15657
rect 31205 15691 31263 15697
rect 31205 15657 31217 15691
rect 31251 15688 31263 15691
rect 31662 15688 31668 15700
rect 31251 15660 31668 15688
rect 31251 15657 31263 15660
rect 31205 15651 31263 15657
rect 31662 15648 31668 15660
rect 31720 15648 31726 15700
rect 31941 15691 31999 15697
rect 31941 15657 31953 15691
rect 31987 15688 31999 15691
rect 32214 15688 32220 15700
rect 31987 15660 32220 15688
rect 31987 15657 31999 15660
rect 31941 15651 31999 15657
rect 32214 15648 32220 15660
rect 32272 15648 32278 15700
rect 32398 15688 32404 15700
rect 32324 15660 32404 15688
rect 26605 15623 26663 15629
rect 26605 15620 26617 15623
rect 25924 15592 26617 15620
rect 25924 15580 25930 15592
rect 26605 15589 26617 15592
rect 26651 15589 26663 15623
rect 26605 15583 26663 15589
rect 26697 15623 26755 15629
rect 26697 15589 26709 15623
rect 26743 15620 26755 15623
rect 28626 15620 28632 15632
rect 26743 15592 28632 15620
rect 26743 15589 26755 15592
rect 26697 15583 26755 15589
rect 28626 15580 28632 15592
rect 28684 15580 28690 15632
rect 32030 15620 32036 15632
rect 31036 15592 32036 15620
rect 24210 15552 24216 15564
rect 24171 15524 24216 15552
rect 24210 15512 24216 15524
rect 24268 15512 24274 15564
rect 24765 15555 24823 15561
rect 24765 15521 24777 15555
rect 24811 15552 24823 15555
rect 24854 15552 24860 15564
rect 24811 15524 24860 15552
rect 24811 15521 24823 15524
rect 24765 15515 24823 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 29089 15555 29147 15561
rect 29089 15521 29101 15555
rect 29135 15521 29147 15555
rect 29362 15552 29368 15564
rect 29323 15524 29368 15552
rect 29089 15515 29147 15521
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 18966 15484 18972 15496
rect 18647 15456 18972 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18966 15444 18972 15456
rect 19024 15444 19030 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 23382 15484 23388 15496
rect 23295 15456 23388 15484
rect 23382 15444 23388 15456
rect 23440 15456 23474 15496
rect 27062 15484 27068 15496
rect 27023 15456 27068 15484
rect 23440 15444 23446 15456
rect 27062 15444 27068 15456
rect 27120 15484 27126 15496
rect 27525 15487 27583 15493
rect 27525 15484 27537 15487
rect 27120 15456 27537 15484
rect 27120 15444 27126 15456
rect 27525 15453 27537 15456
rect 27571 15453 27583 15487
rect 27525 15447 27583 15453
rect 28718 15444 28724 15496
rect 28776 15484 28782 15496
rect 29104 15484 29132 15515
rect 29362 15512 29368 15524
rect 29420 15512 29426 15564
rect 31036 15561 31064 15592
rect 32030 15580 32036 15592
rect 32088 15620 32094 15632
rect 32125 15623 32183 15629
rect 32125 15620 32137 15623
rect 32088 15592 32137 15620
rect 32088 15580 32094 15592
rect 32125 15589 32137 15592
rect 32171 15589 32183 15623
rect 32125 15583 32183 15589
rect 31021 15555 31079 15561
rect 31021 15521 31033 15555
rect 31067 15521 31079 15555
rect 31570 15552 31576 15564
rect 31483 15524 31576 15552
rect 31021 15515 31079 15521
rect 31570 15512 31576 15524
rect 31628 15552 31634 15564
rect 32324 15552 32352 15660
rect 32398 15648 32404 15660
rect 32456 15688 32462 15700
rect 34330 15688 34336 15700
rect 32456 15660 34336 15688
rect 32456 15648 32462 15660
rect 34330 15648 34336 15660
rect 34388 15648 34394 15700
rect 34422 15648 34428 15700
rect 34480 15688 34486 15700
rect 35434 15688 35440 15700
rect 34480 15660 35440 15688
rect 34480 15648 34486 15660
rect 35434 15648 35440 15660
rect 35492 15648 35498 15700
rect 36906 15688 36912 15700
rect 36867 15660 36912 15688
rect 36906 15648 36912 15660
rect 36964 15648 36970 15700
rect 37553 15691 37611 15697
rect 37553 15657 37565 15691
rect 37599 15688 37611 15691
rect 37826 15688 37832 15700
rect 37599 15660 37832 15688
rect 37599 15657 37611 15660
rect 37553 15651 37611 15657
rect 37826 15648 37832 15660
rect 37884 15648 37890 15700
rect 37918 15648 37924 15700
rect 37976 15688 37982 15700
rect 38013 15691 38071 15697
rect 38013 15688 38025 15691
rect 37976 15660 38025 15688
rect 37976 15648 37982 15660
rect 38013 15657 38025 15660
rect 38059 15688 38071 15691
rect 38749 15691 38807 15697
rect 38749 15688 38761 15691
rect 38059 15660 38761 15688
rect 38059 15657 38071 15660
rect 38013 15651 38071 15657
rect 38749 15657 38761 15660
rect 38795 15657 38807 15691
rect 41138 15688 41144 15700
rect 41099 15660 41144 15688
rect 38749 15651 38807 15657
rect 41138 15648 41144 15660
rect 41196 15648 41202 15700
rect 44266 15648 44272 15700
rect 44324 15688 44330 15700
rect 47489 15691 47547 15697
rect 47489 15688 47501 15691
rect 44324 15660 47501 15688
rect 44324 15648 44330 15660
rect 47489 15657 47501 15660
rect 47535 15657 47547 15691
rect 47489 15651 47547 15657
rect 33502 15580 33508 15632
rect 33560 15620 33566 15632
rect 33689 15623 33747 15629
rect 33689 15620 33701 15623
rect 33560 15592 33701 15620
rect 33560 15580 33566 15592
rect 33689 15589 33701 15592
rect 33735 15620 33747 15623
rect 35526 15620 35532 15632
rect 33735 15592 35532 15620
rect 33735 15589 33747 15592
rect 33689 15583 33747 15589
rect 35526 15580 35532 15592
rect 35584 15580 35590 15632
rect 36924 15620 36952 15648
rect 36924 15592 38240 15620
rect 32766 15552 32772 15564
rect 31628 15524 32352 15552
rect 32727 15524 32772 15552
rect 31628 15512 31634 15524
rect 32766 15512 32772 15524
rect 32824 15512 32830 15564
rect 33873 15555 33931 15561
rect 33873 15521 33885 15555
rect 33919 15552 33931 15555
rect 33962 15552 33968 15564
rect 33919 15524 33968 15552
rect 33919 15521 33931 15524
rect 33873 15515 33931 15521
rect 33962 15512 33968 15524
rect 34020 15512 34026 15564
rect 34330 15512 34336 15564
rect 34388 15552 34394 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 34388 15524 34897 15552
rect 34388 15512 34394 15524
rect 34885 15521 34897 15524
rect 34931 15521 34943 15555
rect 34885 15515 34943 15521
rect 35115 15555 35173 15561
rect 35115 15521 35127 15555
rect 35161 15552 35173 15555
rect 35434 15552 35440 15564
rect 35161 15524 35440 15552
rect 35161 15521 35173 15524
rect 35115 15515 35173 15521
rect 35434 15512 35440 15524
rect 35492 15512 35498 15564
rect 35621 15555 35679 15561
rect 35621 15521 35633 15555
rect 35667 15552 35679 15555
rect 36446 15552 36452 15564
rect 35667 15524 36452 15552
rect 35667 15521 35679 15524
rect 35621 15515 35679 15521
rect 36446 15512 36452 15524
rect 36504 15512 36510 15564
rect 37734 15552 37740 15564
rect 37695 15524 37740 15552
rect 37734 15512 37740 15524
rect 37792 15512 37798 15564
rect 38212 15561 38240 15592
rect 39942 15580 39948 15632
rect 40000 15620 40006 15632
rect 40037 15623 40095 15629
rect 40037 15620 40049 15623
rect 40000 15592 40049 15620
rect 40000 15580 40006 15592
rect 40037 15589 40049 15592
rect 40083 15589 40095 15623
rect 40037 15583 40095 15589
rect 42886 15580 42892 15632
rect 42944 15620 42950 15632
rect 43530 15620 43536 15632
rect 42944 15592 43536 15620
rect 42944 15580 42950 15592
rect 43530 15580 43536 15592
rect 43588 15580 43594 15632
rect 45925 15623 45983 15629
rect 45925 15589 45937 15623
rect 45971 15620 45983 15623
rect 46106 15620 46112 15632
rect 45971 15592 46112 15620
rect 45971 15589 45983 15592
rect 45925 15583 45983 15589
rect 46106 15580 46112 15592
rect 46164 15580 46170 15632
rect 38197 15555 38255 15561
rect 38197 15521 38209 15555
rect 38243 15552 38255 15555
rect 38286 15552 38292 15564
rect 38243 15524 38292 15552
rect 38243 15521 38255 15524
rect 38197 15515 38255 15521
rect 38286 15512 38292 15524
rect 38344 15512 38350 15564
rect 42245 15555 42303 15561
rect 42245 15521 42257 15555
rect 42291 15552 42303 15555
rect 42334 15552 42340 15564
rect 42291 15524 42340 15552
rect 42291 15521 42303 15524
rect 42245 15515 42303 15521
rect 42334 15512 42340 15524
rect 42392 15512 42398 15564
rect 47302 15552 47308 15564
rect 47263 15524 47308 15552
rect 47302 15512 47308 15524
rect 47360 15512 47366 15564
rect 29178 15484 29184 15496
rect 28776 15456 29184 15484
rect 28776 15444 28782 15456
rect 29178 15444 29184 15456
rect 29236 15484 29242 15496
rect 33778 15484 33784 15496
rect 29236 15456 33784 15484
rect 29236 15444 29242 15456
rect 33778 15444 33784 15456
rect 33836 15444 33842 15496
rect 34238 15444 34244 15496
rect 34296 15484 34302 15496
rect 35253 15487 35311 15493
rect 35253 15484 35265 15487
rect 34296 15456 35265 15484
rect 34296 15444 34302 15456
rect 35253 15453 35265 15456
rect 35299 15484 35311 15487
rect 36538 15484 36544 15496
rect 35299 15456 36544 15484
rect 35299 15453 35311 15456
rect 35253 15447 35311 15453
rect 36538 15444 36544 15456
rect 36596 15444 36602 15496
rect 39574 15444 39580 15496
rect 39632 15484 39638 15496
rect 39945 15487 40003 15493
rect 39945 15484 39957 15487
rect 39632 15456 39957 15484
rect 39632 15444 39638 15456
rect 39945 15453 39957 15456
rect 39991 15484 40003 15487
rect 40310 15484 40316 15496
rect 39991 15456 40316 15484
rect 39991 15453 40003 15456
rect 39945 15447 40003 15453
rect 40310 15444 40316 15456
rect 40368 15444 40374 15496
rect 40589 15487 40647 15493
rect 40589 15453 40601 15487
rect 40635 15484 40647 15487
rect 40862 15484 40868 15496
rect 40635 15456 40868 15484
rect 40635 15453 40647 15456
rect 40589 15447 40647 15453
rect 40862 15444 40868 15456
rect 40920 15444 40926 15496
rect 43438 15484 43444 15496
rect 43399 15456 43444 15484
rect 43438 15444 43444 15456
rect 43496 15444 43502 15496
rect 45830 15484 45836 15496
rect 45791 15456 45836 15484
rect 45830 15444 45836 15456
rect 45888 15444 45894 15496
rect 46474 15484 46480 15496
rect 46435 15456 46480 15484
rect 46474 15444 46480 15456
rect 46532 15444 46538 15496
rect 19935 15419 19993 15425
rect 19935 15385 19947 15419
rect 19981 15416 19993 15419
rect 21818 15416 21824 15428
rect 19981 15388 21824 15416
rect 19981 15385 19993 15388
rect 19935 15379 19993 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 33134 15376 33140 15428
rect 33192 15416 33198 15428
rect 34057 15419 34115 15425
rect 34057 15416 34069 15419
rect 33192 15388 34069 15416
rect 33192 15376 33198 15388
rect 34057 15385 34069 15388
rect 34103 15385 34115 15419
rect 34057 15379 34115 15385
rect 34514 15376 34520 15428
rect 34572 15416 34578 15428
rect 34701 15419 34759 15425
rect 34701 15416 34713 15419
rect 34572 15388 34713 15416
rect 34572 15376 34578 15388
rect 34701 15385 34713 15388
rect 34747 15385 34759 15419
rect 34701 15379 34759 15385
rect 35050 15419 35108 15425
rect 35050 15385 35062 15419
rect 35096 15416 35108 15419
rect 38470 15416 38476 15428
rect 35096 15388 38476 15416
rect 35096 15385 35108 15388
rect 35050 15379 35108 15385
rect 35268 15360 35296 15388
rect 38470 15376 38476 15388
rect 38528 15376 38534 15428
rect 43990 15416 43996 15428
rect 43951 15388 43996 15416
rect 43990 15376 43996 15388
rect 44048 15376 44054 15428
rect 23750 15348 23756 15360
rect 23711 15320 23756 15348
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 25222 15348 25228 15360
rect 25183 15320 25228 15348
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 33226 15348 33232 15360
rect 33187 15320 33232 15348
rect 33226 15308 33232 15320
rect 33284 15308 33290 15360
rect 34330 15348 34336 15360
rect 34291 15320 34336 15348
rect 34330 15308 34336 15320
rect 34388 15308 34394 15360
rect 35250 15308 35256 15360
rect 35308 15308 35314 15360
rect 36633 15351 36691 15357
rect 36633 15317 36645 15351
rect 36679 15348 36691 15351
rect 36814 15348 36820 15360
rect 36679 15320 36820 15348
rect 36679 15317 36691 15320
rect 36633 15311 36691 15317
rect 36814 15308 36820 15320
rect 36872 15308 36878 15360
rect 42061 15351 42119 15357
rect 42061 15317 42073 15351
rect 42107 15348 42119 15351
rect 42242 15348 42248 15360
rect 42107 15320 42248 15348
rect 42107 15317 42119 15320
rect 42061 15311 42119 15317
rect 42242 15308 42248 15320
rect 42300 15308 42306 15360
rect 46198 15308 46204 15360
rect 46256 15348 46262 15360
rect 46753 15351 46811 15357
rect 46753 15348 46765 15351
rect 46256 15320 46765 15348
rect 46256 15308 46262 15320
rect 46753 15317 46765 15320
rect 46799 15317 46811 15351
rect 46753 15311 46811 15317
rect 1104 15258 48852 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 48852 15258
rect 1104 15184 48852 15206
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18196 15116 18245 15144
rect 18196 15104 18202 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 18506 15104 18512 15156
rect 18564 15144 18570 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 18564 15116 18613 15144
rect 18564 15104 18570 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 18601 15107 18659 15113
rect 19015 15147 19073 15153
rect 19015 15113 19027 15147
rect 19061 15144 19073 15147
rect 21082 15144 21088 15156
rect 19061 15116 21088 15144
rect 19061 15113 19073 15116
rect 19015 15107 19073 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 22741 15147 22799 15153
rect 22741 15144 22753 15147
rect 22704 15116 22753 15144
rect 22704 15104 22710 15116
rect 22741 15113 22753 15116
rect 22787 15113 22799 15147
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 22741 15107 22799 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 25866 15144 25872 15156
rect 25827 15116 25872 15144
rect 25866 15104 25872 15116
rect 25924 15104 25930 15156
rect 26142 15144 26148 15156
rect 26103 15116 26148 15144
rect 26142 15104 26148 15116
rect 26200 15104 26206 15156
rect 28258 15104 28264 15156
rect 28316 15144 28322 15156
rect 30193 15147 30251 15153
rect 30193 15144 30205 15147
rect 28316 15116 30205 15144
rect 28316 15104 28322 15116
rect 30193 15113 30205 15116
rect 30239 15113 30251 15147
rect 30193 15107 30251 15113
rect 31573 15147 31631 15153
rect 31573 15113 31585 15147
rect 31619 15144 31631 15147
rect 32030 15144 32036 15156
rect 31619 15116 32036 15144
rect 31619 15113 31631 15116
rect 31573 15107 31631 15113
rect 32030 15104 32036 15116
rect 32088 15104 32094 15156
rect 33394 15147 33452 15153
rect 33394 15113 33406 15147
rect 33440 15144 33452 15147
rect 33778 15144 33784 15156
rect 33440 15116 33784 15144
rect 33440 15113 33452 15116
rect 33394 15107 33452 15113
rect 33778 15104 33784 15116
rect 33836 15144 33842 15156
rect 34238 15144 34244 15156
rect 33836 15116 34244 15144
rect 33836 15104 33842 15116
rect 34238 15104 34244 15116
rect 34296 15104 34302 15156
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 34609 15147 34667 15153
rect 34609 15144 34621 15147
rect 34480 15116 34621 15144
rect 34480 15104 34486 15116
rect 34609 15113 34621 15116
rect 34655 15113 34667 15147
rect 34609 15107 34667 15113
rect 35161 15147 35219 15153
rect 35161 15113 35173 15147
rect 35207 15144 35219 15147
rect 35526 15144 35532 15156
rect 35207 15116 35532 15144
rect 35207 15113 35219 15116
rect 35161 15107 35219 15113
rect 35526 15104 35532 15116
rect 35584 15104 35590 15156
rect 36538 15104 36544 15156
rect 36596 15144 36602 15156
rect 36633 15147 36691 15153
rect 36633 15144 36645 15147
rect 36596 15116 36645 15144
rect 36596 15104 36602 15116
rect 36633 15113 36645 15116
rect 36679 15113 36691 15147
rect 38286 15144 38292 15156
rect 38247 15116 38292 15144
rect 36633 15107 36691 15113
rect 38286 15104 38292 15116
rect 38344 15104 38350 15156
rect 39574 15144 39580 15156
rect 39535 15116 39580 15144
rect 39574 15104 39580 15116
rect 39632 15104 39638 15156
rect 40218 15144 40224 15156
rect 40179 15116 40224 15144
rect 40218 15104 40224 15116
rect 40276 15104 40282 15156
rect 41693 15147 41751 15153
rect 41693 15113 41705 15147
rect 41739 15144 41751 15147
rect 42334 15144 42340 15156
rect 41739 15116 42340 15144
rect 41739 15113 41751 15116
rect 41693 15107 41751 15113
rect 42334 15104 42340 15116
rect 42392 15104 42398 15156
rect 42886 15144 42892 15156
rect 42847 15116 42892 15144
rect 42886 15104 42892 15116
rect 42944 15104 42950 15156
rect 45833 15147 45891 15153
rect 45833 15113 45845 15147
rect 45879 15144 45891 15147
rect 46106 15144 46112 15156
rect 45879 15116 46112 15144
rect 45879 15113 45891 15116
rect 45833 15107 45891 15113
rect 46106 15104 46112 15116
rect 46164 15104 46170 15156
rect 47302 15144 47308 15156
rect 47263 15116 47308 15144
rect 47302 15104 47308 15116
rect 47360 15104 47366 15156
rect 19150 15036 19156 15088
rect 19208 15076 19214 15088
rect 19208 15048 19748 15076
rect 19208 15036 19214 15048
rect 18944 14943 19002 14949
rect 18944 14909 18956 14943
rect 18990 14940 19002 14943
rect 19058 14940 19064 14952
rect 18990 14912 19064 14940
rect 18990 14909 19002 14912
rect 18944 14903 19002 14909
rect 19058 14900 19064 14912
rect 19116 14940 19122 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 19116 14912 19349 14940
rect 19116 14900 19122 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19720 14940 19748 15048
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 24210 15076 24216 15088
rect 23532 15048 24216 15076
rect 23532 15036 23538 15048
rect 24210 15036 24216 15048
rect 24268 15076 24274 15088
rect 24673 15079 24731 15085
rect 24673 15076 24685 15079
rect 24268 15048 24685 15076
rect 24268 15036 24274 15048
rect 24673 15045 24685 15048
rect 24719 15045 24731 15079
rect 25363 15079 25421 15085
rect 25363 15076 25375 15079
rect 24673 15039 24731 15045
rect 24958 15048 25375 15076
rect 19886 15008 19892 15020
rect 19847 14980 19892 15008
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 22002 15008 22008 15020
rect 21315 14980 22008 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 22002 14968 22008 14980
rect 22060 15008 22066 15020
rect 23750 15008 23756 15020
rect 22060 14980 22232 15008
rect 23663 14980 23756 15008
rect 22060 14968 22066 14980
rect 21637 14943 21695 14949
rect 19720 14912 19840 14940
rect 19337 14903 19395 14909
rect 17586 14804 17592 14816
rect 17547 14776 17592 14804
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 19812 14813 19840 14912
rect 21637 14909 21649 14943
rect 21683 14940 21695 14943
rect 21910 14940 21916 14952
rect 21683 14912 21916 14940
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22204 14949 22232 14980
rect 23750 14968 23756 14980
rect 23808 15008 23814 15020
rect 24958 15008 24986 15048
rect 25363 15045 25375 15048
rect 25409 15045 25421 15079
rect 25363 15039 25421 15045
rect 25498 15036 25504 15088
rect 25556 15076 25562 15088
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 25556 15048 27261 15076
rect 25556 15036 25562 15048
rect 27249 15045 27261 15048
rect 27295 15045 27307 15079
rect 28718 15076 28724 15088
rect 28679 15048 28724 15076
rect 27249 15039 27307 15045
rect 28718 15036 28724 15048
rect 28776 15036 28782 15088
rect 29086 15076 29092 15088
rect 28999 15048 29092 15076
rect 29086 15036 29092 15048
rect 29144 15076 29150 15088
rect 29454 15076 29460 15088
rect 29144 15048 29460 15076
rect 29144 15036 29150 15048
rect 29454 15036 29460 15048
rect 29512 15036 29518 15088
rect 33502 15076 33508 15088
rect 33463 15048 33508 15076
rect 33502 15036 33508 15048
rect 33560 15036 33566 15088
rect 34514 15036 34520 15088
rect 34572 15076 34578 15088
rect 34974 15076 34980 15088
rect 34572 15048 34980 15076
rect 34572 15036 34578 15048
rect 34974 15036 34980 15048
rect 35032 15085 35038 15088
rect 35032 15079 35081 15085
rect 35032 15045 35035 15079
rect 35069 15045 35081 15079
rect 35032 15039 35081 15045
rect 35032 15036 35038 15039
rect 38102 15036 38108 15088
rect 38160 15076 38166 15088
rect 38657 15079 38715 15085
rect 38657 15076 38669 15079
rect 38160 15048 38669 15076
rect 38160 15036 38166 15048
rect 38657 15045 38669 15048
rect 38703 15045 38715 15079
rect 38657 15039 38715 15045
rect 39025 15079 39083 15085
rect 39025 15045 39037 15079
rect 39071 15076 39083 15079
rect 40034 15076 40040 15088
rect 39071 15048 40040 15076
rect 39071 15045 39083 15048
rect 39025 15039 39083 15045
rect 28077 15011 28135 15017
rect 28077 15008 28089 15011
rect 23808 14980 24986 15008
rect 26068 14980 28089 15008
rect 23808 14968 23814 14980
rect 22189 14943 22247 14949
rect 22189 14909 22201 14943
rect 22235 14909 22247 14943
rect 22189 14903 22247 14909
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 25222 14940 25228 14952
rect 25280 14949 25286 14952
rect 25280 14943 25318 14949
rect 24820 14912 25228 14940
rect 24820 14900 24826 14912
rect 25222 14900 25228 14912
rect 25306 14909 25318 14943
rect 25280 14903 25318 14909
rect 25280 14900 25286 14903
rect 20251 14875 20309 14881
rect 20251 14841 20263 14875
rect 20297 14872 20309 14875
rect 20622 14872 20628 14884
rect 20297 14844 20628 14872
rect 20297 14841 20309 14844
rect 20251 14835 20309 14841
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 20272 14804 20300 14835
rect 20622 14832 20628 14844
rect 20680 14832 20686 14884
rect 23382 14832 23388 14884
rect 23440 14872 23446 14884
rect 23845 14875 23903 14881
rect 23440 14844 23520 14872
rect 23440 14832 23446 14844
rect 20806 14804 20812 14816
rect 19843 14776 20300 14804
rect 20767 14776 20812 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 23492 14804 23520 14844
rect 23845 14841 23857 14875
rect 23891 14841 23903 14875
rect 24394 14872 24400 14884
rect 24355 14844 24400 14872
rect 23845 14835 23903 14841
rect 23860 14804 23888 14835
rect 24394 14832 24400 14844
rect 24452 14832 24458 14884
rect 24578 14832 24584 14884
rect 24636 14872 24642 14884
rect 24854 14872 24860 14884
rect 24636 14844 24860 14872
rect 24636 14832 24642 14844
rect 24854 14832 24860 14844
rect 24912 14872 24918 14884
rect 25133 14875 25191 14881
rect 25133 14872 25145 14875
rect 24912 14844 25145 14872
rect 24912 14832 24918 14844
rect 25133 14841 25145 14844
rect 25179 14872 25191 14875
rect 26068 14872 26096 14980
rect 28077 14977 28089 14980
rect 28123 15008 28135 15011
rect 29362 15008 29368 15020
rect 28123 14980 29368 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 29362 14968 29368 14980
rect 29420 14968 29426 15020
rect 33226 15008 33232 15020
rect 32232 14980 33232 15008
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14940 26387 14943
rect 26510 14940 26516 14952
rect 26375 14912 26516 14940
rect 26375 14909 26387 14912
rect 26329 14903 26387 14909
rect 26510 14900 26516 14912
rect 26568 14940 26574 14952
rect 27525 14943 27583 14949
rect 27525 14940 27537 14943
rect 26568 14912 27537 14940
rect 26568 14900 26574 14912
rect 27525 14909 27537 14912
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 28169 14943 28227 14949
rect 28169 14909 28181 14943
rect 28215 14940 28227 14943
rect 28258 14940 28264 14952
rect 28215 14912 28264 14940
rect 28215 14909 28227 14912
rect 28169 14903 28227 14909
rect 28258 14900 28264 14912
rect 28316 14900 28322 14952
rect 29270 14940 29276 14952
rect 29231 14912 29276 14940
rect 29270 14900 29276 14912
rect 29328 14900 29334 14952
rect 30929 14943 30987 14949
rect 30929 14909 30941 14943
rect 30975 14940 30987 14943
rect 31088 14943 31146 14949
rect 31088 14940 31100 14943
rect 30975 14912 31100 14940
rect 30975 14909 30987 14912
rect 30929 14903 30987 14909
rect 31088 14909 31100 14912
rect 31134 14940 31146 14943
rect 31478 14940 31484 14952
rect 31134 14912 31484 14940
rect 31134 14909 31146 14912
rect 31088 14903 31146 14909
rect 31478 14900 31484 14912
rect 31536 14900 31542 14952
rect 32232 14949 32260 14980
rect 33226 14968 33232 14980
rect 33284 15008 33290 15020
rect 33597 15011 33655 15017
rect 33597 15008 33609 15011
rect 33284 14980 33609 15008
rect 33284 14968 33290 14980
rect 33597 14977 33609 14980
rect 33643 15008 33655 15011
rect 35250 15008 35256 15020
rect 33643 14980 35256 15008
rect 33643 14977 33655 14980
rect 33597 14971 33655 14977
rect 35250 14968 35256 14980
rect 35308 15008 35314 15020
rect 35897 15011 35955 15017
rect 35897 15008 35909 15011
rect 35308 14980 35909 15008
rect 35308 14968 35314 14980
rect 35897 14977 35909 14980
rect 35943 14977 35955 15011
rect 35897 14971 35955 14977
rect 32125 14943 32183 14949
rect 32125 14909 32137 14943
rect 32171 14940 32183 14943
rect 32217 14943 32275 14949
rect 32217 14940 32229 14943
rect 32171 14912 32229 14940
rect 32171 14909 32183 14912
rect 32125 14903 32183 14909
rect 32217 14909 32229 14912
rect 32263 14909 32275 14943
rect 32766 14940 32772 14952
rect 32679 14912 32772 14940
rect 32217 14903 32275 14909
rect 32766 14900 32772 14912
rect 32824 14940 32830 14952
rect 33137 14943 33195 14949
rect 33137 14940 33149 14943
rect 32824 14912 33149 14940
rect 32824 14900 32830 14912
rect 33137 14909 33149 14912
rect 33183 14940 33195 14943
rect 34422 14940 34428 14952
rect 33183 14912 34428 14940
rect 33183 14909 33195 14912
rect 33137 14903 33195 14909
rect 25179 14844 26096 14872
rect 25179 14841 25191 14844
rect 25133 14835 25191 14841
rect 26142 14832 26148 14884
rect 26200 14872 26206 14884
rect 26650 14875 26708 14881
rect 26650 14872 26662 14875
rect 26200 14844 26662 14872
rect 26200 14832 26206 14844
rect 26650 14841 26662 14844
rect 26696 14841 26708 14875
rect 26650 14835 26708 14841
rect 29454 14832 29460 14884
rect 29512 14872 29518 14884
rect 33244 14881 33272 14912
rect 34422 14900 34428 14912
rect 34480 14900 34486 14952
rect 34606 14900 34612 14952
rect 34664 14940 34670 14952
rect 34885 14943 34943 14949
rect 34885 14940 34897 14943
rect 34664 14912 34897 14940
rect 34664 14900 34670 14912
rect 34885 14909 34897 14912
rect 34931 14940 34943 14943
rect 35434 14940 35440 14952
rect 34931 14912 35440 14940
rect 34931 14909 34943 14912
rect 34885 14903 34943 14909
rect 35434 14900 35440 14912
rect 35492 14940 35498 14952
rect 36265 14943 36323 14949
rect 36265 14940 36277 14943
rect 35492 14912 36277 14940
rect 35492 14900 35498 14912
rect 36265 14909 36277 14912
rect 36311 14909 36323 14943
rect 36906 14940 36912 14952
rect 36867 14912 36912 14940
rect 36265 14903 36323 14909
rect 36906 14900 36912 14912
rect 36964 14900 36970 14952
rect 37274 14900 37280 14952
rect 37332 14940 37338 14952
rect 37461 14943 37519 14949
rect 37461 14940 37473 14943
rect 37332 14912 37473 14940
rect 37332 14900 37338 14912
rect 37461 14909 37473 14912
rect 37507 14940 37519 14943
rect 38286 14940 38292 14952
rect 37507 14912 38292 14940
rect 37507 14909 37519 14912
rect 37461 14903 37519 14909
rect 38286 14900 38292 14912
rect 38344 14900 38350 14952
rect 38470 14940 38476 14952
rect 38383 14912 38476 14940
rect 38470 14900 38476 14912
rect 38528 14940 38534 14952
rect 39040 14940 39068 15039
rect 40034 15036 40040 15048
rect 40092 15036 40098 15088
rect 42199 15079 42257 15085
rect 42199 15076 42211 15079
rect 40604 15048 42211 15076
rect 40604 15020 40632 15048
rect 42199 15045 42211 15048
rect 42245 15045 42257 15079
rect 42199 15039 42257 15045
rect 43257 15079 43315 15085
rect 43257 15045 43269 15079
rect 43303 15076 43315 15079
rect 43530 15076 43536 15088
rect 43303 15048 43536 15076
rect 43303 15045 43315 15048
rect 43257 15039 43315 15045
rect 43530 15036 43536 15048
rect 43588 15036 43594 15088
rect 43990 15076 43996 15088
rect 43951 15048 43996 15076
rect 43990 15036 43996 15048
rect 44048 15036 44054 15088
rect 44913 15079 44971 15085
rect 44913 15045 44925 15079
rect 44959 15076 44971 15079
rect 44959 15048 46520 15076
rect 44959 15045 44971 15048
rect 44913 15039 44971 15045
rect 40586 15008 40592 15020
rect 40499 14980 40592 15008
rect 40586 14968 40592 14980
rect 40644 14968 40650 15020
rect 40862 15008 40868 15020
rect 40823 14980 40868 15008
rect 40862 14968 40868 14980
rect 40920 15008 40926 15020
rect 43441 15011 43499 15017
rect 43441 15008 43453 15011
rect 40920 14980 43453 15008
rect 40920 14968 40926 14980
rect 43441 14977 43453 14980
rect 43487 15008 43499 15011
rect 44361 15011 44419 15017
rect 44361 15008 44373 15011
rect 43487 14980 44373 15008
rect 43487 14977 43499 14980
rect 43441 14971 43499 14977
rect 44361 14977 44373 14980
rect 44407 14977 44419 15011
rect 44361 14971 44419 14977
rect 38528 14912 39068 14940
rect 38528 14900 38534 14912
rect 41966 14900 41972 14952
rect 42024 14940 42030 14952
rect 42096 14943 42154 14949
rect 42096 14940 42108 14943
rect 42024 14912 42108 14940
rect 42024 14900 42030 14912
rect 42096 14909 42108 14912
rect 42142 14909 42154 14943
rect 42096 14903 42154 14909
rect 45056 14943 45114 14949
rect 45056 14909 45068 14943
rect 45102 14940 45114 14943
rect 45296 14940 45324 15048
rect 46492 15020 46520 15048
rect 46198 15008 46204 15020
rect 46159 14980 46204 15008
rect 46198 14968 46204 14980
rect 46256 14968 46262 15020
rect 46474 15008 46480 15020
rect 46435 14980 46480 15008
rect 46474 14968 46480 14980
rect 46532 14968 46538 15020
rect 45102 14912 45324 14940
rect 45102 14909 45114 14912
rect 45056 14903 45114 14909
rect 29594 14875 29652 14881
rect 29594 14872 29606 14875
rect 29512 14844 29606 14872
rect 29512 14832 29518 14844
rect 29594 14841 29606 14844
rect 29640 14841 29652 14875
rect 33229 14875 33287 14881
rect 33229 14872 33241 14875
rect 33207 14844 33241 14872
rect 29594 14835 29652 14841
rect 33229 14841 33241 14844
rect 33275 14841 33287 14875
rect 33962 14872 33968 14884
rect 33923 14844 33968 14872
rect 33229 14835 33287 14841
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 34333 14875 34391 14881
rect 34333 14841 34345 14875
rect 34379 14872 34391 14875
rect 35158 14872 35164 14884
rect 34379 14844 35164 14872
rect 34379 14841 34391 14844
rect 34333 14835 34391 14841
rect 35158 14832 35164 14844
rect 35216 14832 35222 14884
rect 35618 14872 35624 14884
rect 35579 14844 35624 14872
rect 35618 14832 35624 14844
rect 35676 14832 35682 14884
rect 37645 14875 37703 14881
rect 37645 14841 37657 14875
rect 37691 14872 37703 14875
rect 37826 14872 37832 14884
rect 37691 14844 37832 14872
rect 37691 14841 37703 14844
rect 37645 14835 37703 14841
rect 37826 14832 37832 14844
rect 37884 14832 37890 14884
rect 40218 14832 40224 14884
rect 40276 14872 40282 14884
rect 40681 14875 40739 14881
rect 40681 14872 40693 14875
rect 40276 14844 40693 14872
rect 40276 14832 40282 14844
rect 40681 14841 40693 14844
rect 40727 14872 40739 14875
rect 41690 14872 41696 14884
rect 40727 14844 41696 14872
rect 40727 14841 40739 14844
rect 40681 14835 40739 14841
rect 41690 14832 41696 14844
rect 41748 14832 41754 14884
rect 42242 14872 42248 14884
rect 41800 14844 42248 14872
rect 23492 14776 23888 14804
rect 28307 14807 28365 14813
rect 28307 14773 28319 14807
rect 28353 14804 28365 14807
rect 28534 14804 28540 14816
rect 28353 14776 28540 14804
rect 28353 14773 28365 14776
rect 28307 14767 28365 14773
rect 28534 14764 28540 14776
rect 28592 14764 28598 14816
rect 30282 14764 30288 14816
rect 30340 14804 30346 14816
rect 31159 14807 31217 14813
rect 31159 14804 31171 14807
rect 30340 14776 31171 14804
rect 30340 14764 30346 14776
rect 31159 14773 31171 14776
rect 31205 14773 31217 14807
rect 32398 14804 32404 14816
rect 32359 14776 32404 14804
rect 31159 14767 31217 14773
rect 32398 14764 32404 14776
rect 32456 14764 32462 14816
rect 36814 14764 36820 14816
rect 36872 14804 36878 14816
rect 37734 14804 37740 14816
rect 36872 14776 37740 14804
rect 36872 14764 36878 14776
rect 37734 14764 37740 14776
rect 37792 14804 37798 14816
rect 37921 14807 37979 14813
rect 37921 14804 37933 14807
rect 37792 14776 37933 14804
rect 37792 14764 37798 14776
rect 37921 14773 37933 14776
rect 37967 14773 37979 14807
rect 39942 14804 39948 14816
rect 39855 14776 39948 14804
rect 37921 14767 37979 14773
rect 39942 14764 39948 14776
rect 40000 14804 40006 14816
rect 41800 14804 41828 14844
rect 42242 14832 42248 14844
rect 42300 14832 42306 14884
rect 43530 14832 43536 14884
rect 43588 14872 43594 14884
rect 43588 14844 43633 14872
rect 43588 14832 43594 14844
rect 46290 14832 46296 14884
rect 46348 14872 46354 14884
rect 46348 14844 46393 14872
rect 46348 14832 46354 14844
rect 40000 14776 41828 14804
rect 40000 14764 40006 14776
rect 41874 14764 41880 14816
rect 41932 14804 41938 14816
rect 45143 14807 45201 14813
rect 45143 14804 45155 14807
rect 41932 14776 45155 14804
rect 41932 14764 41938 14776
rect 45143 14773 45155 14776
rect 45189 14773 45201 14807
rect 45143 14767 45201 14773
rect 1104 14714 48852 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 48852 14714
rect 1104 14640 48852 14662
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21232 14572 21925 14600
rect 21232 14560 21238 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 21913 14563 21971 14569
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 25222 14600 25228 14612
rect 23624 14572 25228 14600
rect 23624 14560 23630 14572
rect 25222 14560 25228 14572
rect 25280 14560 25286 14612
rect 30558 14600 30564 14612
rect 30519 14572 30564 14600
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 33778 14600 33784 14612
rect 33739 14572 33784 14600
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 33962 14560 33968 14612
rect 34020 14600 34026 14612
rect 34057 14603 34115 14609
rect 34057 14600 34069 14603
rect 34020 14572 34069 14600
rect 34020 14560 34026 14572
rect 34057 14569 34069 14572
rect 34103 14569 34115 14603
rect 35526 14600 35532 14612
rect 35487 14572 35532 14600
rect 34057 14563 34115 14569
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 36446 14600 36452 14612
rect 36407 14572 36452 14600
rect 36446 14560 36452 14572
rect 36504 14560 36510 14612
rect 38749 14603 38807 14609
rect 38749 14569 38761 14603
rect 38795 14600 38807 14603
rect 40586 14600 40592 14612
rect 38795 14572 40080 14600
rect 40547 14572 40592 14600
rect 38795 14569 38807 14572
rect 38749 14563 38807 14569
rect 17420 14464 17448 14560
rect 18690 14492 18696 14544
rect 18748 14492 18754 14544
rect 19886 14492 19892 14544
rect 19944 14532 19950 14544
rect 20165 14535 20223 14541
rect 20165 14532 20177 14535
rect 19944 14504 20177 14532
rect 19944 14492 19950 14504
rect 20165 14501 20177 14504
rect 20211 14501 20223 14535
rect 20165 14495 20223 14501
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 21085 14535 21143 14541
rect 21085 14532 21097 14535
rect 20864 14504 21097 14532
rect 20864 14492 20870 14504
rect 21085 14501 21097 14504
rect 21131 14501 21143 14535
rect 21085 14495 21143 14501
rect 21637 14535 21695 14541
rect 21637 14501 21649 14535
rect 21683 14532 21695 14535
rect 21726 14532 21732 14544
rect 21683 14504 21732 14532
rect 21683 14501 21695 14504
rect 21637 14495 21695 14501
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 23290 14492 23296 14544
rect 23348 14532 23354 14544
rect 23385 14535 23443 14541
rect 23385 14532 23397 14535
rect 23348 14504 23397 14532
rect 23348 14492 23354 14504
rect 23385 14501 23397 14504
rect 23431 14501 23443 14535
rect 24946 14532 24952 14544
rect 24907 14504 24952 14532
rect 23385 14495 23443 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 25501 14535 25559 14541
rect 25501 14501 25513 14535
rect 25547 14532 25559 14535
rect 26694 14532 26700 14544
rect 25547 14504 26700 14532
rect 25547 14501 25559 14504
rect 25501 14495 25559 14501
rect 26694 14492 26700 14504
rect 26752 14492 26758 14544
rect 26786 14492 26792 14544
rect 26844 14532 26850 14544
rect 27065 14535 27123 14541
rect 27065 14532 27077 14535
rect 26844 14504 27077 14532
rect 26844 14492 26850 14504
rect 27065 14501 27077 14504
rect 27111 14501 27123 14535
rect 27065 14495 27123 14501
rect 29270 14492 29276 14544
rect 29328 14532 29334 14544
rect 29457 14535 29515 14541
rect 29457 14532 29469 14535
rect 29328 14504 29469 14532
rect 29328 14492 29334 14504
rect 29457 14501 29469 14504
rect 29503 14532 29515 14535
rect 29733 14535 29791 14541
rect 29733 14532 29745 14535
rect 29503 14504 29745 14532
rect 29503 14501 29515 14504
rect 29457 14495 29515 14501
rect 29733 14501 29745 14504
rect 29779 14501 29791 14535
rect 32858 14532 32864 14544
rect 32819 14504 32864 14532
rect 29733 14495 29791 14501
rect 32858 14492 32864 14504
rect 32916 14492 32922 14544
rect 33502 14532 33508 14544
rect 33060 14504 33508 14532
rect 17957 14467 18015 14473
rect 17957 14464 17969 14467
rect 17420 14436 17969 14464
rect 17957 14433 17969 14436
rect 18003 14433 18015 14467
rect 17957 14427 18015 14433
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 19300 14436 19441 14464
rect 19300 14424 19306 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 28718 14464 28724 14476
rect 28679 14436 28724 14464
rect 19429 14427 19487 14433
rect 28718 14424 28724 14436
rect 28776 14424 28782 14476
rect 29181 14467 29239 14473
rect 29181 14433 29193 14467
rect 29227 14464 29239 14467
rect 29362 14464 29368 14476
rect 29227 14436 29368 14464
rect 29227 14433 29239 14436
rect 29181 14427 29239 14433
rect 29362 14424 29368 14436
rect 29420 14424 29426 14476
rect 30561 14467 30619 14473
rect 30561 14433 30573 14467
rect 30607 14433 30619 14467
rect 30561 14427 30619 14433
rect 30837 14467 30895 14473
rect 30837 14433 30849 14467
rect 30883 14464 30895 14467
rect 31754 14464 31760 14476
rect 30883 14436 31760 14464
rect 30883 14433 30895 14436
rect 30837 14427 30895 14433
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 20990 14396 20996 14408
rect 20951 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 23290 14396 23296 14408
rect 23251 14368 23296 14396
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 23937 14399 23995 14405
rect 23937 14365 23949 14399
rect 23983 14396 23995 14399
rect 24394 14396 24400 14408
rect 23983 14368 24400 14396
rect 23983 14365 23995 14368
rect 23937 14359 23995 14365
rect 24394 14356 24400 14368
rect 24452 14396 24458 14408
rect 24854 14396 24860 14408
rect 24452 14368 24860 14396
rect 24452 14356 24458 14368
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 26418 14356 26424 14408
rect 26476 14396 26482 14408
rect 26697 14399 26755 14405
rect 26697 14396 26709 14399
rect 26476 14368 26709 14396
rect 26476 14356 26482 14368
rect 26697 14365 26709 14368
rect 26743 14365 26755 14399
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 26697 14359 26755 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27338 14396 27344 14408
rect 27299 14368 27344 14396
rect 27338 14356 27344 14368
rect 27396 14356 27402 14408
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 30576 14396 30604 14427
rect 31754 14424 31760 14436
rect 31812 14424 31818 14476
rect 33060 14473 33088 14504
rect 33502 14492 33508 14504
rect 33560 14492 33566 14544
rect 35161 14535 35219 14541
rect 35161 14501 35173 14535
rect 35207 14532 35219 14535
rect 35250 14532 35256 14544
rect 35207 14504 35256 14532
rect 35207 14501 35219 14504
rect 35161 14495 35219 14501
rect 35250 14492 35256 14504
rect 35308 14492 35314 14544
rect 38010 14492 38016 14544
rect 38068 14532 38074 14544
rect 38150 14535 38208 14541
rect 38150 14532 38162 14535
rect 38068 14504 38162 14532
rect 38068 14492 38074 14504
rect 38150 14501 38162 14504
rect 38196 14501 38208 14535
rect 38150 14495 38208 14501
rect 39761 14535 39819 14541
rect 39761 14501 39773 14535
rect 39807 14532 39819 14535
rect 39942 14532 39948 14544
rect 39807 14504 39948 14532
rect 39807 14501 39819 14504
rect 39761 14495 39819 14501
rect 39942 14492 39948 14504
rect 40000 14492 40006 14544
rect 40052 14532 40080 14572
rect 40586 14560 40592 14572
rect 40644 14560 40650 14612
rect 43165 14603 43223 14609
rect 43165 14600 43177 14603
rect 42766 14572 43177 14600
rect 41966 14532 41972 14544
rect 40052 14504 41972 14532
rect 41966 14492 41972 14504
rect 42024 14532 42030 14544
rect 42613 14535 42671 14541
rect 42613 14532 42625 14535
rect 42024 14504 42625 14532
rect 42024 14492 42030 14504
rect 42613 14501 42625 14504
rect 42659 14501 42671 14535
rect 42613 14495 42671 14501
rect 33045 14467 33103 14473
rect 33045 14433 33057 14467
rect 33091 14433 33103 14467
rect 33045 14427 33103 14433
rect 35069 14467 35127 14473
rect 35069 14433 35081 14467
rect 35115 14433 35127 14467
rect 35069 14427 35127 14433
rect 33134 14396 33140 14408
rect 30156 14368 33140 14396
rect 30156 14356 30162 14368
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 33410 14396 33416 14408
rect 33371 14368 33416 14396
rect 33410 14356 33416 14368
rect 33468 14356 33474 14408
rect 34606 14356 34612 14408
rect 34664 14396 34670 14408
rect 35084 14396 35112 14427
rect 35618 14424 35624 14476
rect 35676 14464 35682 14476
rect 35989 14467 36047 14473
rect 35989 14464 36001 14467
rect 35676 14436 36001 14464
rect 35676 14424 35682 14436
rect 35989 14433 36001 14436
rect 36035 14464 36047 14467
rect 36262 14464 36268 14476
rect 36035 14436 36268 14464
rect 36035 14433 36047 14436
rect 35989 14427 36047 14433
rect 36262 14424 36268 14436
rect 36320 14424 36326 14476
rect 40313 14467 40371 14473
rect 40313 14433 40325 14467
rect 40359 14464 40371 14467
rect 40770 14464 40776 14476
rect 40359 14436 40776 14464
rect 40359 14433 40371 14436
rect 40313 14427 40371 14433
rect 40770 14424 40776 14436
rect 40828 14424 40834 14476
rect 41208 14467 41266 14473
rect 41208 14433 41220 14467
rect 41254 14464 41266 14467
rect 41598 14464 41604 14476
rect 41254 14436 41604 14464
rect 41254 14433 41266 14436
rect 41208 14427 41266 14433
rect 41598 14424 41604 14436
rect 41656 14424 41662 14476
rect 42058 14424 42064 14476
rect 42116 14464 42122 14476
rect 42188 14467 42246 14473
rect 42188 14464 42200 14467
rect 42116 14436 42200 14464
rect 42116 14424 42122 14436
rect 42188 14433 42200 14436
rect 42234 14433 42246 14467
rect 42188 14427 42246 14433
rect 35158 14396 35164 14408
rect 34664 14368 35164 14396
rect 34664 14356 34670 14368
rect 35158 14356 35164 14368
rect 35216 14356 35222 14408
rect 37826 14396 37832 14408
rect 37787 14368 37832 14396
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 39666 14396 39672 14408
rect 39627 14368 39672 14396
rect 39666 14356 39672 14368
rect 39724 14356 39730 14408
rect 40788 14396 40816 14424
rect 42766 14396 42794 14572
rect 43165 14569 43177 14572
rect 43211 14600 43223 14603
rect 43438 14600 43444 14612
rect 43211 14572 43444 14600
rect 43211 14569 43223 14572
rect 43165 14563 43223 14569
rect 43438 14560 43444 14572
rect 43496 14560 43502 14612
rect 43530 14560 43536 14612
rect 43588 14600 43594 14612
rect 43717 14603 43775 14609
rect 43717 14600 43729 14603
rect 43588 14572 43729 14600
rect 43588 14560 43594 14572
rect 43717 14569 43729 14572
rect 43763 14569 43775 14603
rect 43717 14563 43775 14569
rect 46201 14603 46259 14609
rect 46201 14569 46213 14603
rect 46247 14600 46259 14603
rect 46290 14600 46296 14612
rect 46247 14572 46296 14600
rect 46247 14569 46259 14572
rect 46201 14563 46259 14569
rect 46290 14560 46296 14572
rect 46348 14560 46354 14612
rect 43990 14492 43996 14544
rect 44048 14532 44054 14544
rect 45186 14532 45192 14544
rect 44048 14504 45192 14532
rect 44048 14492 44054 14504
rect 45186 14492 45192 14504
rect 45244 14492 45250 14544
rect 45281 14535 45339 14541
rect 45281 14501 45293 14535
rect 45327 14532 45339 14535
rect 45554 14532 45560 14544
rect 45327 14504 45560 14532
rect 45327 14501 45339 14504
rect 45281 14495 45339 14501
rect 45554 14492 45560 14504
rect 45612 14492 45618 14544
rect 45830 14532 45836 14544
rect 45791 14504 45836 14532
rect 45830 14492 45836 14504
rect 45888 14532 45894 14544
rect 46477 14535 46535 14541
rect 46477 14532 46489 14535
rect 45888 14504 46489 14532
rect 45888 14492 45894 14504
rect 46477 14501 46489 14504
rect 46523 14501 46535 14535
rect 46477 14495 46535 14501
rect 43714 14464 43720 14476
rect 43675 14436 43720 14464
rect 43714 14424 43720 14436
rect 43772 14424 43778 14476
rect 46014 14424 46020 14476
rect 46072 14464 46078 14476
rect 46696 14467 46754 14473
rect 46696 14464 46708 14467
rect 46072 14436 46708 14464
rect 46072 14424 46078 14436
rect 46696 14433 46708 14436
rect 46742 14464 46754 14467
rect 46842 14464 46848 14476
rect 46742 14436 46848 14464
rect 46742 14433 46754 14436
rect 46696 14427 46754 14433
rect 46842 14424 46848 14436
rect 46900 14424 46906 14476
rect 40788 14368 42794 14396
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19889 14331 19947 14337
rect 19889 14328 19901 14331
rect 19484 14300 19901 14328
rect 19484 14288 19490 14300
rect 19889 14297 19901 14300
rect 19935 14297 19947 14331
rect 33152 14328 33180 14356
rect 34330 14328 34336 14340
rect 33152 14300 34336 14328
rect 19889 14291 19947 14297
rect 34330 14288 34336 14300
rect 34388 14288 34394 14340
rect 28258 14260 28264 14272
rect 28219 14232 28264 14260
rect 28258 14220 28264 14232
rect 28316 14220 28322 14272
rect 35802 14220 35808 14272
rect 35860 14260 35866 14272
rect 36173 14263 36231 14269
rect 36173 14260 36185 14263
rect 35860 14232 36185 14260
rect 35860 14220 35866 14232
rect 36173 14229 36185 14232
rect 36219 14229 36231 14263
rect 36173 14223 36231 14229
rect 36354 14220 36360 14272
rect 36412 14260 36418 14272
rect 36906 14260 36912 14272
rect 36412 14232 36912 14260
rect 36412 14220 36418 14232
rect 36906 14220 36912 14232
rect 36964 14220 36970 14272
rect 41279 14263 41337 14269
rect 41279 14229 41291 14263
rect 41325 14260 41337 14263
rect 41414 14260 41420 14272
rect 41325 14232 41420 14260
rect 41325 14229 41337 14232
rect 41279 14223 41337 14229
rect 41414 14220 41420 14232
rect 41472 14220 41478 14272
rect 41598 14260 41604 14272
rect 41559 14232 41604 14260
rect 41598 14220 41604 14232
rect 41656 14220 41662 14272
rect 42291 14263 42349 14269
rect 42291 14229 42303 14263
rect 42337 14260 42349 14263
rect 42426 14260 42432 14272
rect 42337 14232 42432 14260
rect 42337 14229 42349 14232
rect 42291 14223 42349 14229
rect 42426 14220 42432 14232
rect 42484 14220 42490 14272
rect 46799 14263 46857 14269
rect 46799 14229 46811 14263
rect 46845 14260 46857 14263
rect 46934 14260 46940 14272
rect 46845 14232 46940 14260
rect 46845 14229 46857 14232
rect 46799 14223 46857 14229
rect 46934 14220 46940 14232
rect 46992 14220 46998 14272
rect 1104 14170 48852 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 48852 14170
rect 1104 14096 48852 14118
rect 16485 14059 16543 14065
rect 16485 14025 16497 14059
rect 16531 14056 16543 14059
rect 17586 14056 17592 14068
rect 16531 14028 17592 14056
rect 16531 14025 16543 14028
rect 16485 14019 16543 14025
rect 17586 14016 17592 14028
rect 17644 14056 17650 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17644 14028 17693 14056
rect 17644 14016 17650 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 17696 13920 17724 14019
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20864 14028 20913 14056
rect 20864 14016 20870 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 23198 14056 23204 14068
rect 23159 14028 23204 14056
rect 20901 14019 20959 14025
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23348 14028 23857 14056
rect 23348 14016 23354 14028
rect 23845 14025 23857 14028
rect 23891 14025 23903 14059
rect 23845 14019 23903 14025
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25777 14059 25835 14065
rect 25777 14056 25789 14059
rect 24912 14028 25789 14056
rect 24912 14016 24918 14028
rect 25777 14025 25789 14028
rect 25823 14025 25835 14059
rect 25777 14019 25835 14025
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 26786 14056 26792 14068
rect 26375 14028 26792 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 26786 14016 26792 14028
rect 26844 14016 26850 14068
rect 29457 14059 29515 14065
rect 29457 14025 29469 14059
rect 29503 14025 29515 14059
rect 30098 14056 30104 14068
rect 30059 14028 30104 14056
rect 29457 14019 29515 14025
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 21637 13991 21695 13997
rect 21637 13988 21649 13991
rect 20680 13960 21649 13988
rect 20680 13948 20686 13960
rect 21637 13957 21649 13960
rect 21683 13988 21695 13991
rect 24302 13988 24308 14000
rect 21683 13960 22140 13988
rect 24215 13960 24308 13988
rect 21683 13957 21695 13960
rect 21637 13951 21695 13957
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 17696 13892 18061 13920
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13920 18475 13923
rect 19058 13920 19064 13932
rect 18463 13892 19064 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 21818 13920 21824 13932
rect 21407 13892 21824 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22112 13920 22140 13960
rect 24302 13948 24308 13960
rect 24360 13988 24366 14000
rect 24946 13988 24952 14000
rect 24360 13960 24952 13988
rect 24360 13948 24366 13960
rect 24946 13948 24952 13960
rect 25004 13988 25010 14000
rect 25317 13991 25375 13997
rect 25317 13988 25329 13991
rect 25004 13960 25329 13988
rect 25004 13948 25010 13960
rect 25317 13957 25329 13960
rect 25363 13957 25375 13991
rect 25317 13951 25375 13957
rect 29270 13948 29276 14000
rect 29328 13988 29334 14000
rect 29472 13988 29500 14019
rect 30098 14016 30104 14028
rect 30156 14016 30162 14068
rect 31478 14056 31484 14068
rect 31439 14028 31484 14056
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 31754 14056 31760 14068
rect 31715 14028 31760 14056
rect 31754 14016 31760 14028
rect 31812 14016 31818 14068
rect 32858 14016 32864 14068
rect 32916 14056 32922 14068
rect 33505 14059 33563 14065
rect 33505 14056 33517 14059
rect 32916 14028 33517 14056
rect 32916 14016 32922 14028
rect 33505 14025 33517 14028
rect 33551 14025 33563 14059
rect 33505 14019 33563 14025
rect 34333 14059 34391 14065
rect 34333 14025 34345 14059
rect 34379 14056 34391 14059
rect 34606 14056 34612 14068
rect 34379 14028 34612 14056
rect 34379 14025 34391 14028
rect 34333 14019 34391 14025
rect 34606 14016 34612 14028
rect 34664 14016 34670 14068
rect 34698 14016 34704 14068
rect 34756 14056 34762 14068
rect 35345 14059 35403 14065
rect 35345 14056 35357 14059
rect 34756 14028 35357 14056
rect 34756 14016 34762 14028
rect 35345 14025 35357 14028
rect 35391 14025 35403 14059
rect 36262 14056 36268 14068
rect 36223 14028 36268 14056
rect 35345 14019 35403 14025
rect 36262 14016 36268 14028
rect 36320 14016 36326 14068
rect 37826 14016 37832 14068
rect 37884 14056 37890 14068
rect 38565 14059 38623 14065
rect 38565 14056 38577 14059
rect 37884 14028 38577 14056
rect 37884 14016 37890 14028
rect 38565 14025 38577 14028
rect 38611 14025 38623 14059
rect 38565 14019 38623 14025
rect 39666 14016 39672 14068
rect 39724 14056 39730 14068
rect 39945 14059 40003 14065
rect 39945 14056 39957 14059
rect 39724 14028 39957 14056
rect 39724 14016 39730 14028
rect 39945 14025 39957 14028
rect 39991 14056 40003 14059
rect 40635 14059 40693 14065
rect 40635 14056 40647 14059
rect 39991 14028 40647 14056
rect 39991 14025 40003 14028
rect 39945 14019 40003 14025
rect 40635 14025 40647 14028
rect 40681 14025 40693 14059
rect 40635 14019 40693 14025
rect 43165 14059 43223 14065
rect 43165 14025 43177 14059
rect 43211 14056 43223 14059
rect 43714 14056 43720 14068
rect 43211 14028 43720 14056
rect 43211 14025 43223 14028
rect 43165 14019 43223 14025
rect 43714 14016 43720 14028
rect 43772 14016 43778 14068
rect 45186 14016 45192 14068
rect 45244 14056 45250 14068
rect 45465 14059 45523 14065
rect 45465 14056 45477 14059
rect 45244 14028 45477 14056
rect 45244 14016 45250 14028
rect 45465 14025 45477 14028
rect 45511 14025 45523 14059
rect 46842 14056 46848 14068
rect 46803 14028 46848 14056
rect 45465 14019 45523 14025
rect 46842 14016 46848 14028
rect 46900 14056 46906 14068
rect 47213 14059 47271 14065
rect 47213 14056 47225 14059
rect 46900 14028 47225 14056
rect 46900 14016 46906 14028
rect 47213 14025 47225 14028
rect 47259 14025 47271 14059
rect 47213 14019 47271 14025
rect 31772 13988 31800 14016
rect 29328 13960 31800 13988
rect 34624 13988 34652 14016
rect 35023 13991 35081 13997
rect 35023 13988 35035 13991
rect 34624 13960 35035 13988
rect 29328 13948 29334 13960
rect 35023 13957 35035 13960
rect 35069 13957 35081 13991
rect 35023 13951 35081 13957
rect 35161 13991 35219 13997
rect 35161 13957 35173 13991
rect 35207 13988 35219 13991
rect 35434 13988 35440 14000
rect 35207 13960 35440 13988
rect 35207 13957 35219 13960
rect 35161 13951 35219 13957
rect 35434 13948 35440 13960
rect 35492 13988 35498 14000
rect 35897 13991 35955 13997
rect 35897 13988 35909 13991
rect 35492 13960 35909 13988
rect 35492 13948 35498 13960
rect 35897 13957 35909 13960
rect 35943 13957 35955 13991
rect 35897 13951 35955 13957
rect 37921 13991 37979 13997
rect 37921 13957 37933 13991
rect 37967 13988 37979 13991
rect 37967 13960 40575 13988
rect 37967 13957 37979 13960
rect 37921 13951 37979 13957
rect 25133 13923 25191 13929
rect 22112 13892 22232 13920
rect 17862 13852 17868 13864
rect 17823 13824 17868 13852
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 19889 13855 19947 13861
rect 19889 13852 19901 13855
rect 19392 13824 19901 13852
rect 19392 13812 19398 13824
rect 19889 13821 19901 13824
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 22204 13796 22232 13892
rect 25133 13889 25145 13923
rect 25179 13920 25191 13923
rect 25774 13920 25780 13932
rect 25179 13892 25780 13920
rect 25179 13889 25191 13892
rect 25133 13883 25191 13889
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 27062 13920 27068 13932
rect 26620 13892 27068 13920
rect 26620 13861 26648 13892
rect 27062 13880 27068 13892
rect 27120 13880 27126 13932
rect 27338 13920 27344 13932
rect 27299 13892 27344 13920
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 30558 13920 30564 13932
rect 30519 13892 30564 13920
rect 30558 13880 30564 13892
rect 30616 13880 30622 13932
rect 32861 13923 32919 13929
rect 32861 13889 32873 13923
rect 32907 13920 32919 13923
rect 35250 13920 35256 13932
rect 32907 13892 35112 13920
rect 35211 13892 35256 13920
rect 32907 13889 32919 13892
rect 32861 13883 32919 13889
rect 25317 13855 25375 13861
rect 25317 13821 25329 13855
rect 25363 13852 25375 13855
rect 25409 13855 25467 13861
rect 25409 13852 25421 13855
rect 25363 13824 25421 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 25409 13821 25421 13824
rect 25455 13852 25467 13855
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 25455 13824 26617 13852
rect 25455 13821 25467 13824
rect 25409 13815 25467 13821
rect 26605 13821 26617 13824
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 28445 13855 28503 13861
rect 28445 13821 28457 13855
rect 28491 13852 28503 13855
rect 29273 13855 29331 13861
rect 29273 13852 29285 13855
rect 28491 13824 29285 13852
rect 28491 13821 28503 13824
rect 28445 13815 28503 13821
rect 29273 13821 29285 13824
rect 29319 13852 29331 13855
rect 29362 13852 29368 13864
rect 29319 13824 29368 13852
rect 29319 13821 29331 13824
rect 29273 13815 29331 13821
rect 29362 13812 29368 13824
rect 29420 13812 29426 13864
rect 29917 13855 29975 13861
rect 29917 13821 29929 13855
rect 29963 13852 29975 13855
rect 30469 13855 30527 13861
rect 30469 13852 30481 13855
rect 29963 13824 30481 13852
rect 29963 13821 29975 13824
rect 29917 13815 29975 13821
rect 30469 13821 30481 13824
rect 30515 13852 30527 13855
rect 30515 13824 30947 13852
rect 30515 13821 30527 13824
rect 30469 13815 30527 13821
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 17129 13787 17187 13793
rect 17129 13784 17141 13787
rect 16264 13756 17141 13784
rect 16264 13744 16270 13756
rect 17129 13753 17141 13756
rect 17175 13784 17187 13787
rect 17497 13787 17555 13793
rect 17497 13784 17509 13787
rect 17175 13756 17509 13784
rect 17175 13753 17187 13756
rect 17129 13747 17187 13753
rect 17497 13753 17509 13756
rect 17543 13784 17555 13787
rect 17954 13784 17960 13796
rect 17543 13756 17960 13784
rect 17543 13753 17555 13756
rect 17497 13747 17555 13753
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18782 13744 18788 13796
rect 18840 13744 18846 13796
rect 22186 13793 22192 13796
rect 22183 13747 22192 13793
rect 22244 13784 22250 13796
rect 24486 13784 24492 13796
rect 22244 13756 22337 13784
rect 24447 13756 24492 13784
rect 22186 13744 22192 13747
rect 22244 13744 22250 13756
rect 24486 13744 24492 13756
rect 24544 13744 24550 13796
rect 24581 13787 24639 13793
rect 24581 13753 24593 13787
rect 24627 13753 24639 13787
rect 24581 13747 24639 13753
rect 26881 13787 26939 13793
rect 26881 13753 26893 13787
rect 26927 13753 26939 13787
rect 26881 13747 26939 13753
rect 26973 13787 27031 13793
rect 26973 13753 26985 13787
rect 27019 13784 27031 13787
rect 27062 13784 27068 13796
rect 27019 13756 27068 13784
rect 27019 13753 27031 13756
rect 26973 13747 27031 13753
rect 16853 13719 16911 13725
rect 16853 13685 16865 13719
rect 16899 13716 16911 13719
rect 17034 13716 17040 13728
rect 16899 13688 17040 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 20349 13719 20407 13725
rect 20349 13685 20361 13719
rect 20395 13716 20407 13719
rect 20898 13716 20904 13728
rect 20395 13688 20904 13716
rect 20395 13685 20407 13688
rect 20349 13679 20407 13685
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 22738 13716 22744 13728
rect 22699 13688 22744 13716
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 24302 13676 24308 13728
rect 24360 13716 24366 13728
rect 24596 13716 24624 13747
rect 24360 13688 24624 13716
rect 26896 13716 26924 13747
rect 27062 13744 27068 13756
rect 27120 13744 27126 13796
rect 28718 13784 28724 13796
rect 28679 13756 28724 13784
rect 28718 13744 28724 13756
rect 28776 13784 28782 13796
rect 30919 13793 30947 13824
rect 31938 13812 31944 13864
rect 31996 13852 32002 13864
rect 32217 13855 32275 13861
rect 32217 13852 32229 13855
rect 31996 13824 32229 13852
rect 31996 13812 32002 13824
rect 32217 13821 32229 13824
rect 32263 13852 32275 13855
rect 32309 13855 32367 13861
rect 32309 13852 32321 13855
rect 32263 13824 32321 13852
rect 32263 13821 32275 13824
rect 32217 13815 32275 13821
rect 32309 13821 32321 13824
rect 32355 13821 32367 13855
rect 32309 13815 32367 13821
rect 32398 13812 32404 13864
rect 32456 13852 32462 13864
rect 32493 13855 32551 13861
rect 32493 13852 32505 13855
rect 32456 13824 32505 13852
rect 32456 13812 32462 13824
rect 32493 13821 32505 13824
rect 32539 13852 32551 13855
rect 32766 13852 32772 13864
rect 32539 13824 32772 13852
rect 32539 13821 32551 13824
rect 32493 13815 32551 13821
rect 32766 13812 32772 13824
rect 32824 13852 32830 13864
rect 33137 13855 33195 13861
rect 33137 13852 33149 13855
rect 32824 13824 33149 13852
rect 32824 13812 32830 13824
rect 33137 13821 33149 13824
rect 33183 13821 33195 13855
rect 33137 13815 33195 13821
rect 33410 13812 33416 13864
rect 33468 13852 33474 13864
rect 33689 13855 33747 13861
rect 33689 13852 33701 13855
rect 33468 13824 33701 13852
rect 33468 13812 33474 13824
rect 33689 13821 33701 13824
rect 33735 13821 33747 13855
rect 33689 13815 33747 13821
rect 30902 13787 30960 13793
rect 28776 13756 30788 13784
rect 28776 13744 28782 13756
rect 27798 13716 27804 13728
rect 26896 13688 27804 13716
rect 24360 13676 24366 13688
rect 27798 13676 27804 13688
rect 27856 13676 27862 13728
rect 28534 13676 28540 13728
rect 28592 13716 28598 13728
rect 29454 13716 29460 13728
rect 28592 13688 29460 13716
rect 28592 13676 28598 13688
rect 29454 13676 29460 13688
rect 29512 13716 29518 13728
rect 29917 13719 29975 13725
rect 29917 13716 29929 13719
rect 29512 13688 29929 13716
rect 29512 13676 29518 13688
rect 29917 13685 29929 13688
rect 29963 13685 29975 13719
rect 30760 13716 30788 13756
rect 30902 13753 30914 13787
rect 30948 13753 30960 13787
rect 30902 13747 30960 13753
rect 34514 13744 34520 13796
rect 34572 13784 34578 13796
rect 34885 13787 34943 13793
rect 34885 13784 34897 13787
rect 34572 13756 34897 13784
rect 34572 13744 34578 13756
rect 34885 13753 34897 13756
rect 34931 13753 34943 13787
rect 35084 13784 35112 13892
rect 35250 13880 35256 13892
rect 35308 13880 35314 13932
rect 36909 13923 36967 13929
rect 36909 13889 36921 13923
rect 36955 13920 36967 13923
rect 37182 13920 37188 13932
rect 36955 13892 37188 13920
rect 36955 13889 36967 13892
rect 36909 13883 36967 13889
rect 37182 13880 37188 13892
rect 37240 13920 37246 13932
rect 38010 13920 38016 13932
rect 37240 13892 38016 13920
rect 37240 13880 37246 13892
rect 38010 13880 38016 13892
rect 38068 13920 38074 13932
rect 38197 13923 38255 13929
rect 38197 13920 38209 13923
rect 38068 13892 38209 13920
rect 38068 13880 38074 13892
rect 38197 13889 38209 13892
rect 38243 13889 38255 13923
rect 38197 13883 38255 13889
rect 39669 13923 39727 13929
rect 39669 13889 39681 13923
rect 39715 13920 39727 13923
rect 39942 13920 39948 13932
rect 39715 13892 39948 13920
rect 39715 13889 39727 13892
rect 39669 13883 39727 13889
rect 39942 13880 39948 13892
rect 40000 13880 40006 13932
rect 36998 13852 37004 13864
rect 36959 13824 37004 13852
rect 36998 13812 37004 13824
rect 37056 13812 37062 13864
rect 40547 13861 40575 13960
rect 42886 13948 42892 14000
rect 42944 13988 42950 14000
rect 43441 13991 43499 13997
rect 43441 13988 43453 13991
rect 42944 13960 43453 13988
rect 42944 13948 42950 13960
rect 43441 13957 43453 13960
rect 43487 13988 43499 13991
rect 43806 13988 43812 14000
rect 43487 13960 43812 13988
rect 43487 13957 43499 13960
rect 43441 13951 43499 13957
rect 43806 13948 43812 13960
rect 43864 13948 43870 14000
rect 41414 13880 41420 13932
rect 41472 13920 41478 13932
rect 41693 13923 41751 13929
rect 41693 13920 41705 13923
rect 41472 13892 41705 13920
rect 41472 13880 41478 13892
rect 41693 13889 41705 13892
rect 41739 13889 41751 13923
rect 41693 13883 41751 13889
rect 38749 13855 38807 13861
rect 38749 13852 38761 13855
rect 37108 13824 38761 13852
rect 37108 13784 37136 13824
rect 38749 13821 38761 13824
rect 38795 13852 38807 13855
rect 39209 13855 39267 13861
rect 39209 13852 39221 13855
rect 38795 13824 39221 13852
rect 38795 13821 38807 13824
rect 38749 13815 38807 13821
rect 39209 13821 39221 13824
rect 39255 13821 39267 13855
rect 39209 13815 39267 13821
rect 40532 13855 40590 13861
rect 40532 13821 40544 13855
rect 40578 13852 40590 13855
rect 40957 13855 41015 13861
rect 40957 13852 40969 13855
rect 40578 13824 40969 13852
rect 40578 13821 40590 13824
rect 40532 13815 40590 13821
rect 40957 13821 40969 13824
rect 41003 13821 41015 13855
rect 40957 13815 41015 13821
rect 46385 13855 46443 13861
rect 46385 13821 46397 13855
rect 46431 13852 46443 13855
rect 46842 13852 46848 13864
rect 46431 13824 46848 13852
rect 46431 13821 46443 13824
rect 46385 13815 46443 13821
rect 46842 13812 46848 13824
rect 46900 13812 46906 13864
rect 35084 13756 37136 13784
rect 41785 13787 41843 13793
rect 34885 13747 34943 13753
rect 41785 13753 41797 13787
rect 41831 13753 41843 13787
rect 42334 13784 42340 13796
rect 42295 13756 42340 13784
rect 41785 13747 41843 13753
rect 32398 13716 32404 13728
rect 30760 13688 32404 13716
rect 29917 13679 29975 13685
rect 32398 13676 32404 13688
rect 32456 13676 32462 13728
rect 33870 13716 33876 13728
rect 33831 13688 33876 13716
rect 33870 13676 33876 13688
rect 33928 13676 33934 13728
rect 37182 13676 37188 13728
rect 37240 13716 37246 13728
rect 37363 13719 37421 13725
rect 37363 13716 37375 13719
rect 37240 13688 37375 13716
rect 37240 13676 37246 13688
rect 37363 13685 37375 13688
rect 37409 13685 37421 13719
rect 38930 13716 38936 13728
rect 38891 13688 38936 13716
rect 37363 13679 37421 13685
rect 38930 13676 38936 13688
rect 38988 13676 38994 13728
rect 41509 13719 41567 13725
rect 41509 13685 41521 13719
rect 41555 13716 41567 13719
rect 41690 13716 41696 13728
rect 41555 13688 41696 13716
rect 41555 13685 41567 13688
rect 41509 13679 41567 13685
rect 41690 13676 41696 13688
rect 41748 13716 41754 13728
rect 41800 13716 41828 13747
rect 42334 13744 42340 13756
rect 42392 13784 42398 13796
rect 43717 13787 43775 13793
rect 43717 13784 43729 13787
rect 42392 13756 43729 13784
rect 42392 13744 42398 13756
rect 43717 13753 43729 13756
rect 43763 13753 43775 13787
rect 43717 13747 43775 13753
rect 41966 13716 41972 13728
rect 41748 13688 41972 13716
rect 41748 13676 41754 13688
rect 41966 13676 41972 13688
rect 42024 13676 42030 13728
rect 42058 13676 42064 13728
rect 42116 13716 42122 13728
rect 42613 13719 42671 13725
rect 42613 13716 42625 13719
rect 42116 13688 42625 13716
rect 42116 13676 42122 13688
rect 42613 13685 42625 13688
rect 42659 13685 42671 13719
rect 43732 13716 43760 13747
rect 43806 13744 43812 13796
rect 43864 13784 43870 13796
rect 44358 13784 44364 13796
rect 43864 13756 43909 13784
rect 44319 13756 44364 13784
rect 43864 13744 43870 13756
rect 44358 13744 44364 13756
rect 44416 13744 44422 13796
rect 44637 13719 44695 13725
rect 44637 13716 44649 13719
rect 43732 13688 44649 13716
rect 42613 13679 42671 13685
rect 44637 13685 44649 13688
rect 44683 13685 44695 13719
rect 44637 13679 44695 13685
rect 45189 13719 45247 13725
rect 45189 13685 45201 13719
rect 45235 13716 45247 13719
rect 45462 13716 45468 13728
rect 45235 13688 45468 13716
rect 45235 13685 45247 13688
rect 45189 13679 45247 13685
rect 45462 13676 45468 13688
rect 45520 13676 45526 13728
rect 46566 13716 46572 13728
rect 46527 13688 46572 13716
rect 46566 13676 46572 13688
rect 46624 13676 46630 13728
rect 1104 13626 48852 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 48852 13626
rect 1104 13552 48852 13574
rect 18414 13512 18420 13524
rect 18375 13484 18420 13512
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 19058 13512 19064 13524
rect 19019 13484 19064 13512
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 20990 13512 20996 13524
rect 20949 13484 20996 13512
rect 20990 13472 20996 13484
rect 21048 13521 21054 13524
rect 21048 13515 21097 13521
rect 21048 13481 21051 13515
rect 21085 13512 21097 13515
rect 21361 13515 21419 13521
rect 21361 13512 21373 13515
rect 21085 13484 21373 13512
rect 21085 13481 21097 13484
rect 21048 13475 21097 13481
rect 21361 13481 21373 13484
rect 21407 13481 21419 13515
rect 24486 13512 24492 13524
rect 24447 13484 24492 13512
rect 21361 13475 21419 13481
rect 21048 13472 21054 13475
rect 24486 13472 24492 13484
rect 24544 13472 24550 13524
rect 25130 13512 25136 13524
rect 25043 13484 25136 13512
rect 17126 13404 17132 13456
rect 17184 13404 17190 13456
rect 22186 13404 22192 13456
rect 22244 13444 22250 13456
rect 22510 13447 22568 13453
rect 22510 13444 22522 13447
rect 22244 13416 22522 13444
rect 22244 13404 22250 13416
rect 22510 13413 22522 13416
rect 22556 13444 22568 13447
rect 22830 13444 22836 13456
rect 22556 13416 22836 13444
rect 22556 13413 22568 13416
rect 22510 13407 22568 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 25056 13453 25084 13484
rect 25130 13472 25136 13484
rect 25188 13512 25194 13524
rect 25188 13484 26740 13512
rect 25188 13472 25194 13484
rect 25041 13447 25099 13453
rect 25041 13413 25053 13447
rect 25087 13413 25099 13447
rect 25041 13407 25099 13413
rect 25593 13447 25651 13453
rect 25593 13413 25605 13447
rect 25639 13444 25651 13447
rect 25774 13444 25780 13456
rect 25639 13416 25780 13444
rect 25639 13413 25651 13416
rect 25593 13407 25651 13413
rect 25774 13404 25780 13416
rect 25832 13404 25838 13456
rect 26712 13453 26740 13484
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 29549 13515 29607 13521
rect 29549 13512 29561 13515
rect 29420 13484 29561 13512
rect 29420 13472 29426 13484
rect 29549 13481 29561 13484
rect 29595 13481 29607 13515
rect 29549 13475 29607 13481
rect 30558 13472 30564 13524
rect 30616 13512 30622 13524
rect 31205 13515 31263 13521
rect 31205 13512 31217 13515
rect 30616 13484 31217 13512
rect 30616 13472 30622 13484
rect 31205 13481 31217 13484
rect 31251 13481 31263 13515
rect 31205 13475 31263 13481
rect 33410 13472 33416 13524
rect 33468 13512 33474 13524
rect 33781 13515 33839 13521
rect 33781 13512 33793 13515
rect 33468 13484 33793 13512
rect 33468 13472 33474 13484
rect 33781 13481 33793 13484
rect 33827 13481 33839 13515
rect 34514 13512 34520 13524
rect 34475 13484 34520 13512
rect 33781 13475 33839 13481
rect 34514 13472 34520 13484
rect 34572 13472 34578 13524
rect 35250 13472 35256 13524
rect 35308 13512 35314 13524
rect 35437 13515 35495 13521
rect 35437 13512 35449 13515
rect 35308 13484 35449 13512
rect 35308 13472 35314 13484
rect 35437 13481 35449 13484
rect 35483 13481 35495 13515
rect 35437 13475 35495 13481
rect 41506 13472 41512 13524
rect 41564 13512 41570 13524
rect 41693 13515 41751 13521
rect 41693 13512 41705 13515
rect 41564 13484 41705 13512
rect 41564 13472 41570 13484
rect 41693 13481 41705 13484
rect 41739 13481 41751 13515
rect 41693 13475 41751 13481
rect 26697 13447 26755 13453
rect 26697 13413 26709 13447
rect 26743 13444 26755 13447
rect 26786 13444 26792 13456
rect 26743 13416 26792 13444
rect 26743 13413 26755 13416
rect 26697 13407 26755 13413
rect 26786 13404 26792 13416
rect 26844 13404 26850 13456
rect 28534 13404 28540 13456
rect 28592 13444 28598 13456
rect 28674 13447 28732 13453
rect 28674 13444 28686 13447
rect 28592 13416 28686 13444
rect 28592 13404 28598 13416
rect 28674 13413 28686 13416
rect 28720 13413 28732 13447
rect 28674 13407 28732 13413
rect 30098 13404 30104 13456
rect 30156 13444 30162 13456
rect 30374 13444 30380 13456
rect 30156 13416 30380 13444
rect 30156 13404 30162 13416
rect 30374 13404 30380 13416
rect 30432 13404 30438 13456
rect 32585 13447 32643 13453
rect 32585 13413 32597 13447
rect 32631 13444 32643 13447
rect 32858 13444 32864 13456
rect 32631 13416 32864 13444
rect 32631 13413 32643 13416
rect 32585 13407 32643 13413
rect 32858 13404 32864 13416
rect 32916 13404 32922 13456
rect 33137 13447 33195 13453
rect 33137 13413 33149 13447
rect 33183 13444 33195 13447
rect 36725 13447 36783 13453
rect 33183 13416 36445 13444
rect 33183 13413 33195 13416
rect 33137 13407 33195 13413
rect 17954 13376 17960 13388
rect 17915 13348 17960 13376
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13376 20867 13379
rect 20898 13376 20904 13388
rect 20855 13348 20904 13376
rect 20855 13345 20867 13348
rect 20809 13339 20867 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 23109 13379 23167 13385
rect 23109 13345 23121 13379
rect 23155 13376 23167 13379
rect 24762 13376 24768 13388
rect 23155 13348 24768 13376
rect 23155 13345 23167 13348
rect 23109 13339 23167 13345
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 28258 13336 28264 13388
rect 28316 13376 28322 13388
rect 29273 13379 29331 13385
rect 29273 13376 29285 13379
rect 28316 13348 29285 13376
rect 28316 13336 28322 13348
rect 29273 13345 29285 13348
rect 29319 13345 29331 13379
rect 32766 13376 32772 13388
rect 32679 13348 32772 13376
rect 29273 13339 29331 13345
rect 32766 13336 32772 13348
rect 32824 13336 32830 13388
rect 34609 13379 34667 13385
rect 34609 13345 34621 13379
rect 34655 13376 34667 13379
rect 34698 13376 34704 13388
rect 34655 13348 34704 13376
rect 34655 13345 34667 13348
rect 34609 13339 34667 13345
rect 34698 13336 34704 13348
rect 34756 13336 34762 13388
rect 34790 13336 34796 13388
rect 34848 13376 34854 13388
rect 35986 13376 35992 13388
rect 34848 13348 34893 13376
rect 35947 13348 35992 13376
rect 34848 13336 34854 13348
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 16942 13308 16948 13320
rect 16531 13280 16948 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13308 19395 13311
rect 20990 13308 20996 13320
rect 19383 13280 20996 13308
rect 19383 13277 19395 13280
rect 19337 13271 19395 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 24946 13308 24952 13320
rect 24907 13280 24952 13308
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 26602 13308 26608 13320
rect 26563 13280 26608 13308
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 26881 13311 26939 13317
rect 26881 13308 26893 13311
rect 26752 13280 26893 13308
rect 26752 13268 26758 13280
rect 26881 13277 26893 13280
rect 26927 13277 26939 13311
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 26881 13271 26939 13277
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 30282 13308 30288 13320
rect 30195 13280 30288 13308
rect 30282 13268 30288 13280
rect 30340 13308 30346 13320
rect 30650 13308 30656 13320
rect 30340 13280 30656 13308
rect 30340 13268 30346 13280
rect 30650 13268 30656 13280
rect 30708 13268 30714 13320
rect 32582 13268 32588 13320
rect 32640 13308 32646 13320
rect 32784 13308 32812 13336
rect 32640 13280 32812 13308
rect 35161 13311 35219 13317
rect 32640 13268 32646 13280
rect 35161 13277 35173 13311
rect 35207 13308 35219 13311
rect 36170 13308 36176 13320
rect 35207 13280 36176 13308
rect 35207 13277 35219 13280
rect 35161 13271 35219 13277
rect 36170 13268 36176 13280
rect 36228 13268 36234 13320
rect 36417 13308 36445 13416
rect 36725 13413 36737 13447
rect 36771 13444 36783 13447
rect 36998 13444 37004 13456
rect 36771 13416 37004 13444
rect 36771 13413 36783 13416
rect 36725 13407 36783 13413
rect 36998 13404 37004 13416
rect 37056 13404 37062 13456
rect 39114 13444 39120 13456
rect 38396 13416 39120 13444
rect 36541 13379 36599 13385
rect 36541 13345 36553 13379
rect 36587 13376 36599 13379
rect 37274 13376 37280 13388
rect 36587 13348 37280 13376
rect 36587 13345 36599 13348
rect 36541 13339 36599 13345
rect 37274 13336 37280 13348
rect 37332 13336 37338 13388
rect 37918 13376 37924 13388
rect 37879 13348 37924 13376
rect 37918 13336 37924 13348
rect 37976 13336 37982 13388
rect 38396 13385 38424 13416
rect 39114 13404 39120 13416
rect 39172 13404 39178 13456
rect 40859 13447 40917 13453
rect 40859 13413 40871 13447
rect 40905 13444 40917 13447
rect 40954 13444 40960 13456
rect 40905 13416 40960 13444
rect 40905 13413 40917 13416
rect 40859 13407 40917 13413
rect 40954 13404 40960 13416
rect 41012 13404 41018 13456
rect 43438 13404 43444 13456
rect 43496 13444 43502 13456
rect 43809 13447 43867 13453
rect 43809 13444 43821 13447
rect 43496 13416 43821 13444
rect 43496 13404 43502 13416
rect 43809 13413 43821 13416
rect 43855 13413 43867 13447
rect 45370 13444 45376 13456
rect 45331 13416 45376 13444
rect 43809 13407 43867 13413
rect 45370 13404 45376 13416
rect 45428 13404 45434 13456
rect 45462 13404 45468 13456
rect 45520 13444 45526 13456
rect 46753 13447 46811 13453
rect 46753 13444 46765 13447
rect 45520 13416 46765 13444
rect 45520 13404 45526 13416
rect 46753 13413 46765 13416
rect 46799 13413 46811 13447
rect 46753 13407 46811 13413
rect 38381 13379 38439 13385
rect 38381 13345 38393 13379
rect 38427 13345 38439 13379
rect 39485 13379 39543 13385
rect 39485 13376 39497 13379
rect 38381 13339 38439 13345
rect 38488 13348 39497 13376
rect 38488 13308 38516 13348
rect 39485 13345 39497 13348
rect 39531 13376 39543 13379
rect 39850 13376 39856 13388
rect 39531 13348 39856 13376
rect 39531 13345 39543 13348
rect 39485 13339 39543 13345
rect 39850 13336 39856 13348
rect 39908 13336 39914 13388
rect 41417 13379 41475 13385
rect 41417 13345 41429 13379
rect 41463 13376 41475 13379
rect 42312 13379 42370 13385
rect 42312 13376 42324 13379
rect 41463 13348 42324 13376
rect 41463 13345 41475 13348
rect 41417 13339 41475 13345
rect 42312 13345 42324 13348
rect 42358 13376 42370 13379
rect 42610 13376 42616 13388
rect 42358 13348 42616 13376
rect 42358 13345 42370 13348
rect 42312 13339 42370 13345
rect 42610 13336 42616 13348
rect 42668 13336 42674 13388
rect 46934 13336 46940 13388
rect 46992 13376 46998 13388
rect 47118 13376 47124 13388
rect 46992 13348 47124 13376
rect 46992 13336 46998 13348
rect 47118 13336 47124 13348
rect 47176 13336 47182 13388
rect 38654 13308 38660 13320
rect 36417 13280 38516 13308
rect 38567 13280 38660 13308
rect 38654 13268 38660 13280
rect 38712 13308 38718 13320
rect 38933 13311 38991 13317
rect 38933 13308 38945 13311
rect 38712 13280 38945 13308
rect 38712 13268 38718 13280
rect 38933 13277 38945 13280
rect 38979 13277 38991 13311
rect 38933 13271 38991 13277
rect 40310 13268 40316 13320
rect 40368 13308 40374 13320
rect 40497 13311 40555 13317
rect 40497 13308 40509 13311
rect 40368 13280 40509 13308
rect 40368 13268 40374 13280
rect 40497 13277 40509 13280
rect 40543 13277 40555 13311
rect 43714 13308 43720 13320
rect 43675 13280 43720 13308
rect 40497 13271 40555 13277
rect 43714 13268 43720 13280
rect 43772 13268 43778 13320
rect 44358 13308 44364 13320
rect 44271 13280 44364 13308
rect 44358 13268 44364 13280
rect 44416 13308 44422 13320
rect 45278 13308 45284 13320
rect 44416 13280 45284 13308
rect 44416 13268 44422 13280
rect 45278 13268 45284 13280
rect 45336 13268 45342 13320
rect 27798 13200 27804 13252
rect 27856 13240 27862 13252
rect 30742 13240 30748 13252
rect 27856 13212 30748 13240
rect 27856 13200 27862 13212
rect 30742 13200 30748 13212
rect 30800 13240 30806 13252
rect 30837 13243 30895 13249
rect 30837 13240 30849 13243
rect 30800 13212 30849 13240
rect 30800 13200 30806 13212
rect 30837 13209 30849 13212
rect 30883 13209 30895 13243
rect 45830 13240 45836 13252
rect 45791 13212 45836 13240
rect 30837 13203 30895 13209
rect 45830 13200 45836 13212
rect 45888 13200 45894 13252
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 17184 13144 18705 13172
rect 17184 13132 17190 13144
rect 18693 13141 18705 13144
rect 18739 13172 18751 13175
rect 18782 13172 18788 13184
rect 18739 13144 18788 13172
rect 18739 13141 18751 13144
rect 18693 13135 18751 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 21913 13175 21971 13181
rect 21913 13141 21925 13175
rect 21959 13172 21971 13175
rect 22002 13172 22008 13184
rect 21959 13144 22008 13172
rect 21959 13141 21971 13144
rect 21913 13135 21971 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 26329 13175 26387 13181
rect 26329 13141 26341 13175
rect 26375 13172 26387 13175
rect 27062 13172 27068 13184
rect 26375 13144 27068 13172
rect 26375 13141 26387 13144
rect 26329 13135 26387 13141
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 27709 13175 27767 13181
rect 27709 13141 27721 13175
rect 27755 13172 27767 13175
rect 28074 13172 28080 13184
rect 27755 13144 28080 13172
rect 27755 13141 27767 13144
rect 27709 13135 27767 13141
rect 28074 13132 28080 13144
rect 28132 13172 28138 13184
rect 29270 13172 29276 13184
rect 28132 13144 29276 13172
rect 28132 13132 28138 13144
rect 29270 13132 29276 13144
rect 29328 13132 29334 13184
rect 33502 13172 33508 13184
rect 33463 13144 33508 13172
rect 33502 13132 33508 13144
rect 33560 13132 33566 13184
rect 39666 13172 39672 13184
rect 39627 13144 39672 13172
rect 39666 13132 39672 13144
rect 39724 13132 39730 13184
rect 40405 13175 40463 13181
rect 40405 13141 40417 13175
rect 40451 13172 40463 13175
rect 40954 13172 40960 13184
rect 40451 13144 40960 13172
rect 40451 13141 40463 13144
rect 40405 13135 40463 13141
rect 40954 13132 40960 13144
rect 41012 13132 41018 13184
rect 42150 13172 42156 13184
rect 42111 13144 42156 13172
rect 42150 13132 42156 13144
rect 42208 13132 42214 13184
rect 42383 13175 42441 13181
rect 42383 13141 42395 13175
rect 42429 13172 42441 13175
rect 43530 13172 43536 13184
rect 42429 13144 43536 13172
rect 42429 13141 42441 13144
rect 42383 13135 42441 13141
rect 43530 13132 43536 13144
rect 43588 13132 43594 13184
rect 46290 13172 46296 13184
rect 46251 13144 46296 13172
rect 46290 13132 46296 13144
rect 46348 13132 46354 13184
rect 1104 13082 48852 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 48852 13082
rect 1104 13008 48852 13030
rect 15841 12971 15899 12977
rect 15841 12937 15853 12971
rect 15887 12968 15899 12971
rect 16114 12968 16120 12980
rect 15887 12940 16120 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 17773 12971 17831 12977
rect 17773 12937 17785 12971
rect 17819 12968 17831 12971
rect 17862 12968 17868 12980
rect 17819 12940 17868 12968
rect 17819 12937 17831 12940
rect 17773 12931 17831 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 22830 12968 22836 12980
rect 22791 12940 22836 12968
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 24578 12968 24584 12980
rect 24539 12940 24584 12968
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 25130 12968 25136 12980
rect 25091 12940 25136 12968
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 26786 12928 26792 12980
rect 26844 12968 26850 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 26844 12940 26985 12968
rect 26844 12928 26850 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 30650 12968 30656 12980
rect 30611 12940 30656 12968
rect 26973 12931 27031 12937
rect 30650 12928 30656 12940
rect 30708 12928 30714 12980
rect 32217 12971 32275 12977
rect 32217 12937 32229 12971
rect 32263 12968 32275 12971
rect 33597 12971 33655 12977
rect 33597 12968 33609 12971
rect 32263 12940 33609 12968
rect 32263 12937 32275 12940
rect 32217 12931 32275 12937
rect 18248 12832 18276 12928
rect 27062 12860 27068 12912
rect 27120 12900 27126 12912
rect 30006 12900 30012 12912
rect 27120 12872 30012 12900
rect 27120 12860 27126 12872
rect 30006 12860 30012 12872
rect 30064 12860 30070 12912
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18248 12804 18797 12832
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22244 12804 22385 12832
rect 22244 12792 22250 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23799 12835 23857 12841
rect 23799 12832 23811 12835
rect 23348 12804 23811 12832
rect 23348 12792 23354 12804
rect 23799 12801 23811 12804
rect 23845 12801 23857 12835
rect 26326 12832 26332 12844
rect 23799 12795 23857 12801
rect 26252 12804 26332 12832
rect 21729 12767 21787 12773
rect 21729 12733 21741 12767
rect 21775 12764 21787 12767
rect 22094 12764 22100 12776
rect 21775 12736 22100 12764
rect 21775 12733 21787 12736
rect 21729 12727 21787 12733
rect 22094 12724 22100 12736
rect 22152 12724 22158 12776
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 16577 12699 16635 12705
rect 16577 12665 16589 12699
rect 16623 12696 16635 12699
rect 17126 12696 17132 12708
rect 16623 12668 17132 12696
rect 16623 12665 16635 12668
rect 16577 12659 16635 12665
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 19242 12656 19248 12708
rect 19300 12696 19306 12708
rect 19334 12696 19340 12708
rect 19300 12668 19340 12696
rect 19300 12656 19306 12668
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 22002 12656 22008 12708
rect 22060 12696 22066 12708
rect 22296 12696 22324 12727
rect 22738 12724 22744 12776
rect 22796 12764 22802 12776
rect 23712 12767 23770 12773
rect 23712 12764 23724 12767
rect 22796 12736 23724 12764
rect 22796 12724 22802 12736
rect 23712 12733 23724 12736
rect 23758 12764 23770 12767
rect 24121 12767 24179 12773
rect 24121 12764 24133 12767
rect 23758 12736 24133 12764
rect 23758 12733 23770 12736
rect 23712 12727 23770 12733
rect 24121 12733 24133 12736
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 24578 12724 24584 12776
rect 24636 12764 24642 12776
rect 24673 12767 24731 12773
rect 24673 12764 24685 12767
rect 24636 12736 24685 12764
rect 24636 12724 24642 12736
rect 24673 12733 24685 12736
rect 24719 12764 24731 12767
rect 24719 12736 25636 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 25608 12696 25636 12736
rect 25682 12724 25688 12776
rect 25740 12764 25746 12776
rect 26252 12773 26280 12804
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 26510 12832 26516 12844
rect 26471 12804 26516 12832
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 28350 12832 28356 12844
rect 28311 12804 28356 12832
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 28626 12792 28632 12844
rect 28684 12832 28690 12844
rect 29362 12832 29368 12844
rect 28684 12804 29368 12832
rect 28684 12792 28690 12804
rect 29362 12792 29368 12804
rect 29420 12792 29426 12844
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 25740 12736 25881 12764
rect 25740 12724 25746 12736
rect 25869 12733 25881 12736
rect 25915 12764 25927 12767
rect 26237 12767 26295 12773
rect 26237 12764 26249 12767
rect 25915 12736 26249 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 26237 12733 26249 12736
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 26421 12767 26479 12773
rect 26421 12733 26433 12767
rect 26467 12733 26479 12767
rect 26421 12727 26479 12733
rect 27525 12767 27583 12773
rect 27525 12733 27537 12767
rect 27571 12764 27583 12767
rect 27890 12764 27896 12776
rect 27571 12736 27896 12764
rect 27571 12733 27583 12736
rect 27525 12727 27583 12733
rect 26050 12696 26056 12708
rect 22060 12668 24900 12696
rect 25608 12668 26056 12696
rect 22060 12656 22066 12668
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16942 12628 16948 12640
rect 16855 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12628 17006 12640
rect 17954 12628 17960 12640
rect 17000 12600 17960 12628
rect 17000 12588 17006 12600
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 18564 12600 18705 12628
rect 18564 12588 18570 12600
rect 18693 12597 18705 12600
rect 18739 12628 18751 12631
rect 19153 12631 19211 12637
rect 19153 12628 19165 12631
rect 18739 12600 19165 12628
rect 18739 12597 18751 12600
rect 18693 12591 18751 12597
rect 19153 12597 19165 12600
rect 19199 12628 19211 12631
rect 19260 12628 19288 12656
rect 24872 12640 24900 12668
rect 26050 12656 26056 12668
rect 26108 12696 26114 12708
rect 26436 12696 26464 12727
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 28074 12764 28080 12776
rect 28035 12736 28080 12764
rect 28074 12724 28080 12736
rect 28132 12724 28138 12776
rect 32324 12773 32352 12940
rect 33597 12937 33609 12940
rect 33643 12937 33655 12971
rect 37274 12968 37280 12980
rect 37235 12940 37280 12968
rect 33597 12931 33655 12937
rect 37274 12928 37280 12940
rect 37332 12928 37338 12980
rect 39577 12971 39635 12977
rect 39577 12937 39589 12971
rect 39623 12968 39635 12971
rect 41598 12968 41604 12980
rect 39623 12940 41604 12968
rect 39623 12937 39635 12940
rect 39577 12931 39635 12937
rect 41598 12928 41604 12940
rect 41656 12928 41662 12980
rect 43165 12971 43223 12977
rect 43165 12937 43177 12971
rect 43211 12968 43223 12971
rect 43438 12968 43444 12980
rect 43211 12940 43444 12968
rect 43211 12937 43223 12940
rect 43165 12931 43223 12937
rect 43438 12928 43444 12940
rect 43496 12928 43502 12980
rect 47118 12968 47124 12980
rect 47079 12940 47124 12968
rect 47118 12928 47124 12940
rect 47176 12928 47182 12980
rect 32398 12860 32404 12912
rect 32456 12900 32462 12912
rect 32493 12903 32551 12909
rect 32493 12900 32505 12903
rect 32456 12872 32505 12900
rect 32456 12860 32462 12872
rect 32493 12869 32505 12872
rect 32539 12869 32551 12903
rect 32493 12863 32551 12869
rect 30904 12767 30962 12773
rect 30904 12733 30916 12767
rect 30950 12764 30962 12767
rect 32309 12767 32367 12773
rect 30950 12736 31340 12764
rect 30950 12733 30962 12736
rect 30904 12727 30962 12733
rect 29086 12696 29092 12708
rect 26108 12668 26464 12696
rect 28999 12668 29092 12696
rect 26108 12656 26114 12668
rect 19199 12600 19288 12628
rect 19705 12631 19763 12637
rect 19199 12597 19211 12600
rect 19153 12591 19211 12597
rect 19705 12597 19717 12631
rect 19751 12628 19763 12631
rect 21082 12628 21088 12640
rect 19751 12600 21088 12628
rect 19751 12597 19763 12600
rect 19705 12591 19763 12597
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 24854 12628 24860 12640
rect 24815 12600 24860 12628
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 28534 12588 28540 12640
rect 28592 12628 28598 12640
rect 28629 12631 28687 12637
rect 28629 12628 28641 12631
rect 28592 12600 28641 12628
rect 28592 12588 28598 12600
rect 28629 12597 28641 12600
rect 28675 12597 28687 12631
rect 28629 12591 28687 12597
rect 28902 12588 28908 12640
rect 28960 12628 28966 12640
rect 29012 12637 29040 12668
rect 29086 12656 29092 12668
rect 29144 12696 29150 12708
rect 29457 12699 29515 12705
rect 29457 12696 29469 12699
rect 29144 12668 29469 12696
rect 29144 12656 29150 12668
rect 29457 12665 29469 12668
rect 29503 12665 29515 12699
rect 30006 12696 30012 12708
rect 29967 12668 30012 12696
rect 29457 12659 29515 12665
rect 30006 12656 30012 12668
rect 30064 12656 30070 12708
rect 31312 12640 31340 12736
rect 32309 12733 32321 12767
rect 32355 12733 32367 12767
rect 32309 12727 32367 12733
rect 32508 12696 32536 12863
rect 32858 12860 32864 12912
rect 32916 12900 32922 12912
rect 33137 12903 33195 12909
rect 33137 12900 33149 12903
rect 32916 12872 33149 12900
rect 32916 12860 32922 12872
rect 33137 12869 33149 12872
rect 33183 12869 33195 12903
rect 35986 12900 35992 12912
rect 33137 12863 33195 12869
rect 34992 12872 35992 12900
rect 34992 12832 35020 12872
rect 35986 12860 35992 12872
rect 36044 12900 36050 12912
rect 36265 12903 36323 12909
rect 36265 12900 36277 12903
rect 36044 12872 36277 12900
rect 36044 12860 36050 12872
rect 36265 12869 36277 12872
rect 36311 12869 36323 12903
rect 39850 12900 39856 12912
rect 39811 12872 39856 12900
rect 36265 12863 36323 12869
rect 39850 12860 39856 12872
rect 39908 12860 39914 12912
rect 40313 12903 40371 12909
rect 40313 12869 40325 12903
rect 40359 12900 40371 12903
rect 40862 12900 40868 12912
rect 40359 12872 40868 12900
rect 40359 12869 40371 12872
rect 40313 12863 40371 12869
rect 40862 12860 40868 12872
rect 40920 12860 40926 12912
rect 35342 12832 35348 12844
rect 33106 12804 35020 12832
rect 35084 12804 35348 12832
rect 32950 12696 32956 12708
rect 32508 12668 32956 12696
rect 32950 12656 32956 12668
rect 33008 12696 33014 12708
rect 33106 12696 33134 12804
rect 33318 12764 33324 12776
rect 33279 12736 33324 12764
rect 33318 12724 33324 12736
rect 33376 12724 33382 12776
rect 33502 12764 33508 12776
rect 33415 12736 33508 12764
rect 33502 12724 33508 12736
rect 33560 12764 33566 12776
rect 35084 12773 35112 12804
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 35897 12835 35955 12841
rect 35897 12801 35909 12835
rect 35943 12832 35955 12835
rect 38102 12832 38108 12844
rect 35943 12804 38108 12832
rect 35943 12801 35955 12804
rect 35897 12795 35955 12801
rect 35069 12767 35127 12773
rect 33560 12736 34744 12764
rect 33560 12724 33566 12736
rect 33008 12668 33134 12696
rect 33336 12696 33364 12724
rect 34716 12705 34744 12736
rect 35069 12733 35081 12767
rect 35115 12733 35127 12767
rect 35069 12727 35127 12733
rect 35253 12767 35311 12773
rect 35253 12733 35265 12767
rect 35299 12764 35311 12767
rect 35912 12764 35940 12795
rect 38102 12792 38108 12804
rect 38160 12792 38166 12844
rect 38654 12832 38660 12844
rect 38615 12804 38660 12832
rect 38654 12792 38660 12804
rect 38712 12792 38718 12844
rect 41509 12835 41567 12841
rect 41509 12832 41521 12835
rect 40512 12804 41521 12832
rect 35299 12736 35940 12764
rect 35299 12733 35311 12736
rect 35253 12727 35311 12733
rect 34149 12699 34207 12705
rect 34149 12696 34161 12699
rect 33336 12668 34161 12696
rect 33008 12656 33014 12668
rect 34149 12665 34161 12668
rect 34195 12665 34207 12699
rect 34149 12659 34207 12665
rect 34701 12699 34759 12705
rect 34701 12665 34713 12699
rect 34747 12696 34759 12699
rect 34790 12696 34796 12708
rect 34747 12668 34796 12696
rect 34747 12665 34759 12668
rect 34701 12659 34759 12665
rect 34790 12656 34796 12668
rect 34848 12696 34854 12708
rect 35268 12696 35296 12727
rect 36170 12724 36176 12776
rect 36228 12764 36234 12776
rect 36449 12767 36507 12773
rect 36449 12764 36461 12767
rect 36228 12736 36461 12764
rect 36228 12724 36234 12736
rect 36449 12733 36461 12736
rect 36495 12764 36507 12767
rect 36909 12767 36967 12773
rect 36909 12764 36921 12767
rect 36495 12736 36921 12764
rect 36495 12733 36507 12736
rect 36449 12727 36507 12733
rect 36909 12733 36921 12736
rect 36955 12733 36967 12767
rect 36909 12727 36967 12733
rect 37274 12724 37280 12776
rect 37332 12764 37338 12776
rect 37461 12767 37519 12773
rect 37461 12764 37473 12767
rect 37332 12736 37473 12764
rect 37332 12724 37338 12736
rect 37461 12733 37473 12736
rect 37507 12733 37519 12767
rect 37461 12727 37519 12733
rect 38838 12724 38844 12776
rect 38896 12764 38902 12776
rect 40512 12773 40540 12804
rect 41509 12801 41521 12804
rect 41555 12801 41567 12835
rect 42150 12832 42156 12844
rect 42111 12804 42156 12832
rect 41509 12795 41567 12801
rect 42150 12792 42156 12804
rect 42208 12792 42214 12844
rect 42242 12792 42248 12844
rect 42300 12832 42306 12844
rect 42518 12832 42524 12844
rect 42300 12804 42524 12832
rect 42300 12792 42306 12804
rect 42518 12792 42524 12804
rect 42576 12792 42582 12844
rect 42797 12835 42855 12841
rect 42797 12801 42809 12835
rect 42843 12832 42855 12835
rect 43714 12832 43720 12844
rect 42843 12804 43720 12832
rect 42843 12801 42855 12804
rect 42797 12795 42855 12801
rect 43714 12792 43720 12804
rect 43772 12832 43778 12844
rect 43993 12835 44051 12841
rect 43993 12832 44005 12835
rect 43772 12804 44005 12832
rect 43772 12792 43778 12804
rect 43993 12801 44005 12804
rect 44039 12832 44051 12835
rect 44637 12835 44695 12841
rect 44637 12832 44649 12835
rect 44039 12804 44649 12832
rect 44039 12801 44051 12804
rect 43993 12795 44051 12801
rect 44637 12801 44649 12804
rect 44683 12801 44695 12835
rect 44637 12795 44695 12801
rect 46014 12792 46020 12844
rect 46072 12832 46078 12844
rect 46198 12832 46204 12844
rect 46072 12804 46204 12832
rect 46072 12792 46078 12804
rect 46198 12792 46204 12804
rect 46256 12832 46262 12844
rect 46477 12835 46535 12841
rect 46477 12832 46489 12835
rect 46256 12804 46489 12832
rect 46256 12792 46262 12804
rect 46477 12801 46489 12804
rect 46523 12801 46535 12835
rect 46477 12795 46535 12801
rect 40497 12767 40555 12773
rect 40497 12764 40509 12767
rect 38896 12736 40509 12764
rect 38896 12724 38902 12736
rect 40497 12733 40509 12736
rect 40543 12733 40555 12767
rect 40954 12764 40960 12776
rect 40915 12736 40960 12764
rect 40497 12727 40555 12733
rect 40954 12724 40960 12736
rect 41012 12724 41018 12776
rect 34848 12668 35296 12696
rect 35621 12699 35679 12705
rect 34848 12656 34854 12668
rect 35621 12665 35633 12699
rect 35667 12696 35679 12699
rect 36538 12696 36544 12708
rect 35667 12668 36544 12696
rect 35667 12665 35679 12668
rect 35621 12659 35679 12665
rect 36538 12656 36544 12668
rect 36596 12656 36602 12708
rect 37550 12696 37556 12708
rect 36648 12668 37556 12696
rect 28997 12631 29055 12637
rect 28997 12628 29009 12631
rect 28960 12600 29009 12628
rect 28960 12588 28966 12600
rect 28997 12597 29009 12600
rect 29043 12597 29055 12631
rect 28997 12591 29055 12597
rect 30098 12588 30104 12640
rect 30156 12628 30162 12640
rect 30285 12631 30343 12637
rect 30285 12628 30297 12631
rect 30156 12600 30297 12628
rect 30156 12588 30162 12600
rect 30285 12597 30297 12600
rect 30331 12597 30343 12631
rect 30285 12591 30343 12597
rect 30374 12588 30380 12640
rect 30432 12628 30438 12640
rect 30975 12631 31033 12637
rect 30975 12628 30987 12631
rect 30432 12600 30987 12628
rect 30432 12588 30438 12600
rect 30975 12597 30987 12600
rect 31021 12597 31033 12631
rect 31294 12628 31300 12640
rect 31255 12600 31300 12628
rect 30975 12591 31033 12597
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 32582 12588 32588 12640
rect 32640 12628 32646 12640
rect 36648 12637 36676 12668
rect 37550 12656 37556 12668
rect 37608 12696 37614 12708
rect 37918 12696 37924 12708
rect 37608 12668 37924 12696
rect 37608 12656 37614 12668
rect 37918 12656 37924 12668
rect 37976 12656 37982 12708
rect 38978 12699 39036 12705
rect 38978 12665 38990 12699
rect 39024 12665 39036 12699
rect 42245 12699 42303 12705
rect 42245 12696 42257 12699
rect 38978 12659 39036 12665
rect 41984 12668 42257 12696
rect 32769 12631 32827 12637
rect 32769 12628 32781 12631
rect 32640 12600 32781 12628
rect 32640 12588 32646 12600
rect 32769 12597 32781 12600
rect 32815 12597 32827 12631
rect 32769 12591 32827 12597
rect 36633 12631 36691 12637
rect 36633 12597 36645 12631
rect 36679 12597 36691 12631
rect 37642 12628 37648 12640
rect 37603 12600 37648 12628
rect 36633 12591 36691 12597
rect 37642 12588 37648 12600
rect 37700 12588 37706 12640
rect 38010 12588 38016 12640
rect 38068 12628 38074 12640
rect 38473 12631 38531 12637
rect 38473 12628 38485 12631
rect 38068 12600 38485 12628
rect 38068 12588 38074 12600
rect 38473 12597 38485 12600
rect 38519 12628 38531 12631
rect 38993 12628 39021 12659
rect 41984 12640 42012 12668
rect 42245 12665 42257 12668
rect 42291 12665 42303 12699
rect 43441 12699 43499 12705
rect 43441 12696 43453 12699
rect 42245 12659 42303 12665
rect 42996 12668 43453 12696
rect 38519 12600 39021 12628
rect 38519 12597 38531 12600
rect 38473 12591 38531 12597
rect 40310 12588 40316 12640
rect 40368 12628 40374 12640
rect 40589 12631 40647 12637
rect 40589 12628 40601 12631
rect 40368 12600 40601 12628
rect 40368 12588 40374 12600
rect 40589 12597 40601 12600
rect 40635 12597 40647 12631
rect 41966 12628 41972 12640
rect 41927 12600 41972 12628
rect 40589 12591 40647 12597
rect 41966 12588 41972 12600
rect 42024 12588 42030 12640
rect 42518 12588 42524 12640
rect 42576 12628 42582 12640
rect 42996 12628 43024 12668
rect 43441 12665 43453 12668
rect 43487 12665 43499 12699
rect 43441 12659 43499 12665
rect 42576 12600 43024 12628
rect 43456 12628 43484 12659
rect 43530 12656 43536 12708
rect 43588 12696 43594 12708
rect 43717 12699 43775 12705
rect 43717 12696 43729 12699
rect 43588 12668 43729 12696
rect 43588 12656 43594 12668
rect 43717 12665 43729 12668
rect 43763 12665 43775 12699
rect 43717 12659 43775 12665
rect 43809 12699 43867 12705
rect 43809 12665 43821 12699
rect 43855 12665 43867 12699
rect 43809 12659 43867 12665
rect 43824 12628 43852 12659
rect 44450 12656 44456 12708
rect 44508 12696 44514 12708
rect 46198 12696 46204 12708
rect 44508 12668 46204 12696
rect 44508 12656 44514 12668
rect 46198 12656 46204 12668
rect 46256 12656 46262 12708
rect 46293 12699 46351 12705
rect 46293 12665 46305 12699
rect 46339 12696 46351 12699
rect 46842 12696 46848 12708
rect 46339 12668 46848 12696
rect 46339 12665 46351 12668
rect 46293 12659 46351 12665
rect 43456 12600 43852 12628
rect 45281 12631 45339 12637
rect 42576 12588 42582 12600
rect 45281 12597 45293 12631
rect 45327 12628 45339 12631
rect 45370 12628 45376 12640
rect 45327 12600 45376 12628
rect 45327 12597 45339 12600
rect 45281 12591 45339 12597
rect 45370 12588 45376 12600
rect 45428 12628 45434 12640
rect 45925 12631 45983 12637
rect 45925 12628 45937 12631
rect 45428 12600 45937 12628
rect 45428 12588 45434 12600
rect 45925 12597 45937 12600
rect 45971 12628 45983 12631
rect 46308 12628 46336 12659
rect 46842 12656 46848 12668
rect 46900 12656 46906 12708
rect 45971 12600 46336 12628
rect 45971 12597 45983 12600
rect 45925 12591 45983 12597
rect 1104 12538 48852 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 48852 12538
rect 1104 12464 48852 12486
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 18417 12427 18475 12433
rect 18417 12424 18429 12427
rect 17920 12396 18429 12424
rect 17920 12384 17926 12396
rect 18417 12393 18429 12396
rect 18463 12393 18475 12427
rect 19334 12424 19340 12436
rect 19295 12396 19340 12424
rect 18417 12387 18475 12393
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 22186 12424 22192 12436
rect 22147 12396 22192 12424
rect 22186 12384 22192 12396
rect 22244 12384 22250 12436
rect 24762 12424 24768 12436
rect 24723 12396 24768 12424
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 26050 12424 26056 12436
rect 26011 12396 26056 12424
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 26697 12427 26755 12433
rect 26697 12424 26709 12427
rect 26660 12396 26709 12424
rect 26660 12384 26666 12396
rect 26697 12393 26709 12396
rect 26743 12424 26755 12427
rect 28350 12424 28356 12436
rect 26743 12396 27844 12424
rect 28311 12396 28356 12424
rect 26743 12393 26755 12396
rect 26697 12387 26755 12393
rect 27816 12368 27844 12396
rect 28350 12384 28356 12396
rect 28408 12384 28414 12436
rect 29362 12424 29368 12436
rect 29323 12396 29368 12424
rect 29362 12384 29368 12396
rect 29420 12384 29426 12436
rect 33318 12424 33324 12436
rect 33279 12396 33324 12424
rect 33318 12384 33324 12396
rect 33376 12384 33382 12436
rect 34698 12424 34704 12436
rect 34659 12396 34704 12424
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 35161 12427 35219 12433
rect 35161 12393 35173 12427
rect 35207 12424 35219 12427
rect 35342 12424 35348 12436
rect 35207 12396 35348 12424
rect 35207 12393 35219 12396
rect 35161 12387 35219 12393
rect 35342 12384 35348 12396
rect 35400 12384 35406 12436
rect 36078 12384 36084 12436
rect 36136 12424 36142 12436
rect 36173 12427 36231 12433
rect 36173 12424 36185 12427
rect 36136 12396 36185 12424
rect 36136 12384 36142 12396
rect 36173 12393 36185 12396
rect 36219 12424 36231 12427
rect 37274 12424 37280 12436
rect 36219 12396 37280 12424
rect 36219 12393 36231 12396
rect 36173 12387 36231 12393
rect 37274 12384 37280 12396
rect 37332 12384 37338 12436
rect 40310 12424 40316 12436
rect 40271 12396 40316 12424
rect 40310 12384 40316 12396
rect 40368 12384 40374 12436
rect 41325 12427 41383 12433
rect 41325 12393 41337 12427
rect 41371 12424 41383 12427
rect 42058 12424 42064 12436
rect 41371 12396 42064 12424
rect 41371 12393 41383 12396
rect 41325 12387 41383 12393
rect 42058 12384 42064 12396
rect 42116 12384 42122 12436
rect 42150 12384 42156 12436
rect 42208 12424 42214 12436
rect 42291 12427 42349 12433
rect 42291 12424 42303 12427
rect 42208 12396 42303 12424
rect 42208 12384 42214 12396
rect 42291 12393 42303 12396
rect 42337 12393 42349 12427
rect 42610 12424 42616 12436
rect 42571 12396 42616 12424
rect 42291 12387 42349 12393
rect 42610 12384 42616 12396
rect 42668 12384 42674 12436
rect 43530 12384 43536 12436
rect 43588 12424 43594 12436
rect 43809 12427 43867 12433
rect 43809 12424 43821 12427
rect 43588 12396 43821 12424
rect 43588 12384 43594 12396
rect 43809 12393 43821 12396
rect 43855 12393 43867 12427
rect 43809 12387 43867 12393
rect 45189 12427 45247 12433
rect 45189 12393 45201 12427
rect 45235 12424 45247 12427
rect 45278 12424 45284 12436
rect 45235 12396 45284 12424
rect 45235 12393 45247 12396
rect 45189 12387 45247 12393
rect 45278 12384 45284 12396
rect 45336 12384 45342 12436
rect 21082 12356 21088 12368
rect 21043 12328 21088 12356
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 23109 12359 23167 12365
rect 23109 12325 23121 12359
rect 23155 12356 23167 12359
rect 23198 12356 23204 12368
rect 23155 12328 23204 12356
rect 23155 12325 23167 12328
rect 23109 12319 23167 12325
rect 23198 12316 23204 12328
rect 23256 12316 23262 12368
rect 26786 12316 26792 12368
rect 26844 12356 26850 12368
rect 27249 12359 27307 12365
rect 27249 12356 27261 12359
rect 26844 12328 27261 12356
rect 26844 12316 26850 12328
rect 27249 12325 27261 12328
rect 27295 12325 27307 12359
rect 27798 12356 27804 12368
rect 27711 12328 27804 12356
rect 27249 12319 27307 12325
rect 27798 12316 27804 12328
rect 27856 12316 27862 12368
rect 28902 12316 28908 12368
rect 28960 12356 28966 12368
rect 30101 12359 30159 12365
rect 30101 12356 30113 12359
rect 28960 12328 30113 12356
rect 28960 12316 28966 12328
rect 30101 12325 30113 12328
rect 30147 12325 30159 12359
rect 30101 12319 30159 12325
rect 30653 12359 30711 12365
rect 30653 12325 30665 12359
rect 30699 12356 30711 12359
rect 30742 12356 30748 12368
rect 30699 12328 30748 12356
rect 30699 12325 30711 12328
rect 30653 12319 30711 12325
rect 30742 12316 30748 12328
rect 30800 12316 30806 12368
rect 32490 12356 32496 12368
rect 32451 12328 32496 12356
rect 32490 12316 32496 12328
rect 32548 12316 32554 12368
rect 33686 12316 33692 12368
rect 33744 12356 33750 12368
rect 33873 12359 33931 12365
rect 33873 12356 33885 12359
rect 33744 12328 33885 12356
rect 33744 12316 33750 12328
rect 33873 12325 33885 12328
rect 33919 12325 33931 12359
rect 33873 12319 33931 12325
rect 38010 12316 38016 12368
rect 38068 12356 38074 12368
rect 38150 12359 38208 12365
rect 38150 12356 38162 12359
rect 38068 12328 38162 12356
rect 38068 12316 38074 12328
rect 38150 12325 38162 12328
rect 38196 12325 38208 12359
rect 38150 12319 38208 12325
rect 40767 12359 40825 12365
rect 40767 12325 40779 12359
rect 40813 12356 40825 12359
rect 40862 12356 40868 12368
rect 40813 12328 40868 12356
rect 40813 12325 40825 12328
rect 40767 12319 40825 12325
rect 40862 12316 40868 12328
rect 40920 12316 40926 12368
rect 45462 12356 45468 12368
rect 45423 12328 45468 12356
rect 45462 12316 45468 12328
rect 45520 12316 45526 12368
rect 46014 12356 46020 12368
rect 45975 12328 46020 12356
rect 46014 12316 46020 12328
rect 46072 12316 46078 12368
rect 46842 12356 46848 12368
rect 46803 12328 46848 12356
rect 46842 12316 46848 12328
rect 46900 12316 46906 12368
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17402 12288 17408 12300
rect 17175 12260 17408 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 18966 12288 18972 12300
rect 18927 12260 18972 12288
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 24578 12288 24584 12300
rect 24539 12260 24584 12288
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24912 12260 25053 12288
rect 24912 12248 24918 12260
rect 25041 12257 25053 12260
rect 25087 12288 25099 12291
rect 26234 12288 26240 12300
rect 25087 12260 26240 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 26234 12248 26240 12260
rect 26292 12248 26298 12300
rect 28442 12248 28448 12300
rect 28500 12288 28506 12300
rect 28664 12291 28722 12297
rect 28664 12288 28676 12291
rect 28500 12260 28676 12288
rect 28500 12248 28506 12260
rect 28664 12257 28676 12260
rect 28710 12257 28722 12291
rect 28664 12251 28722 12257
rect 32582 12248 32588 12300
rect 32640 12288 32646 12300
rect 32677 12291 32735 12297
rect 32677 12288 32689 12291
rect 32640 12260 32689 12288
rect 32640 12248 32646 12260
rect 32677 12257 32689 12260
rect 32723 12257 32735 12291
rect 32677 12251 32735 12257
rect 34057 12291 34115 12297
rect 34057 12257 34069 12291
rect 34103 12288 34115 12291
rect 34790 12288 34796 12300
rect 34103 12260 34796 12288
rect 34103 12257 34115 12260
rect 34057 12251 34115 12257
rect 20990 12220 20996 12232
rect 20951 12192 20996 12220
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21266 12220 21272 12232
rect 21227 12192 21272 12220
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 28166 12220 28172 12232
rect 27203 12192 28172 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 28166 12180 28172 12192
rect 28224 12220 28230 12232
rect 28767 12223 28825 12229
rect 28767 12220 28779 12223
rect 28224 12192 28779 12220
rect 28224 12180 28230 12192
rect 28767 12189 28779 12192
rect 28813 12189 28825 12223
rect 28767 12183 28825 12189
rect 29086 12180 29092 12232
rect 29144 12220 29150 12232
rect 30009 12223 30067 12229
rect 30009 12220 30021 12223
rect 29144 12192 30021 12220
rect 29144 12180 29150 12192
rect 30009 12189 30021 12192
rect 30055 12220 30067 12223
rect 30374 12220 30380 12232
rect 30055 12192 30380 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 30374 12180 30380 12192
rect 30432 12180 30438 12232
rect 33045 12223 33103 12229
rect 33045 12189 33057 12223
rect 33091 12189 33103 12223
rect 33045 12183 33103 12189
rect 33781 12223 33839 12229
rect 33781 12189 33793 12223
rect 33827 12220 33839 12223
rect 33870 12220 33876 12232
rect 33827 12192 33876 12220
rect 33827 12189 33839 12192
rect 33781 12183 33839 12189
rect 23569 12155 23627 12161
rect 23569 12121 23581 12155
rect 23615 12152 23627 12155
rect 24486 12152 24492 12164
rect 23615 12124 24492 12152
rect 23615 12121 23627 12124
rect 23569 12115 23627 12121
rect 24486 12112 24492 12124
rect 24544 12112 24550 12164
rect 33060 12152 33088 12183
rect 33870 12180 33876 12192
rect 33928 12220 33934 12232
rect 34072 12220 34100 12251
rect 34790 12248 34796 12260
rect 34848 12248 34854 12300
rect 35621 12291 35679 12297
rect 35621 12257 35633 12291
rect 35667 12288 35679 12291
rect 36078 12288 36084 12300
rect 35667 12260 36084 12288
rect 35667 12257 35679 12260
rect 35621 12251 35679 12257
rect 36078 12248 36084 12260
rect 36136 12248 36142 12300
rect 36538 12248 36544 12300
rect 36596 12288 36602 12300
rect 36633 12291 36691 12297
rect 36633 12288 36645 12291
rect 36596 12260 36645 12288
rect 36596 12248 36602 12260
rect 36633 12257 36645 12260
rect 36679 12257 36691 12291
rect 36633 12251 36691 12257
rect 38749 12291 38807 12297
rect 38749 12257 38761 12291
rect 38795 12288 38807 12291
rect 42150 12288 42156 12300
rect 42208 12297 42214 12300
rect 42208 12291 42246 12297
rect 38795 12260 42156 12288
rect 38795 12257 38807 12260
rect 38749 12251 38807 12257
rect 42150 12248 42156 12260
rect 42234 12257 42246 12291
rect 42208 12251 42246 12257
rect 42208 12248 42214 12251
rect 43254 12248 43260 12300
rect 43312 12288 43318 12300
rect 43384 12291 43442 12297
rect 43384 12288 43396 12291
rect 43312 12260 43396 12288
rect 43312 12248 43318 12260
rect 43384 12257 43396 12260
rect 43430 12257 43442 12291
rect 43384 12251 43442 12257
rect 46566 12248 46572 12300
rect 46624 12288 46630 12300
rect 46937 12291 46995 12297
rect 46937 12288 46949 12291
rect 46624 12260 46949 12288
rect 46624 12248 46630 12260
rect 46937 12257 46949 12260
rect 46983 12257 46995 12291
rect 46937 12251 46995 12257
rect 34422 12220 34428 12232
rect 33928 12192 34100 12220
rect 34383 12192 34428 12220
rect 33928 12180 33934 12192
rect 34422 12180 34428 12192
rect 34480 12180 34486 12232
rect 37829 12223 37887 12229
rect 37829 12189 37841 12223
rect 37875 12220 37887 12223
rect 37918 12220 37924 12232
rect 37875 12192 37924 12220
rect 37875 12189 37887 12192
rect 37829 12183 37887 12189
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 40405 12223 40463 12229
rect 40405 12189 40417 12223
rect 40451 12220 40463 12223
rect 40586 12220 40592 12232
rect 40451 12192 40592 12220
rect 40451 12189 40463 12192
rect 40405 12183 40463 12189
rect 40586 12180 40592 12192
rect 40644 12180 40650 12232
rect 43622 12180 43628 12232
rect 43680 12220 43686 12232
rect 44726 12220 44732 12232
rect 43680 12192 44732 12220
rect 43680 12180 43686 12192
rect 44726 12180 44732 12192
rect 44784 12180 44790 12232
rect 45370 12220 45376 12232
rect 45331 12192 45376 12220
rect 45370 12180 45376 12192
rect 45428 12180 45434 12232
rect 36446 12152 36452 12164
rect 33060 12124 36452 12152
rect 36446 12112 36452 12124
rect 36504 12112 36510 12164
rect 36630 12112 36636 12164
rect 36688 12152 36694 12164
rect 36817 12155 36875 12161
rect 36817 12152 36829 12155
rect 36688 12124 36829 12152
rect 36688 12112 36694 12124
rect 36817 12121 36829 12124
rect 36863 12152 36875 12155
rect 38838 12152 38844 12164
rect 36863 12124 38844 12152
rect 36863 12121 36875 12124
rect 36817 12115 36875 12121
rect 38838 12112 38844 12124
rect 38896 12112 38902 12164
rect 19886 12084 19892 12096
rect 19847 12056 19892 12084
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 24397 12087 24455 12093
rect 24397 12053 24409 12087
rect 24443 12084 24455 12087
rect 24670 12084 24676 12096
rect 24443 12056 24676 12084
rect 24443 12053 24455 12056
rect 24397 12047 24455 12053
rect 24670 12044 24676 12056
rect 24728 12084 24734 12096
rect 24946 12084 24952 12096
rect 24728 12056 24952 12084
rect 24728 12044 24734 12056
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 25314 12044 25320 12096
rect 25372 12084 25378 12096
rect 25501 12087 25559 12093
rect 25501 12084 25513 12087
rect 25372 12056 25513 12084
rect 25372 12044 25378 12056
rect 25501 12053 25513 12056
rect 25547 12053 25559 12087
rect 35526 12084 35532 12096
rect 35439 12056 35532 12084
rect 25501 12047 25559 12053
rect 35526 12044 35532 12056
rect 35584 12084 35590 12096
rect 35805 12087 35863 12093
rect 35805 12084 35817 12087
rect 35584 12056 35817 12084
rect 35584 12044 35590 12056
rect 35805 12053 35817 12056
rect 35851 12053 35863 12087
rect 35805 12047 35863 12053
rect 37553 12087 37611 12093
rect 37553 12053 37565 12087
rect 37599 12084 37611 12087
rect 37642 12084 37648 12096
rect 37599 12056 37648 12084
rect 37599 12053 37611 12056
rect 37553 12047 37611 12053
rect 37642 12044 37648 12056
rect 37700 12044 37706 12096
rect 39114 12084 39120 12096
rect 39075 12056 39120 12084
rect 39114 12044 39120 12056
rect 39172 12044 39178 12096
rect 41782 12044 41788 12096
rect 41840 12084 41846 12096
rect 43487 12087 43545 12093
rect 43487 12084 43499 12087
rect 41840 12056 43499 12084
rect 41840 12044 41846 12056
rect 43487 12053 43499 12056
rect 43533 12053 43545 12087
rect 43487 12047 43545 12053
rect 43622 12044 43628 12096
rect 43680 12084 43686 12096
rect 44177 12087 44235 12093
rect 44177 12084 44189 12087
rect 43680 12056 44189 12084
rect 43680 12044 43686 12056
rect 44177 12053 44189 12056
rect 44223 12053 44235 12087
rect 44177 12047 44235 12053
rect 1104 11994 48852 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 48852 11994
rect 1104 11920 48852 11942
rect 18506 11880 18512 11892
rect 18467 11852 18512 11880
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 20165 11883 20223 11889
rect 20165 11880 20177 11883
rect 19024 11852 20177 11880
rect 19024 11840 19030 11852
rect 20165 11849 20177 11852
rect 20211 11849 20223 11883
rect 20530 11880 20536 11892
rect 20491 11852 20536 11880
rect 20165 11843 20223 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 23017 11883 23075 11889
rect 23017 11849 23029 11883
rect 23063 11880 23075 11883
rect 23198 11880 23204 11892
rect 23063 11852 23204 11880
rect 23063 11849 23075 11852
rect 23017 11843 23075 11849
rect 23198 11840 23204 11852
rect 23256 11840 23262 11892
rect 23382 11880 23388 11892
rect 23343 11852 23388 11880
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 26234 11880 26240 11892
rect 26195 11852 26240 11880
rect 26234 11840 26240 11852
rect 26292 11840 26298 11892
rect 26697 11883 26755 11889
rect 26697 11849 26709 11883
rect 26743 11880 26755 11883
rect 26786 11880 26792 11892
rect 26743 11852 26792 11880
rect 26743 11849 26755 11852
rect 26697 11843 26755 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 28166 11880 28172 11892
rect 28127 11852 28172 11880
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 29086 11880 29092 11892
rect 29047 11852 29092 11880
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 33686 11840 33692 11892
rect 33744 11880 33750 11892
rect 34149 11883 34207 11889
rect 34149 11880 34161 11883
rect 33744 11852 34161 11880
rect 33744 11840 33750 11852
rect 34149 11849 34161 11852
rect 34195 11849 34207 11883
rect 36078 11880 36084 11892
rect 36039 11852 36084 11880
rect 34149 11843 34207 11849
rect 36078 11840 36084 11852
rect 36136 11840 36142 11892
rect 36538 11840 36544 11892
rect 36596 11880 36602 11892
rect 36633 11883 36691 11889
rect 36633 11880 36645 11883
rect 36596 11852 36645 11880
rect 36596 11840 36602 11852
rect 36633 11849 36645 11852
rect 36679 11849 36691 11883
rect 36633 11843 36691 11849
rect 40313 11883 40371 11889
rect 40313 11849 40325 11883
rect 40359 11880 40371 11883
rect 40862 11880 40868 11892
rect 40359 11852 40868 11880
rect 40359 11849 40371 11852
rect 40313 11843 40371 11849
rect 40862 11840 40868 11852
rect 40920 11840 40926 11892
rect 42061 11883 42119 11889
rect 42061 11849 42073 11883
rect 42107 11880 42119 11883
rect 42242 11880 42248 11892
rect 42107 11852 42248 11880
rect 42107 11849 42119 11852
rect 42061 11843 42119 11849
rect 42242 11840 42248 11852
rect 42300 11840 42306 11892
rect 43254 11880 43260 11892
rect 43215 11852 43260 11880
rect 43254 11840 43260 11852
rect 43312 11840 43318 11892
rect 43438 11840 43444 11892
rect 43496 11880 43502 11892
rect 43533 11883 43591 11889
rect 43533 11880 43545 11883
rect 43496 11852 43545 11880
rect 43496 11840 43502 11852
rect 43533 11849 43545 11852
rect 43579 11849 43591 11883
rect 43533 11843 43591 11849
rect 45373 11883 45431 11889
rect 45373 11849 45385 11883
rect 45419 11880 45431 11883
rect 45462 11880 45468 11892
rect 45419 11852 45468 11880
rect 45419 11849 45431 11852
rect 45373 11843 45431 11849
rect 45462 11840 45468 11852
rect 45520 11840 45526 11892
rect 46566 11840 46572 11892
rect 46624 11880 46630 11892
rect 46845 11883 46903 11889
rect 46845 11880 46857 11883
rect 46624 11852 46857 11880
rect 46624 11840 46630 11852
rect 46845 11849 46857 11852
rect 46891 11849 46903 11883
rect 46845 11843 46903 11849
rect 19889 11815 19947 11821
rect 19889 11781 19901 11815
rect 19935 11812 19947 11815
rect 20622 11812 20628 11824
rect 19935 11784 20628 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 18922 11611 18980 11617
rect 18922 11577 18934 11611
rect 18968 11608 18980 11611
rect 19904 11608 19932 11775
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 23216 11812 23244 11840
rect 24949 11815 25007 11821
rect 24949 11812 24961 11815
rect 23216 11784 24961 11812
rect 24949 11781 24961 11784
rect 24995 11812 25007 11815
rect 25041 11815 25099 11821
rect 25041 11812 25053 11815
rect 24995 11784 25053 11812
rect 24995 11781 25007 11784
rect 24949 11775 25007 11781
rect 25041 11781 25053 11784
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 41693 11815 41751 11821
rect 41693 11781 41705 11815
rect 41739 11812 41751 11815
rect 42426 11812 42432 11824
rect 41739 11784 42432 11812
rect 41739 11781 41751 11784
rect 41693 11775 41751 11781
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 23753 11747 23811 11753
rect 21223 11716 22048 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 22020 11688 22048 11716
rect 23753 11713 23765 11747
rect 23799 11744 23811 11747
rect 23842 11744 23848 11756
rect 23799 11716 23848 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11744 24455 11747
rect 24486 11744 24492 11756
rect 24443 11716 24492 11744
rect 24443 11713 24455 11716
rect 24397 11707 24455 11713
rect 24486 11704 24492 11716
rect 24544 11704 24550 11756
rect 24670 11704 24676 11756
rect 24728 11744 24734 11756
rect 25961 11747 26019 11753
rect 25961 11744 25973 11747
rect 24728 11716 25973 11744
rect 24728 11704 24734 11716
rect 25961 11713 25973 11716
rect 26007 11744 26019 11747
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26007 11716 27169 11744
rect 26007 11713 26019 11716
rect 25961 11707 26019 11713
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 30006 11704 30012 11756
rect 30064 11744 30070 11756
rect 30285 11747 30343 11753
rect 30285 11744 30297 11747
rect 30064 11716 30297 11744
rect 30064 11704 30070 11716
rect 30285 11713 30297 11716
rect 30331 11713 30343 11747
rect 30285 11707 30343 11713
rect 37642 11704 37648 11756
rect 37700 11744 37706 11756
rect 42260 11753 42288 11784
rect 42426 11772 42432 11784
rect 42484 11772 42490 11824
rect 39945 11747 40003 11753
rect 37700 11716 39160 11744
rect 37700 11704 37706 11716
rect 20438 11685 20444 11688
rect 20416 11679 20444 11685
rect 20416 11676 20428 11679
rect 20351 11648 20428 11676
rect 20416 11645 20428 11648
rect 20496 11676 20502 11688
rect 21266 11676 21272 11688
rect 20496 11648 21272 11676
rect 20416 11639 20444 11645
rect 20438 11636 20444 11639
rect 20496 11636 20502 11648
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 21545 11679 21603 11685
rect 21545 11645 21557 11679
rect 21591 11676 21603 11679
rect 21818 11676 21824 11688
rect 21591 11648 21824 11676
rect 21591 11645 21603 11648
rect 21545 11639 21603 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 22002 11636 22008 11688
rect 22060 11676 22066 11688
rect 22097 11679 22155 11685
rect 22097 11676 22109 11679
rect 22060 11648 22109 11676
rect 22060 11636 22066 11648
rect 22097 11645 22109 11648
rect 22143 11645 22155 11679
rect 22097 11639 22155 11645
rect 27614 11636 27620 11688
rect 27672 11676 27678 11688
rect 28902 11676 28908 11688
rect 27672 11648 28908 11676
rect 27672 11636 27678 11648
rect 28902 11636 28908 11648
rect 28960 11676 28966 11688
rect 29733 11679 29791 11685
rect 29733 11676 29745 11679
rect 28960 11648 29745 11676
rect 28960 11636 28966 11648
rect 29733 11645 29745 11648
rect 29779 11645 29791 11679
rect 29733 11639 29791 11645
rect 31481 11679 31539 11685
rect 31481 11645 31493 11679
rect 31527 11676 31539 11679
rect 31757 11679 31815 11685
rect 31757 11676 31769 11679
rect 31527 11648 31769 11676
rect 31527 11645 31539 11648
rect 31481 11639 31539 11645
rect 31757 11645 31769 11648
rect 31803 11676 31815 11679
rect 32582 11676 32588 11688
rect 31803 11648 32588 11676
rect 31803 11645 31815 11648
rect 31757 11639 31815 11645
rect 32582 11636 32588 11648
rect 32640 11676 32646 11688
rect 33042 11676 33048 11688
rect 32640 11648 33048 11676
rect 32640 11636 32646 11648
rect 33042 11636 33048 11648
rect 33100 11676 33106 11688
rect 33137 11679 33195 11685
rect 33137 11676 33149 11679
rect 33100 11648 33149 11676
rect 33100 11636 33106 11648
rect 33137 11645 33149 11648
rect 33183 11676 33195 11679
rect 33781 11679 33839 11685
rect 33781 11676 33793 11679
rect 33183 11648 33793 11676
rect 33183 11645 33195 11648
rect 33137 11639 33195 11645
rect 33781 11645 33793 11648
rect 33827 11645 33839 11679
rect 33781 11639 33839 11645
rect 35253 11679 35311 11685
rect 35253 11645 35265 11679
rect 35299 11645 35311 11679
rect 35526 11676 35532 11688
rect 35487 11648 35532 11676
rect 35253 11639 35311 11645
rect 18968 11580 19932 11608
rect 18968 11577 18980 11580
rect 18922 11571 18980 11577
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 23845 11611 23903 11617
rect 23440 11580 23520 11608
rect 23440 11568 23446 11580
rect 17221 11543 17279 11549
rect 17221 11509 17233 11543
rect 17267 11540 17279 11543
rect 17402 11540 17408 11552
rect 17267 11512 17408 11540
rect 17267 11509 17279 11512
rect 17221 11503 17279 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 19521 11543 19579 11549
rect 19521 11540 19533 11543
rect 19484 11512 19533 11540
rect 19484 11500 19490 11512
rect 19521 11509 19533 11512
rect 19567 11509 19579 11543
rect 21726 11540 21732 11552
rect 21687 11512 21732 11540
rect 19521 11503 19579 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 23492 11540 23520 11580
rect 23845 11577 23857 11611
rect 23891 11577 23903 11611
rect 25314 11608 25320 11620
rect 25275 11580 25320 11608
rect 23845 11571 23903 11577
rect 23860 11540 23888 11571
rect 25314 11568 25320 11580
rect 25372 11568 25378 11620
rect 25409 11611 25467 11617
rect 25409 11577 25421 11611
rect 25455 11577 25467 11611
rect 25409 11571 25467 11577
rect 26881 11611 26939 11617
rect 26881 11577 26893 11611
rect 26927 11577 26939 11611
rect 26881 11571 26939 11577
rect 23492 11512 23888 11540
rect 24486 11500 24492 11552
rect 24544 11540 24550 11552
rect 24673 11543 24731 11549
rect 24673 11540 24685 11543
rect 24544 11512 24685 11540
rect 24544 11500 24550 11512
rect 24673 11509 24685 11512
rect 24719 11509 24731 11543
rect 24673 11503 24731 11509
rect 24949 11543 25007 11549
rect 24949 11509 24961 11543
rect 24995 11540 25007 11543
rect 25424 11540 25452 11571
rect 26694 11540 26700 11552
rect 24995 11512 26700 11540
rect 24995 11509 25007 11512
rect 24949 11503 25007 11509
rect 26694 11500 26700 11512
rect 26752 11500 26758 11552
rect 26786 11500 26792 11552
rect 26844 11540 26850 11552
rect 26896 11540 26924 11571
rect 26970 11568 26976 11620
rect 27028 11608 27034 11620
rect 27801 11611 27859 11617
rect 27801 11608 27813 11611
rect 27028 11580 27813 11608
rect 27028 11568 27034 11580
rect 27801 11577 27813 11580
rect 27847 11608 27859 11611
rect 29822 11608 29828 11620
rect 27847 11580 29828 11608
rect 27847 11577 27859 11580
rect 27801 11571 27859 11577
rect 29822 11568 29828 11580
rect 29880 11568 29886 11620
rect 30009 11611 30067 11617
rect 30009 11577 30021 11611
rect 30055 11577 30067 11611
rect 30009 11571 30067 11577
rect 26844 11512 26924 11540
rect 26844 11500 26850 11512
rect 28442 11500 28448 11552
rect 28500 11540 28506 11552
rect 28629 11543 28687 11549
rect 28629 11540 28641 11543
rect 28500 11512 28641 11540
rect 28500 11500 28506 11512
rect 28629 11509 28641 11512
rect 28675 11509 28687 11543
rect 30024 11540 30052 11571
rect 30098 11568 30104 11620
rect 30156 11608 30162 11620
rect 31570 11608 31576 11620
rect 30156 11580 30201 11608
rect 31531 11580 31576 11608
rect 30156 11568 30162 11580
rect 31570 11568 31576 11580
rect 31628 11568 31634 11620
rect 32125 11611 32183 11617
rect 32125 11577 32137 11611
rect 32171 11608 32183 11611
rect 32674 11608 32680 11620
rect 32171 11580 32680 11608
rect 32171 11577 32183 11580
rect 32125 11571 32183 11577
rect 32674 11568 32680 11580
rect 32732 11568 32738 11620
rect 32953 11611 33011 11617
rect 32953 11577 32965 11611
rect 32999 11608 33011 11611
rect 33318 11608 33324 11620
rect 32999 11580 33324 11608
rect 32999 11577 33011 11580
rect 32953 11571 33011 11577
rect 33318 11568 33324 11580
rect 33376 11568 33382 11620
rect 33502 11608 33508 11620
rect 33463 11580 33508 11608
rect 33502 11568 33508 11580
rect 33560 11568 33566 11620
rect 30834 11540 30840 11552
rect 30024 11512 30840 11540
rect 28629 11503 28687 11509
rect 30834 11500 30840 11512
rect 30892 11540 30898 11552
rect 30929 11543 30987 11549
rect 30929 11540 30941 11543
rect 30892 11512 30941 11540
rect 30892 11500 30898 11512
rect 30929 11509 30941 11512
rect 30975 11509 30987 11543
rect 30929 11503 30987 11509
rect 34701 11543 34759 11549
rect 34701 11509 34713 11543
rect 34747 11540 34759 11543
rect 35268 11540 35296 11639
rect 35526 11636 35532 11648
rect 35584 11636 35590 11688
rect 36722 11636 36728 11688
rect 36780 11676 36786 11688
rect 37752 11685 37780 11716
rect 39132 11688 39160 11716
rect 39945 11713 39957 11747
rect 39991 11744 40003 11747
rect 42245 11747 42303 11753
rect 39991 11716 41000 11744
rect 39991 11713 40003 11716
rect 39945 11707 40003 11713
rect 37093 11679 37151 11685
rect 37093 11676 37105 11679
rect 36780 11648 37105 11676
rect 36780 11636 36786 11648
rect 37093 11645 37105 11648
rect 37139 11676 37151 11679
rect 37461 11679 37519 11685
rect 37461 11676 37473 11679
rect 37139 11648 37473 11676
rect 37139 11645 37151 11648
rect 37093 11639 37151 11645
rect 37461 11645 37473 11648
rect 37507 11676 37519 11679
rect 37737 11679 37795 11685
rect 37507 11648 37596 11676
rect 37507 11645 37519 11648
rect 37461 11639 37519 11645
rect 35710 11608 35716 11620
rect 35671 11580 35716 11608
rect 35710 11568 35716 11580
rect 35768 11568 35774 11620
rect 35894 11540 35900 11552
rect 34747 11512 35900 11540
rect 34747 11509 34759 11512
rect 34701 11503 34759 11509
rect 35894 11500 35900 11512
rect 35952 11500 35958 11552
rect 37568 11540 37596 11648
rect 37737 11645 37749 11679
rect 37783 11645 37795 11679
rect 38841 11679 38899 11685
rect 38841 11676 38853 11679
rect 37737 11639 37795 11645
rect 38672 11648 38853 11676
rect 37918 11608 37924 11620
rect 37879 11580 37924 11608
rect 37918 11568 37924 11580
rect 37976 11568 37982 11620
rect 37826 11540 37832 11552
rect 37568 11512 37832 11540
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 38010 11500 38016 11552
rect 38068 11540 38074 11552
rect 38197 11543 38255 11549
rect 38197 11540 38209 11543
rect 38068 11512 38209 11540
rect 38068 11500 38074 11512
rect 38197 11509 38209 11512
rect 38243 11509 38255 11543
rect 38197 11503 38255 11509
rect 38562 11500 38568 11552
rect 38620 11540 38626 11552
rect 38672 11549 38700 11648
rect 38841 11645 38853 11648
rect 38887 11676 38899 11679
rect 38930 11676 38936 11688
rect 38887 11648 38936 11676
rect 38887 11645 38899 11648
rect 38841 11639 38899 11645
rect 38930 11636 38936 11648
rect 38988 11636 38994 11688
rect 39114 11636 39120 11688
rect 39172 11676 39178 11688
rect 39393 11679 39451 11685
rect 39393 11676 39405 11679
rect 39172 11648 39405 11676
rect 39172 11636 39178 11648
rect 39393 11645 39405 11648
rect 39439 11676 39451 11679
rect 39960 11676 39988 11707
rect 40972 11688 41000 11716
rect 42245 11713 42257 11747
rect 42291 11713 42303 11747
rect 42245 11707 42303 11713
rect 42334 11704 42340 11756
rect 42392 11744 42398 11756
rect 42521 11747 42579 11753
rect 42521 11744 42533 11747
rect 42392 11716 42533 11744
rect 42392 11704 42398 11716
rect 42521 11713 42533 11716
rect 42567 11713 42579 11747
rect 42521 11707 42579 11713
rect 40494 11676 40500 11688
rect 39439 11648 39988 11676
rect 40455 11648 40500 11676
rect 39439 11645 39451 11648
rect 39393 11639 39451 11645
rect 40494 11636 40500 11648
rect 40552 11636 40558 11688
rect 40954 11676 40960 11688
rect 40915 11648 40960 11676
rect 40954 11636 40960 11648
rect 41012 11636 41018 11688
rect 39574 11608 39580 11620
rect 39535 11580 39580 11608
rect 39574 11568 39580 11580
rect 39632 11568 39638 11620
rect 42242 11568 42248 11620
rect 42300 11608 42306 11620
rect 42337 11611 42395 11617
rect 42337 11608 42349 11611
rect 42300 11580 42349 11608
rect 42300 11568 42306 11580
rect 42337 11577 42349 11580
rect 42383 11577 42395 11611
rect 42337 11571 42395 11577
rect 43622 11568 43628 11620
rect 43680 11608 43686 11620
rect 43809 11611 43867 11617
rect 43809 11608 43821 11611
rect 43680 11580 43821 11608
rect 43680 11568 43686 11580
rect 43809 11577 43821 11580
rect 43855 11577 43867 11611
rect 43809 11571 43867 11577
rect 43901 11611 43959 11617
rect 43901 11577 43913 11611
rect 43947 11577 43959 11611
rect 44450 11608 44456 11620
rect 44411 11580 44456 11608
rect 43901 11571 43959 11577
rect 38657 11543 38715 11549
rect 38657 11540 38669 11543
rect 38620 11512 38669 11540
rect 38620 11500 38626 11512
rect 38657 11509 38669 11512
rect 38703 11509 38715 11543
rect 40586 11540 40592 11552
rect 40547 11512 40592 11540
rect 38657 11503 38715 11509
rect 40586 11500 40592 11512
rect 40644 11500 40650 11552
rect 42058 11500 42064 11552
rect 42116 11540 42122 11552
rect 43254 11540 43260 11552
rect 42116 11512 43260 11540
rect 42116 11500 42122 11512
rect 43254 11500 43260 11512
rect 43312 11500 43318 11552
rect 43438 11500 43444 11552
rect 43496 11540 43502 11552
rect 43916 11540 43944 11571
rect 44450 11568 44456 11580
rect 44508 11568 44514 11620
rect 44542 11568 44548 11620
rect 44600 11608 44606 11620
rect 45370 11608 45376 11620
rect 44600 11580 45376 11608
rect 44600 11568 44606 11580
rect 45370 11568 45376 11580
rect 45428 11608 45434 11620
rect 45649 11611 45707 11617
rect 45649 11608 45661 11611
rect 45428 11580 45661 11608
rect 45428 11568 45434 11580
rect 45649 11577 45661 11580
rect 45695 11577 45707 11611
rect 45649 11571 45707 11577
rect 43990 11540 43996 11552
rect 43496 11512 43996 11540
rect 43496 11500 43502 11512
rect 43990 11500 43996 11512
rect 44048 11500 44054 11552
rect 1104 11450 48852 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 48852 11450
rect 1104 11376 48852 11398
rect 18598 11336 18604 11348
rect 18559 11308 18604 11336
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 20438 11336 20444 11348
rect 20399 11308 20444 11336
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21453 11339 21511 11345
rect 21453 11336 21465 11339
rect 21140 11308 21465 11336
rect 21140 11296 21146 11308
rect 21453 11305 21465 11308
rect 21499 11305 21511 11339
rect 23014 11336 23020 11348
rect 22975 11308 23020 11336
rect 21453 11299 21511 11305
rect 23014 11296 23020 11308
rect 23072 11336 23078 11348
rect 23523 11339 23581 11345
rect 23523 11336 23535 11339
rect 23072 11308 23535 11336
rect 23072 11296 23078 11308
rect 23523 11305 23535 11308
rect 23569 11305 23581 11339
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 23523 11299 23581 11305
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 28718 11336 28724 11348
rect 28679 11308 28724 11336
rect 28718 11296 28724 11308
rect 28776 11296 28782 11348
rect 29822 11296 29828 11348
rect 29880 11336 29886 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 29880 11308 29929 11336
rect 29880 11296 29886 11308
rect 29917 11305 29929 11308
rect 29963 11336 29975 11339
rect 30098 11336 30104 11348
rect 29963 11308 30104 11336
rect 29963 11305 29975 11308
rect 29917 11299 29975 11305
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 31570 11336 31576 11348
rect 31531 11308 31576 11336
rect 31570 11296 31576 11308
rect 31628 11296 31634 11348
rect 32490 11336 32496 11348
rect 32451 11308 32496 11336
rect 32490 11296 32496 11308
rect 32548 11296 32554 11348
rect 33594 11336 33600 11348
rect 32876 11308 33600 11336
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 19208 11240 19257 11268
rect 19208 11228 19214 11240
rect 19245 11237 19257 11240
rect 19291 11268 19303 11271
rect 19886 11268 19892 11280
rect 19291 11240 19892 11268
rect 19291 11237 19303 11240
rect 19245 11231 19303 11237
rect 19886 11228 19892 11240
rect 19944 11228 19950 11280
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18084 11203 18142 11209
rect 18084 11200 18096 11203
rect 17920 11172 18096 11200
rect 17920 11160 17926 11172
rect 18084 11169 18096 11172
rect 18130 11169 18142 11203
rect 18084 11163 18142 11169
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11200 19855 11203
rect 20070 11200 20076 11212
rect 19843 11172 20076 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 20070 11160 20076 11172
rect 20128 11200 20134 11212
rect 20456 11200 20484 11296
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 21266 11268 21272 11280
rect 20680 11240 21272 11268
rect 20680 11228 20686 11240
rect 21266 11228 21272 11240
rect 21324 11268 21330 11280
rect 21958 11271 22016 11277
rect 21958 11268 21970 11271
rect 21324 11240 21970 11268
rect 21324 11228 21330 11240
rect 21958 11237 21970 11240
rect 22004 11237 22016 11271
rect 21958 11231 22016 11237
rect 26694 11228 26700 11280
rect 26752 11268 26758 11280
rect 27249 11271 27307 11277
rect 27249 11268 27261 11271
rect 26752 11240 27261 11268
rect 26752 11228 26758 11240
rect 27249 11237 27261 11240
rect 27295 11268 27307 11271
rect 27614 11268 27620 11280
rect 27295 11240 27620 11268
rect 27295 11237 27307 11240
rect 27249 11231 27307 11237
rect 27614 11228 27620 11240
rect 27672 11228 27678 11280
rect 27798 11268 27804 11280
rect 27759 11240 27804 11268
rect 27798 11228 27804 11240
rect 27856 11228 27862 11280
rect 31588 11268 31616 11296
rect 32876 11277 32904 11308
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 33870 11336 33876 11348
rect 33831 11308 33876 11336
rect 33870 11296 33876 11308
rect 33928 11296 33934 11348
rect 36722 11336 36728 11348
rect 36683 11308 36728 11336
rect 36722 11296 36728 11308
rect 36780 11296 36786 11348
rect 37277 11339 37335 11345
rect 37277 11305 37289 11339
rect 37323 11336 37335 11339
rect 37642 11336 37648 11348
rect 37323 11308 37648 11336
rect 37323 11305 37335 11308
rect 37277 11299 37335 11305
rect 37642 11296 37648 11308
rect 37700 11296 37706 11348
rect 37918 11336 37924 11348
rect 37879 11308 37924 11336
rect 37918 11296 37924 11308
rect 37976 11296 37982 11348
rect 40221 11339 40279 11345
rect 40221 11305 40233 11339
rect 40267 11336 40279 11339
rect 40586 11336 40592 11348
rect 40267 11308 40592 11336
rect 40267 11305 40279 11308
rect 40221 11299 40279 11305
rect 40586 11296 40592 11308
rect 40644 11296 40650 11348
rect 42150 11336 42156 11348
rect 42111 11308 42156 11336
rect 42150 11296 42156 11308
rect 42208 11296 42214 11348
rect 32861 11271 32919 11277
rect 32861 11268 32873 11271
rect 31588 11240 32873 11268
rect 32861 11237 32873 11240
rect 32907 11237 32919 11271
rect 32861 11231 32919 11237
rect 33413 11271 33471 11277
rect 33413 11237 33425 11271
rect 33459 11268 33471 11271
rect 38746 11268 38752 11280
rect 33459 11240 36584 11268
rect 38707 11240 38752 11268
rect 33459 11237 33471 11240
rect 33413 11231 33471 11237
rect 20128 11172 20484 11200
rect 20128 11160 20134 11172
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21085 11203 21143 11209
rect 21085 11200 21097 11203
rect 21048 11172 21097 11200
rect 21048 11160 21054 11172
rect 21085 11169 21097 11172
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 22557 11203 22615 11209
rect 22557 11169 22569 11203
rect 22603 11200 22615 11203
rect 23382 11200 23388 11212
rect 23440 11209 23446 11212
rect 23440 11203 23478 11209
rect 22603 11172 23388 11200
rect 22603 11169 22615 11172
rect 22557 11163 22615 11169
rect 23382 11160 23388 11172
rect 23466 11169 23478 11203
rect 28626 11200 28632 11212
rect 28587 11172 28632 11200
rect 23440 11163 23478 11169
rect 23440 11160 23446 11163
rect 28626 11160 28632 11172
rect 28684 11160 28690 11212
rect 29181 11203 29239 11209
rect 29181 11169 29193 11203
rect 29227 11200 29239 11203
rect 29270 11200 29276 11212
rect 29227 11172 29276 11200
rect 29227 11169 29239 11172
rect 29181 11163 29239 11169
rect 29270 11160 29276 11172
rect 29328 11160 29334 11212
rect 30466 11200 30472 11212
rect 30427 11172 30472 11200
rect 30466 11160 30472 11172
rect 30524 11160 30530 11212
rect 30653 11203 30711 11209
rect 30653 11169 30665 11203
rect 30699 11169 30711 11203
rect 30653 11163 30711 11169
rect 33045 11203 33103 11209
rect 33045 11169 33057 11203
rect 33091 11200 33103 11203
rect 33870 11200 33876 11212
rect 33091 11172 33876 11200
rect 33091 11169 33103 11172
rect 33045 11163 33103 11169
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 19024 11104 19165 11132
rect 19024 11092 19030 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 21634 11132 21640 11144
rect 21595 11104 21640 11132
rect 19153 11095 19211 11101
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 24578 11132 24584 11144
rect 24539 11104 24584 11132
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 27157 11135 27215 11141
rect 27157 11101 27169 11135
rect 27203 11132 27215 11135
rect 27430 11132 27436 11144
rect 27203 11104 27436 11132
rect 27203 11101 27215 11104
rect 27157 11095 27215 11101
rect 27430 11092 27436 11104
rect 27488 11092 27494 11144
rect 29288 11132 29316 11160
rect 30006 11132 30012 11144
rect 29288 11104 30012 11132
rect 30006 11092 30012 11104
rect 30064 11132 30070 11144
rect 30668 11132 30696 11163
rect 33870 11160 33876 11172
rect 33928 11160 33934 11212
rect 34606 11160 34612 11212
rect 34664 11200 34670 11212
rect 34977 11203 35035 11209
rect 34977 11200 34989 11203
rect 34664 11172 34989 11200
rect 34664 11160 34670 11172
rect 34977 11169 34989 11172
rect 35023 11169 35035 11203
rect 35526 11200 35532 11212
rect 35487 11172 35532 11200
rect 34977 11163 35035 11169
rect 35526 11160 35532 11172
rect 35584 11160 35590 11212
rect 36556 11209 36584 11240
rect 38746 11228 38752 11240
rect 38804 11228 38810 11280
rect 40862 11228 40868 11280
rect 40920 11268 40926 11280
rect 41002 11271 41060 11277
rect 41002 11268 41014 11271
rect 40920 11240 41014 11268
rect 40920 11228 40926 11240
rect 41002 11237 41014 11240
rect 41048 11237 41060 11271
rect 43990 11268 43996 11280
rect 43951 11240 43996 11268
rect 41002 11231 41060 11237
rect 43990 11228 43996 11240
rect 44048 11228 44054 11280
rect 36541 11203 36599 11209
rect 36541 11169 36553 11203
rect 36587 11200 36599 11203
rect 37274 11200 37280 11212
rect 36587 11172 37280 11200
rect 36587 11169 36599 11172
rect 36541 11163 36599 11169
rect 37274 11160 37280 11172
rect 37332 11160 37338 11212
rect 45186 11160 45192 11212
rect 45244 11200 45250 11212
rect 45500 11203 45558 11209
rect 45500 11200 45512 11203
rect 45244 11172 45512 11200
rect 45244 11160 45250 11172
rect 45500 11169 45512 11172
rect 45546 11169 45558 11203
rect 45500 11163 45558 11169
rect 30926 11132 30932 11144
rect 30064 11104 30696 11132
rect 30887 11104 30932 11132
rect 30064 11092 30070 11104
rect 30926 11092 30932 11104
rect 30984 11092 30990 11144
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11132 35771 11135
rect 37826 11132 37832 11144
rect 35759 11104 37832 11132
rect 35759 11101 35771 11104
rect 35713 11095 35771 11101
rect 37826 11092 37832 11104
rect 37884 11092 37890 11144
rect 38657 11135 38715 11141
rect 38657 11101 38669 11135
rect 38703 11132 38715 11135
rect 39482 11132 39488 11144
rect 38703 11104 39488 11132
rect 38703 11101 38715 11104
rect 38657 11095 38715 11101
rect 39482 11092 39488 11104
rect 39540 11092 39546 11144
rect 39942 11092 39948 11144
rect 40000 11132 40006 11144
rect 40681 11135 40739 11141
rect 40681 11132 40693 11135
rect 40000 11104 40693 11132
rect 40000 11092 40006 11104
rect 40681 11101 40693 11104
rect 40727 11101 40739 11135
rect 43898 11132 43904 11144
rect 43859 11104 43904 11132
rect 40681 11095 40739 11101
rect 43898 11092 43904 11104
rect 43956 11092 43962 11144
rect 44542 11132 44548 11144
rect 44503 11104 44548 11132
rect 44542 11092 44548 11104
rect 44600 11092 44606 11144
rect 39209 11067 39267 11073
rect 39209 11033 39221 11067
rect 39255 11064 39267 11067
rect 39298 11064 39304 11076
rect 39255 11036 39304 11064
rect 39255 11033 39267 11036
rect 39209 11027 39267 11033
rect 39298 11024 39304 11036
rect 39356 11024 39362 11076
rect 18187 10999 18245 11005
rect 18187 10965 18199 10999
rect 18233 10996 18245 10999
rect 19518 10996 19524 11008
rect 18233 10968 19524 10996
rect 18233 10965 18245 10968
rect 18187 10959 18245 10965
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 23842 10996 23848 11008
rect 23803 10968 23848 10996
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 25498 10996 25504 11008
rect 25459 10968 25504 10996
rect 25498 10956 25504 10968
rect 25556 10956 25562 11008
rect 26786 10996 26792 11008
rect 26747 10968 26792 10996
rect 26786 10956 26792 10968
rect 26844 10956 26850 11008
rect 27522 10956 27528 11008
rect 27580 10996 27586 11008
rect 28077 10999 28135 11005
rect 28077 10996 28089 10999
rect 27580 10968 28089 10996
rect 27580 10956 27586 10968
rect 28077 10965 28089 10968
rect 28123 10965 28135 10999
rect 28077 10959 28135 10965
rect 37734 10956 37740 11008
rect 37792 10996 37798 11008
rect 40494 10996 40500 11008
rect 37792 10968 40500 10996
rect 37792 10956 37798 10968
rect 40494 10956 40500 10968
rect 40552 10956 40558 11008
rect 41598 10996 41604 11008
rect 41559 10968 41604 10996
rect 41598 10956 41604 10968
rect 41656 10956 41662 11008
rect 45603 10999 45661 11005
rect 45603 10965 45615 10999
rect 45649 10996 45661 10999
rect 46014 10996 46020 11008
rect 45649 10968 46020 10996
rect 45649 10965 45661 10968
rect 45603 10959 45661 10965
rect 46014 10956 46020 10968
rect 46072 10956 46078 11008
rect 1104 10906 48852 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 48852 10906
rect 1104 10832 48852 10854
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 16172 10764 16221 10792
rect 16172 10752 16178 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16209 10755 16267 10761
rect 17083 10795 17141 10801
rect 17083 10761 17095 10795
rect 17129 10792 17141 10795
rect 18966 10792 18972 10804
rect 17129 10764 18972 10792
rect 17129 10761 17141 10764
rect 17083 10755 17141 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 19150 10792 19156 10804
rect 19111 10764 19156 10792
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 19260 10764 20821 10792
rect 16761 10727 16819 10733
rect 16761 10693 16773 10727
rect 16807 10724 16819 10727
rect 17770 10724 17776 10736
rect 16807 10696 17776 10724
rect 16807 10693 16819 10696
rect 16761 10687 16819 10693
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16776 10588 16804 10687
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18984 10724 19012 10752
rect 19260 10724 19288 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 20809 10755 20867 10761
rect 21266 10752 21272 10764
rect 21324 10792 21330 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 21324 10764 21557 10792
rect 21324 10752 21330 10764
rect 21545 10761 21557 10764
rect 21591 10761 21603 10795
rect 23382 10792 23388 10804
rect 23343 10764 23388 10792
rect 21545 10755 21603 10761
rect 20070 10724 20076 10736
rect 18984 10696 19288 10724
rect 20031 10696 20076 10724
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 16439 10560 16804 10588
rect 16868 10628 17877 10656
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16298 10480 16304 10532
rect 16356 10520 16362 10532
rect 16868 10520 16896 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 19518 10656 19524 10668
rect 19479 10628 19524 10656
rect 17865 10619 17923 10625
rect 17012 10591 17070 10597
rect 17012 10557 17024 10591
rect 17058 10588 17070 10591
rect 17880 10588 17908 10619
rect 19518 10616 19524 10628
rect 19576 10656 19582 10668
rect 19978 10656 19984 10668
rect 19576 10628 19984 10656
rect 19576 10616 19582 10628
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 18452 10591 18510 10597
rect 18452 10588 18464 10591
rect 17058 10560 17540 10588
rect 17880 10560 18464 10588
rect 17058 10557 17070 10560
rect 17012 10551 17070 10557
rect 16356 10492 16896 10520
rect 16356 10480 16362 10492
rect 17512 10464 17540 10560
rect 18452 10557 18464 10560
rect 18498 10557 18510 10591
rect 18452 10551 18510 10557
rect 19613 10523 19671 10529
rect 19613 10489 19625 10523
rect 19659 10489 19671 10523
rect 21560 10520 21588 10755
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 25314 10752 25320 10804
rect 25372 10792 25378 10804
rect 26467 10795 26525 10801
rect 26467 10792 26479 10795
rect 25372 10764 26479 10792
rect 25372 10752 25378 10764
rect 26467 10761 26479 10764
rect 26513 10761 26525 10795
rect 26467 10755 26525 10761
rect 26694 10752 26700 10804
rect 26752 10792 26758 10804
rect 26881 10795 26939 10801
rect 26881 10792 26893 10795
rect 26752 10764 26893 10792
rect 26752 10752 26758 10764
rect 26881 10761 26893 10764
rect 26927 10761 26939 10795
rect 26881 10755 26939 10761
rect 28994 10752 29000 10804
rect 29052 10792 29058 10804
rect 29089 10795 29147 10801
rect 29089 10792 29101 10795
rect 29052 10764 29101 10792
rect 29052 10752 29058 10764
rect 29089 10761 29101 10764
rect 29135 10792 29147 10795
rect 29270 10792 29276 10804
rect 29135 10764 29276 10792
rect 29135 10761 29147 10764
rect 29089 10755 29147 10761
rect 29270 10752 29276 10764
rect 29328 10752 29334 10804
rect 31294 10792 31300 10804
rect 31255 10764 31300 10792
rect 31294 10752 31300 10764
rect 31352 10752 31358 10804
rect 33413 10795 33471 10801
rect 33413 10761 33425 10795
rect 33459 10792 33471 10795
rect 33594 10792 33600 10804
rect 33459 10764 33600 10792
rect 33459 10761 33471 10764
rect 33413 10755 33471 10761
rect 33594 10752 33600 10764
rect 33652 10752 33658 10804
rect 33781 10795 33839 10801
rect 33781 10761 33793 10795
rect 33827 10792 33839 10795
rect 33870 10792 33876 10804
rect 33827 10764 33876 10792
rect 33827 10761 33839 10764
rect 33781 10755 33839 10761
rect 33870 10752 33876 10764
rect 33928 10752 33934 10804
rect 37274 10792 37280 10804
rect 37235 10764 37280 10792
rect 37274 10752 37280 10764
rect 37332 10752 37338 10804
rect 39850 10752 39856 10804
rect 39908 10792 39914 10804
rect 40313 10795 40371 10801
rect 40313 10792 40325 10795
rect 39908 10764 40325 10792
rect 39908 10752 39914 10764
rect 40313 10761 40325 10764
rect 40359 10792 40371 10795
rect 40773 10795 40831 10801
rect 40773 10792 40785 10795
rect 40359 10764 40785 10792
rect 40359 10761 40371 10764
rect 40313 10755 40371 10761
rect 40773 10761 40785 10764
rect 40819 10792 40831 10795
rect 40862 10792 40868 10804
rect 40819 10764 40868 10792
rect 40819 10761 40831 10764
rect 40773 10755 40831 10761
rect 40862 10752 40868 10764
rect 40920 10752 40926 10804
rect 41598 10752 41604 10804
rect 41656 10792 41662 10804
rect 42429 10795 42487 10801
rect 42429 10792 42441 10795
rect 41656 10764 42441 10792
rect 41656 10752 41662 10764
rect 42429 10761 42441 10764
rect 42475 10761 42487 10795
rect 42429 10755 42487 10761
rect 43441 10795 43499 10801
rect 43441 10761 43453 10795
rect 43487 10792 43499 10795
rect 43714 10792 43720 10804
rect 43487 10764 43720 10792
rect 43487 10761 43499 10764
rect 43441 10755 43499 10761
rect 29549 10727 29607 10733
rect 29549 10693 29561 10727
rect 29595 10724 29607 10727
rect 30466 10724 30472 10736
rect 29595 10696 30472 10724
rect 29595 10693 29607 10696
rect 29549 10687 29607 10693
rect 30466 10684 30472 10696
rect 30524 10684 30530 10736
rect 35069 10727 35127 10733
rect 35069 10693 35081 10727
rect 35115 10693 35127 10727
rect 35069 10687 35127 10693
rect 41785 10727 41843 10733
rect 41785 10693 41797 10727
rect 41831 10724 41843 10727
rect 42058 10724 42064 10736
rect 41831 10696 42064 10724
rect 41831 10693 41843 10696
rect 41785 10687 41843 10693
rect 21726 10656 21732 10668
rect 21687 10628 21732 10656
rect 21726 10616 21732 10628
rect 21784 10616 21790 10668
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 24762 10656 24768 10668
rect 24627 10628 24768 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 32125 10659 32183 10665
rect 32125 10656 32137 10659
rect 30984 10628 32137 10656
rect 30984 10616 30990 10628
rect 32125 10625 32137 10628
rect 32171 10656 32183 10659
rect 32306 10656 32312 10668
rect 32171 10628 32312 10656
rect 32171 10625 32183 10628
rect 32125 10619 32183 10625
rect 32306 10616 32312 10628
rect 32364 10616 32370 10668
rect 34606 10656 34612 10668
rect 34567 10628 34612 10656
rect 34606 10616 34612 10628
rect 34664 10656 34670 10668
rect 35084 10656 35112 10687
rect 42058 10684 42064 10696
rect 42116 10684 42122 10736
rect 34664 10628 35112 10656
rect 34664 10616 34670 10628
rect 35710 10616 35716 10668
rect 35768 10656 35774 10668
rect 36078 10656 36084 10668
rect 35768 10628 36084 10656
rect 35768 10616 35774 10628
rect 36078 10616 36084 10628
rect 36136 10616 36142 10668
rect 37826 10656 37832 10668
rect 37787 10628 37832 10656
rect 37826 10616 37832 10628
rect 37884 10616 37890 10668
rect 39574 10616 39580 10668
rect 39632 10656 39638 10668
rect 40865 10659 40923 10665
rect 40865 10656 40877 10659
rect 39632 10628 40877 10656
rect 39632 10616 39638 10628
rect 40865 10625 40877 10628
rect 40911 10656 40923 10659
rect 41138 10656 41144 10668
rect 40911 10628 41144 10656
rect 40911 10625 40923 10628
rect 40865 10619 40923 10625
rect 41138 10616 41144 10628
rect 41196 10616 41202 10668
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 22925 10591 22983 10597
rect 22925 10588 22937 10591
rect 21692 10560 22937 10588
rect 21692 10548 21698 10560
rect 22925 10557 22937 10560
rect 22971 10557 22983 10591
rect 22925 10551 22983 10557
rect 25501 10591 25559 10597
rect 25501 10557 25513 10591
rect 25547 10588 25559 10591
rect 26145 10591 26203 10597
rect 26145 10588 26157 10591
rect 25547 10560 26157 10588
rect 25547 10557 25559 10560
rect 25501 10551 25559 10557
rect 26145 10557 26157 10560
rect 26191 10588 26203 10591
rect 26364 10591 26422 10597
rect 26364 10588 26376 10591
rect 26191 10560 26376 10588
rect 26191 10557 26203 10560
rect 26145 10551 26203 10557
rect 26364 10557 26376 10560
rect 26410 10557 26422 10591
rect 26364 10551 26422 10557
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10588 27491 10591
rect 27522 10588 27528 10600
rect 27479 10560 27528 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 27522 10548 27528 10560
rect 27580 10548 27586 10600
rect 29365 10591 29423 10597
rect 29365 10557 29377 10591
rect 29411 10588 29423 10591
rect 30374 10588 30380 10600
rect 29411 10560 29960 10588
rect 30335 10560 30380 10588
rect 29411 10557 29423 10560
rect 29365 10551 29423 10557
rect 22050 10523 22108 10529
rect 22050 10520 22062 10523
rect 21560 10492 22062 10520
rect 19613 10483 19671 10489
rect 22050 10489 22062 10492
rect 22096 10520 22108 10523
rect 23566 10520 23572 10532
rect 22096 10492 23572 10520
rect 22096 10489 22108 10492
rect 22050 10483 22108 10489
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 17920 10424 18245 10452
rect 17920 10412 17926 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18233 10415 18291 10421
rect 18555 10455 18613 10461
rect 18555 10421 18567 10455
rect 18601 10452 18613 10455
rect 18782 10452 18788 10464
rect 18601 10424 18788 10452
rect 18601 10421 18613 10424
rect 18555 10415 18613 10421
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19628 10452 19656 10483
rect 23566 10480 23572 10492
rect 23624 10520 23630 10532
rect 24946 10529 24952 10532
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 23624 10492 24041 10520
rect 23624 10480 23630 10492
rect 24029 10489 24041 10492
rect 24075 10520 24087 10523
rect 24397 10523 24455 10529
rect 24397 10520 24409 10523
rect 24075 10492 24409 10520
rect 24075 10489 24087 10492
rect 24029 10483 24087 10489
rect 24397 10489 24409 10492
rect 24443 10520 24455 10523
rect 24902 10523 24952 10529
rect 24902 10520 24914 10523
rect 24443 10492 24914 10520
rect 24443 10489 24455 10492
rect 24397 10483 24455 10489
rect 24902 10489 24914 10492
rect 24948 10489 24952 10523
rect 24902 10483 24952 10489
rect 24946 10480 24952 10483
rect 25004 10520 25010 10532
rect 27062 10520 27068 10532
rect 25004 10492 27068 10520
rect 25004 10480 25010 10492
rect 27062 10480 27068 10492
rect 27120 10520 27126 10532
rect 27249 10523 27307 10529
rect 27249 10520 27261 10523
rect 27120 10492 27261 10520
rect 27120 10480 27126 10492
rect 27249 10489 27261 10492
rect 27295 10520 27307 10523
rect 27754 10523 27812 10529
rect 27754 10520 27766 10523
rect 27295 10492 27766 10520
rect 27295 10489 27307 10492
rect 27249 10483 27307 10489
rect 27754 10489 27766 10492
rect 27800 10520 27812 10523
rect 28534 10520 28540 10532
rect 27800 10492 28540 10520
rect 27800 10489 27812 10492
rect 27754 10483 27812 10489
rect 28534 10480 28540 10492
rect 28592 10480 28598 10532
rect 20441 10455 20499 10461
rect 20441 10452 20453 10455
rect 19484 10424 20453 10452
rect 19484 10412 19490 10424
rect 20441 10421 20453 10424
rect 20487 10421 20499 10455
rect 22646 10452 22652 10464
rect 22607 10424 22652 10452
rect 20441 10415 20499 10421
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 24578 10412 24584 10464
rect 24636 10452 24642 10464
rect 25777 10455 25835 10461
rect 25777 10452 25789 10455
rect 24636 10424 25789 10452
rect 24636 10412 24642 10424
rect 25777 10421 25789 10424
rect 25823 10421 25835 10455
rect 28350 10452 28356 10464
rect 28311 10424 28356 10452
rect 25777 10415 25835 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 28626 10452 28632 10464
rect 28587 10424 28632 10452
rect 28626 10412 28632 10424
rect 28684 10412 28690 10464
rect 29932 10461 29960 10560
rect 30374 10548 30380 10560
rect 30432 10548 30438 10600
rect 30466 10548 30472 10600
rect 30524 10588 30530 10600
rect 31665 10591 31723 10597
rect 31665 10588 31677 10591
rect 30524 10560 31677 10588
rect 30524 10548 30530 10560
rect 31665 10557 31677 10560
rect 31711 10588 31723 10591
rect 33410 10588 33416 10600
rect 31711 10560 33416 10588
rect 31711 10557 31723 10560
rect 31665 10551 31723 10557
rect 33410 10548 33416 10560
rect 33468 10548 33474 10600
rect 33502 10548 33508 10600
rect 33560 10588 33566 10600
rect 34885 10591 34943 10597
rect 34885 10588 34897 10591
rect 33560 10560 34897 10588
rect 33560 10548 33566 10560
rect 34885 10557 34897 10560
rect 34931 10588 34943 10591
rect 35345 10591 35403 10597
rect 35345 10588 35357 10591
rect 34931 10560 35357 10588
rect 34931 10557 34943 10560
rect 34885 10551 34943 10557
rect 35345 10557 35357 10560
rect 35391 10557 35403 10591
rect 35345 10551 35403 10557
rect 38746 10548 38752 10600
rect 38804 10588 38810 10600
rect 39117 10591 39175 10597
rect 39117 10588 39129 10591
rect 38804 10560 39129 10588
rect 38804 10548 38810 10560
rect 39117 10557 39129 10560
rect 39163 10588 39175 10591
rect 42242 10588 42248 10600
rect 39163 10560 42248 10588
rect 39163 10557 39175 10560
rect 39117 10551 39175 10557
rect 42242 10548 42248 10560
rect 42300 10548 42306 10600
rect 42444 10588 42472 10755
rect 43714 10752 43720 10764
rect 43772 10752 43778 10804
rect 43898 10752 43904 10804
rect 43956 10792 43962 10804
rect 44913 10795 44971 10801
rect 44913 10792 44925 10795
rect 43956 10764 44925 10792
rect 43956 10752 43962 10764
rect 44913 10761 44925 10764
rect 44959 10761 44971 10795
rect 44913 10755 44971 10761
rect 45186 10752 45192 10804
rect 45244 10792 45250 10804
rect 45465 10795 45523 10801
rect 45465 10792 45477 10795
rect 45244 10764 45477 10792
rect 45244 10752 45250 10764
rect 45465 10761 45477 10764
rect 45511 10792 45523 10795
rect 47486 10792 47492 10804
rect 45511 10764 47492 10792
rect 45511 10761 45523 10764
rect 45465 10755 45523 10761
rect 47486 10752 47492 10764
rect 47544 10752 47550 10804
rect 43732 10656 43760 10752
rect 43809 10727 43867 10733
rect 43809 10693 43821 10727
rect 43855 10724 43867 10727
rect 43990 10724 43996 10736
rect 43855 10696 43996 10724
rect 43855 10693 43867 10696
rect 43809 10687 43867 10693
rect 43990 10684 43996 10696
rect 44048 10684 44054 10736
rect 44542 10724 44548 10736
rect 44503 10696 44548 10724
rect 44542 10684 44548 10696
rect 44600 10684 44606 10736
rect 44082 10656 44088 10668
rect 43732 10628 44088 10656
rect 44082 10616 44088 10628
rect 44140 10616 44146 10668
rect 42648 10591 42706 10597
rect 42648 10588 42660 10591
rect 42444 10560 42660 10588
rect 42648 10557 42660 10560
rect 42694 10557 42706 10591
rect 42648 10551 42706 10557
rect 45925 10591 45983 10597
rect 45925 10557 45937 10591
rect 45971 10588 45983 10591
rect 46750 10588 46756 10600
rect 45971 10560 46756 10588
rect 45971 10557 45983 10560
rect 45925 10551 45983 10557
rect 46750 10548 46756 10560
rect 46808 10548 46814 10600
rect 30285 10523 30343 10529
rect 30285 10489 30297 10523
rect 30331 10520 30343 10523
rect 30698 10523 30756 10529
rect 30698 10520 30710 10523
rect 30331 10492 30710 10520
rect 30331 10489 30343 10492
rect 30285 10483 30343 10489
rect 30698 10489 30710 10492
rect 30744 10520 30756 10523
rect 31941 10523 31999 10529
rect 31941 10520 31953 10523
rect 30744 10492 31953 10520
rect 30744 10489 30756 10492
rect 30698 10483 30756 10489
rect 31941 10489 31953 10492
rect 31987 10520 31999 10523
rect 32446 10523 32504 10529
rect 32446 10520 32458 10523
rect 31987 10492 32458 10520
rect 31987 10489 31999 10492
rect 31941 10483 31999 10489
rect 32446 10489 32458 10492
rect 32492 10520 32504 10523
rect 35710 10520 35716 10532
rect 32492 10492 35716 10520
rect 32492 10489 32504 10492
rect 32446 10483 32504 10489
rect 35710 10480 35716 10492
rect 35768 10520 35774 10532
rect 35897 10523 35955 10529
rect 35897 10520 35909 10523
rect 35768 10492 35909 10520
rect 35768 10480 35774 10492
rect 35897 10489 35909 10492
rect 35943 10520 35955 10523
rect 36402 10523 36460 10529
rect 36402 10520 36414 10523
rect 35943 10492 36414 10520
rect 35943 10489 35955 10492
rect 35897 10483 35955 10489
rect 36402 10489 36414 10492
rect 36448 10520 36460 10523
rect 37645 10523 37703 10529
rect 37645 10520 37657 10523
rect 36448 10492 37657 10520
rect 36448 10489 36460 10492
rect 36402 10483 36460 10489
rect 37645 10489 37657 10492
rect 37691 10520 37703 10523
rect 38010 10520 38016 10532
rect 37691 10492 38016 10520
rect 37691 10489 37703 10492
rect 37645 10483 37703 10489
rect 38010 10480 38016 10492
rect 38068 10520 38074 10532
rect 38150 10523 38208 10529
rect 38150 10520 38162 10523
rect 38068 10492 38162 10520
rect 38068 10480 38074 10492
rect 38150 10489 38162 10492
rect 38196 10489 38208 10523
rect 38150 10483 38208 10489
rect 40862 10480 40868 10532
rect 40920 10520 40926 10532
rect 41186 10523 41244 10529
rect 41186 10520 41198 10523
rect 40920 10492 41198 10520
rect 40920 10480 40926 10492
rect 41186 10489 41198 10492
rect 41232 10489 41244 10523
rect 41186 10483 41244 10489
rect 43806 10480 43812 10532
rect 43864 10520 43870 10532
rect 43993 10523 44051 10529
rect 43993 10520 44005 10523
rect 43864 10492 44005 10520
rect 43864 10480 43870 10492
rect 43993 10489 44005 10492
rect 44039 10489 44051 10523
rect 43993 10483 44051 10489
rect 44082 10480 44088 10532
rect 44140 10520 44146 10532
rect 46106 10520 46112 10532
rect 44140 10492 44185 10520
rect 46067 10492 46112 10520
rect 44140 10480 44146 10492
rect 46106 10480 46112 10492
rect 46164 10480 46170 10532
rect 29917 10455 29975 10461
rect 29917 10421 29929 10455
rect 29963 10452 29975 10455
rect 30098 10452 30104 10464
rect 29963 10424 30104 10452
rect 29963 10421 29975 10424
rect 29917 10415 29975 10421
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 32122 10412 32128 10464
rect 32180 10452 32186 10464
rect 33045 10455 33103 10461
rect 33045 10452 33057 10455
rect 32180 10424 33057 10452
rect 32180 10412 32186 10424
rect 33045 10421 33057 10424
rect 33091 10421 33103 10455
rect 33045 10415 33103 10421
rect 34333 10455 34391 10461
rect 34333 10421 34345 10455
rect 34379 10452 34391 10455
rect 35526 10452 35532 10464
rect 34379 10424 35532 10452
rect 34379 10421 34391 10424
rect 34333 10415 34391 10421
rect 35526 10412 35532 10424
rect 35584 10412 35590 10464
rect 36998 10452 37004 10464
rect 36959 10424 37004 10452
rect 36998 10412 37004 10424
rect 37056 10412 37062 10464
rect 38746 10452 38752 10464
rect 38707 10424 38752 10452
rect 38746 10412 38752 10424
rect 38804 10412 38810 10464
rect 39482 10452 39488 10464
rect 39443 10424 39488 10452
rect 39482 10412 39488 10424
rect 39540 10412 39546 10464
rect 39942 10452 39948 10464
rect 39903 10424 39948 10452
rect 39942 10412 39948 10424
rect 40000 10412 40006 10464
rect 42518 10412 42524 10464
rect 42576 10452 42582 10464
rect 42751 10455 42809 10461
rect 42751 10452 42763 10455
rect 42576 10424 42763 10452
rect 42576 10412 42582 10424
rect 42751 10421 42763 10424
rect 42797 10421 42809 10455
rect 42751 10415 42809 10421
rect 1104 10362 48852 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 48852 10362
rect 1104 10288 48852 10310
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 17552 10220 19809 10248
rect 17552 10208 17558 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 20036 10220 20085 10248
rect 20036 10208 20042 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 21634 10248 21640 10260
rect 21595 10220 21640 10248
rect 20073 10211 20131 10217
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 22557 10251 22615 10257
rect 22557 10248 22569 10251
rect 21784 10220 22569 10248
rect 21784 10208 21790 10220
rect 22557 10217 22569 10220
rect 22603 10217 22615 10251
rect 22557 10211 22615 10217
rect 23247 10251 23305 10257
rect 23247 10217 23259 10251
rect 23293 10248 23305 10251
rect 23842 10248 23848 10260
rect 23293 10220 23848 10248
rect 23293 10217 23305 10220
rect 23247 10211 23305 10217
rect 23842 10208 23848 10220
rect 23900 10208 23906 10260
rect 24397 10251 24455 10257
rect 24397 10217 24409 10251
rect 24443 10248 24455 10251
rect 24578 10248 24584 10260
rect 24443 10220 24584 10248
rect 24443 10217 24455 10220
rect 24397 10211 24455 10217
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 24762 10208 24768 10260
rect 24820 10248 24826 10260
rect 25133 10251 25191 10257
rect 25133 10248 25145 10251
rect 24820 10220 25145 10248
rect 24820 10208 24826 10220
rect 25133 10217 25145 10220
rect 25179 10217 25191 10251
rect 25133 10211 25191 10217
rect 26651 10251 26709 10257
rect 26651 10217 26663 10251
rect 26697 10248 26709 10251
rect 26786 10248 26792 10260
rect 26697 10220 26792 10248
rect 26697 10217 26709 10220
rect 26651 10211 26709 10217
rect 26786 10208 26792 10220
rect 26844 10208 26850 10260
rect 28442 10248 28448 10260
rect 28403 10220 28448 10248
rect 28442 10208 28448 10220
rect 28500 10208 28506 10260
rect 30006 10248 30012 10260
rect 29967 10220 30012 10248
rect 30006 10208 30012 10220
rect 30064 10208 30070 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 30469 10251 30527 10257
rect 30469 10248 30481 10251
rect 30432 10220 30481 10248
rect 30432 10208 30438 10220
rect 30469 10217 30481 10220
rect 30515 10248 30527 10251
rect 31205 10251 31263 10257
rect 31205 10248 31217 10251
rect 30515 10220 31217 10248
rect 30515 10217 30527 10220
rect 30469 10211 30527 10217
rect 31205 10217 31217 10220
rect 31251 10217 31263 10251
rect 32306 10248 32312 10260
rect 32267 10220 32312 10248
rect 31205 10211 31263 10217
rect 32306 10208 32312 10220
rect 32364 10208 32370 10260
rect 36078 10248 36084 10260
rect 36039 10220 36084 10248
rect 36078 10208 36084 10220
rect 36136 10208 36142 10260
rect 37826 10208 37832 10260
rect 37884 10248 37890 10260
rect 37921 10251 37979 10257
rect 37921 10248 37933 10251
rect 37884 10220 37933 10248
rect 37884 10208 37890 10220
rect 37921 10217 37933 10220
rect 37967 10217 37979 10251
rect 37921 10211 37979 10217
rect 39942 10208 39948 10260
rect 40000 10248 40006 10260
rect 40221 10251 40279 10257
rect 40221 10248 40233 10251
rect 40000 10220 40233 10248
rect 40000 10208 40006 10220
rect 40221 10217 40233 10220
rect 40267 10217 40279 10251
rect 41138 10248 41144 10260
rect 41099 10220 41144 10248
rect 40221 10211 40279 10217
rect 41138 10208 41144 10220
rect 41196 10208 41202 10260
rect 43717 10251 43775 10257
rect 43717 10217 43729 10251
rect 43763 10248 43775 10251
rect 43806 10248 43812 10260
rect 43763 10220 43812 10248
rect 43763 10217 43775 10220
rect 43717 10211 43775 10217
rect 43806 10208 43812 10220
rect 43864 10208 43870 10260
rect 46750 10208 46756 10260
rect 46808 10248 46814 10260
rect 47673 10251 47731 10257
rect 47673 10248 47685 10251
rect 46808 10220 47685 10248
rect 46808 10208 46814 10220
rect 47673 10217 47685 10220
rect 47719 10217 47731 10251
rect 47673 10211 47731 10217
rect 18230 10140 18236 10192
rect 18288 10140 18294 10192
rect 24854 10180 24860 10192
rect 24136 10152 24860 10180
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 16172 10084 17509 10112
rect 16172 10072 16178 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 17497 10075 17555 10081
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 19337 10115 19395 10121
rect 19337 10112 19349 10115
rect 19208 10084 19349 10112
rect 19208 10072 19214 10084
rect 19337 10081 19349 10084
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 21508 10084 21557 10112
rect 21508 10072 21514 10084
rect 21545 10081 21557 10084
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 22097 10115 22155 10121
rect 22097 10081 22109 10115
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 22112 10044 22140 10075
rect 22646 10072 22652 10124
rect 22704 10112 22710 10124
rect 24136 10121 24164 10152
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 27062 10140 27068 10192
rect 27120 10180 27126 10192
rect 27846 10183 27904 10189
rect 27846 10180 27858 10183
rect 27120 10152 27858 10180
rect 27120 10140 27126 10152
rect 27846 10149 27858 10152
rect 27892 10149 27904 10183
rect 27846 10143 27904 10149
rect 32861 10183 32919 10189
rect 32861 10149 32873 10183
rect 32907 10180 32919 10183
rect 33686 10180 33692 10192
rect 32907 10152 33692 10180
rect 32907 10149 32919 10152
rect 32861 10143 32919 10149
rect 33686 10140 33692 10152
rect 33744 10140 33750 10192
rect 38749 10183 38807 10189
rect 38749 10149 38761 10183
rect 38795 10180 38807 10183
rect 39022 10180 39028 10192
rect 38795 10152 39028 10180
rect 38795 10149 38807 10152
rect 38749 10143 38807 10149
rect 39022 10140 39028 10152
rect 39080 10140 39086 10192
rect 41782 10180 41788 10192
rect 41743 10152 41788 10180
rect 41782 10140 41788 10152
rect 41840 10140 41846 10192
rect 41877 10183 41935 10189
rect 41877 10149 41889 10183
rect 41923 10180 41935 10183
rect 42242 10180 42248 10192
rect 41923 10152 42248 10180
rect 41923 10149 41935 10152
rect 41877 10143 41935 10149
rect 42242 10140 42248 10152
rect 42300 10140 42306 10192
rect 42429 10183 42487 10189
rect 42429 10149 42441 10183
rect 42475 10180 42487 10183
rect 43070 10180 43076 10192
rect 42475 10152 43076 10180
rect 42475 10149 42487 10152
rect 42429 10143 42487 10149
rect 43070 10140 43076 10152
rect 43128 10180 43134 10192
rect 43898 10180 43904 10192
rect 43128 10152 43904 10180
rect 43128 10140 43134 10152
rect 43898 10140 43904 10152
rect 43956 10140 43962 10192
rect 43993 10183 44051 10189
rect 43993 10149 44005 10183
rect 44039 10180 44051 10183
rect 44082 10180 44088 10192
rect 44039 10152 44088 10180
rect 44039 10149 44051 10152
rect 43993 10143 44051 10149
rect 44082 10140 44088 10152
rect 44140 10140 44146 10192
rect 23144 10115 23202 10121
rect 23144 10112 23156 10115
rect 22704 10084 23156 10112
rect 22704 10072 22710 10084
rect 23144 10081 23156 10084
rect 23190 10081 23202 10115
rect 23144 10075 23202 10081
rect 24121 10115 24179 10121
rect 24121 10081 24133 10115
rect 24167 10081 24179 10115
rect 24121 10075 24179 10081
rect 24210 10072 24216 10124
rect 24268 10112 24274 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 24268 10084 24593 10112
rect 24268 10072 24274 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 25498 10072 25504 10124
rect 25556 10112 25562 10124
rect 26234 10112 26240 10124
rect 25556 10084 26240 10112
rect 25556 10072 25562 10084
rect 26234 10072 26240 10084
rect 26292 10112 26298 10124
rect 26548 10115 26606 10121
rect 26548 10112 26560 10115
rect 26292 10084 26560 10112
rect 26292 10072 26298 10084
rect 26548 10081 26560 10084
rect 26594 10081 26606 10115
rect 26548 10075 26606 10081
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10112 27583 10115
rect 28166 10112 28172 10124
rect 27571 10084 28172 10112
rect 27571 10081 27583 10084
rect 27525 10075 27583 10081
rect 28166 10072 28172 10084
rect 28224 10112 28230 10124
rect 28718 10112 28724 10124
rect 28224 10084 28724 10112
rect 28224 10072 28230 10084
rect 28718 10072 28724 10084
rect 28776 10072 28782 10124
rect 30374 10112 30380 10124
rect 30335 10084 30380 10112
rect 30374 10072 30380 10084
rect 30432 10072 30438 10124
rect 30745 10115 30803 10121
rect 30745 10081 30757 10115
rect 30791 10081 30803 10115
rect 33042 10112 33048 10124
rect 33003 10084 33048 10112
rect 30745 10075 30803 10081
rect 24228 10044 24256 10072
rect 22060 10016 24256 10044
rect 22060 10004 22066 10016
rect 30006 10004 30012 10056
rect 30064 10044 30070 10056
rect 30650 10044 30656 10056
rect 30064 10016 30656 10044
rect 30064 10004 30070 10016
rect 30650 10004 30656 10016
rect 30708 10044 30714 10056
rect 30760 10044 30788 10075
rect 33042 10072 33048 10084
rect 33100 10072 33106 10124
rect 35161 10115 35219 10121
rect 35161 10081 35173 10115
rect 35207 10081 35219 10115
rect 35161 10075 35219 10081
rect 35437 10115 35495 10121
rect 35437 10081 35449 10115
rect 35483 10112 35495 10115
rect 35526 10112 35532 10124
rect 35483 10084 35532 10112
rect 35483 10081 35495 10084
rect 35437 10075 35495 10081
rect 30708 10016 30788 10044
rect 30708 10004 30714 10016
rect 35176 9976 35204 10075
rect 35526 10072 35532 10084
rect 35584 10072 35590 10124
rect 36446 10112 36452 10124
rect 36407 10084 36452 10112
rect 36446 10072 36452 10084
rect 36504 10072 36510 10124
rect 39666 10072 39672 10124
rect 39724 10112 39730 10124
rect 40126 10112 40132 10124
rect 39724 10084 40132 10112
rect 39724 10072 39730 10084
rect 40126 10072 40132 10084
rect 40184 10072 40190 10124
rect 40681 10115 40739 10121
rect 40681 10081 40693 10115
rect 40727 10112 40739 10115
rect 40954 10112 40960 10124
rect 40727 10084 40960 10112
rect 40727 10081 40739 10084
rect 40681 10075 40739 10081
rect 40954 10072 40960 10084
rect 41012 10072 41018 10124
rect 46014 10112 46020 10124
rect 45975 10084 46020 10112
rect 46014 10072 46020 10084
rect 46072 10072 46078 10124
rect 47486 10112 47492 10124
rect 47447 10084 47492 10112
rect 47486 10072 47492 10084
rect 47544 10072 47550 10124
rect 35618 10044 35624 10056
rect 35579 10016 35624 10044
rect 35618 10004 35624 10016
rect 35676 10004 35682 10056
rect 38654 10044 38660 10056
rect 38615 10016 38660 10044
rect 38654 10004 38660 10016
rect 38712 10004 38718 10056
rect 43898 10044 43904 10056
rect 43859 10016 43904 10044
rect 43898 10004 43904 10016
rect 43956 10004 43962 10056
rect 45922 10044 45928 10056
rect 45883 10016 45928 10044
rect 45922 10004 45928 10016
rect 45980 10004 45986 10056
rect 35250 9976 35256 9988
rect 35163 9948 35256 9976
rect 35250 9936 35256 9948
rect 35308 9976 35314 9988
rect 35802 9976 35808 9988
rect 35308 9948 35808 9976
rect 35308 9936 35314 9948
rect 35802 9936 35808 9948
rect 35860 9936 35866 9988
rect 39209 9979 39267 9985
rect 39209 9945 39221 9979
rect 39255 9945 39267 9979
rect 44450 9976 44456 9988
rect 44411 9948 44456 9976
rect 39209 9939 39267 9945
rect 23842 9908 23848 9920
rect 23803 9880 23848 9908
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 27157 9911 27215 9917
rect 27157 9877 27169 9911
rect 27203 9908 27215 9911
rect 27430 9908 27436 9920
rect 27203 9880 27436 9908
rect 27203 9877 27215 9880
rect 27157 9871 27215 9877
rect 27430 9868 27436 9880
rect 27488 9868 27494 9920
rect 29270 9908 29276 9920
rect 29231 9880 29276 9908
rect 29270 9868 29276 9880
rect 29328 9868 29334 9920
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 33137 9911 33195 9917
rect 33137 9908 33149 9911
rect 30156 9880 33149 9908
rect 30156 9868 30162 9880
rect 33137 9877 33149 9880
rect 33183 9877 33195 9911
rect 33137 9871 33195 9877
rect 35894 9868 35900 9920
rect 35952 9908 35958 9920
rect 36633 9911 36691 9917
rect 36633 9908 36645 9911
rect 35952 9880 36645 9908
rect 35952 9868 35958 9880
rect 36633 9877 36645 9880
rect 36679 9877 36691 9911
rect 39224 9908 39252 9939
rect 44450 9936 44456 9948
rect 44508 9936 44514 9988
rect 39298 9908 39304 9920
rect 39211 9880 39304 9908
rect 36633 9871 36691 9877
rect 39298 9868 39304 9880
rect 39356 9908 39362 9920
rect 43806 9908 43812 9920
rect 39356 9880 43812 9908
rect 39356 9868 39362 9880
rect 43806 9868 43812 9880
rect 43864 9868 43870 9920
rect 1104 9818 48852 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 48852 9818
rect 1104 9744 48852 9766
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 16172 9676 16773 9704
rect 16172 9664 16178 9676
rect 16761 9673 16773 9676
rect 16807 9673 16819 9707
rect 16761 9667 16819 9673
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 19383 9707 19441 9713
rect 19383 9704 19395 9707
rect 17920 9676 19395 9704
rect 17920 9664 17926 9676
rect 19383 9673 19395 9676
rect 19429 9673 19441 9707
rect 22002 9704 22008 9716
rect 21963 9676 22008 9704
rect 19383 9667 19441 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22465 9707 22523 9713
rect 22465 9673 22477 9707
rect 22511 9704 22523 9707
rect 22646 9704 22652 9716
rect 22511 9676 22652 9704
rect 22511 9673 22523 9676
rect 22465 9667 22523 9673
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 25682 9704 25688 9716
rect 25643 9676 25688 9704
rect 25682 9664 25688 9676
rect 25740 9664 25746 9716
rect 29089 9707 29147 9713
rect 29089 9673 29101 9707
rect 29135 9704 29147 9707
rect 29178 9704 29184 9716
rect 29135 9676 29184 9704
rect 29135 9673 29147 9676
rect 29089 9667 29147 9673
rect 29178 9664 29184 9676
rect 29236 9664 29242 9716
rect 30374 9704 30380 9716
rect 30335 9676 30380 9704
rect 30374 9664 30380 9676
rect 30432 9664 30438 9716
rect 30650 9704 30656 9716
rect 30611 9676 30656 9704
rect 30650 9664 30656 9676
rect 30708 9664 30714 9716
rect 32398 9704 32404 9716
rect 32359 9676 32404 9704
rect 32398 9664 32404 9676
rect 32456 9664 32462 9716
rect 32674 9704 32680 9716
rect 32635 9676 32680 9704
rect 32674 9664 32680 9676
rect 32732 9664 32738 9716
rect 33042 9664 33048 9716
rect 33100 9704 33106 9716
rect 33321 9707 33379 9713
rect 33321 9704 33333 9707
rect 33100 9676 33333 9704
rect 33100 9664 33106 9676
rect 33321 9673 33333 9676
rect 33367 9673 33379 9707
rect 33686 9704 33692 9716
rect 33647 9676 33692 9704
rect 33321 9667 33379 9673
rect 33686 9664 33692 9676
rect 33744 9664 33750 9716
rect 34701 9707 34759 9713
rect 34701 9673 34713 9707
rect 34747 9704 34759 9707
rect 35526 9704 35532 9716
rect 34747 9676 35532 9704
rect 34747 9673 34759 9676
rect 34701 9667 34759 9673
rect 35526 9664 35532 9676
rect 35584 9664 35590 9716
rect 36446 9664 36452 9716
rect 36504 9704 36510 9716
rect 37001 9707 37059 9713
rect 37001 9704 37013 9707
rect 36504 9676 37013 9704
rect 36504 9664 36510 9676
rect 37001 9673 37013 9676
rect 37047 9673 37059 9707
rect 37001 9667 37059 9673
rect 38473 9707 38531 9713
rect 38473 9673 38485 9707
rect 38519 9704 38531 9707
rect 38654 9704 38660 9716
rect 38519 9676 38660 9704
rect 38519 9673 38531 9676
rect 38473 9667 38531 9673
rect 38654 9664 38660 9676
rect 38712 9713 38718 9716
rect 38712 9707 38761 9713
rect 38712 9673 38715 9707
rect 38749 9673 38761 9707
rect 39022 9704 39028 9716
rect 38983 9676 39028 9704
rect 38712 9667 38761 9673
rect 38712 9664 38718 9667
rect 39022 9664 39028 9676
rect 39080 9664 39086 9716
rect 39482 9664 39488 9716
rect 39540 9704 39546 9716
rect 40635 9707 40693 9713
rect 40635 9704 40647 9707
rect 39540 9676 40647 9704
rect 39540 9664 39546 9676
rect 40635 9673 40647 9676
rect 40681 9673 40693 9707
rect 40954 9704 40960 9716
rect 40915 9676 40960 9704
rect 40635 9667 40693 9673
rect 40954 9664 40960 9676
rect 41012 9664 41018 9716
rect 41785 9707 41843 9713
rect 41785 9673 41797 9707
rect 41831 9704 41843 9707
rect 41874 9704 41880 9716
rect 41831 9676 41880 9704
rect 41831 9673 41843 9676
rect 41785 9667 41843 9673
rect 41874 9664 41880 9676
rect 41932 9704 41938 9716
rect 42242 9704 42248 9716
rect 41932 9676 42248 9704
rect 41932 9664 41938 9676
rect 42242 9664 42248 9676
rect 42300 9664 42306 9716
rect 43533 9707 43591 9713
rect 43533 9673 43545 9707
rect 43579 9704 43591 9707
rect 44082 9704 44088 9716
rect 43579 9676 44088 9704
rect 43579 9673 43591 9676
rect 43533 9667 43591 9673
rect 44082 9664 44088 9676
rect 44140 9664 44146 9716
rect 45922 9704 45928 9716
rect 45883 9676 45928 9704
rect 45922 9664 45928 9676
rect 45980 9664 45986 9716
rect 47486 9704 47492 9716
rect 47447 9676 47492 9704
rect 47486 9664 47492 9676
rect 47544 9664 47550 9716
rect 19150 9568 19156 9580
rect 17512 9540 19156 9568
rect 16206 9500 16212 9512
rect 13786 9472 16212 9500
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 13786 9432 13814 9472
rect 16206 9460 16212 9472
rect 16264 9500 16270 9512
rect 17512 9509 17540 9540
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19484 9540 20269 9568
rect 19484 9528 19490 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 25700 9568 25728 9664
rect 31021 9639 31079 9645
rect 31021 9636 31033 9639
rect 29748 9608 31033 9636
rect 25700 9540 25820 9568
rect 20257 9531 20315 9537
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 16264 9472 17509 9500
rect 16264 9460 16270 9472
rect 17497 9469 17509 9472
rect 17543 9469 17555 9503
rect 17497 9463 17555 9469
rect 18300 9503 18358 9509
rect 18300 9469 18312 9503
rect 18346 9500 18358 9503
rect 19312 9503 19370 9509
rect 18346 9472 18828 9500
rect 18346 9469 18358 9472
rect 18300 9463 18358 9469
rect 18138 9432 18144 9444
rect 11020 9404 13814 9432
rect 17144 9404 18144 9432
rect 11020 9392 11026 9404
rect 17144 9376 17172 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18800 9376 18828 9472
rect 19312 9469 19324 9503
rect 19358 9500 19370 9503
rect 20162 9500 20168 9512
rect 19358 9472 19840 9500
rect 20075 9472 20168 9500
rect 19358 9469 19370 9472
rect 19312 9463 19370 9469
rect 17126 9364 17132 9376
rect 17087 9336 17132 9364
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 18371 9367 18429 9373
rect 18371 9333 18383 9367
rect 18417 9364 18429 9367
rect 18598 9364 18604 9376
rect 18417 9336 18604 9364
rect 18417 9333 18429 9336
rect 18371 9327 18429 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 18782 9364 18788 9376
rect 18743 9336 18788 9364
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19812 9373 19840 9472
rect 20162 9460 20168 9472
rect 20220 9500 20226 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 20220 9472 20361 9500
rect 20220 9460 20226 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 22624 9503 22682 9509
rect 22624 9469 22636 9503
rect 22670 9500 22682 9503
rect 22670 9472 23152 9500
rect 22670 9469 22682 9472
rect 22624 9463 22682 9469
rect 23124 9376 23152 9472
rect 23474 9460 23480 9512
rect 23532 9500 23538 9512
rect 23750 9500 23756 9512
rect 23532 9472 23756 9500
rect 23532 9460 23538 9472
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 23842 9460 23848 9512
rect 23900 9500 23906 9512
rect 24118 9500 24124 9512
rect 23900 9472 24124 9500
rect 23900 9460 23906 9472
rect 24118 9460 24124 9472
rect 24176 9500 24182 9512
rect 24213 9503 24271 9509
rect 24213 9500 24225 9503
rect 24176 9472 24225 9500
rect 24176 9460 24182 9472
rect 24213 9469 24225 9472
rect 24259 9500 24271 9503
rect 25682 9500 25688 9512
rect 24259 9472 25688 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 25792 9509 25820 9540
rect 25777 9503 25835 9509
rect 25777 9469 25789 9503
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 26237 9503 26295 9509
rect 26237 9469 26249 9503
rect 26283 9469 26295 9503
rect 26237 9463 26295 9469
rect 27893 9503 27951 9509
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 27893 9463 27951 9469
rect 25700 9432 25728 9460
rect 26252 9432 26280 9463
rect 26510 9432 26516 9444
rect 25700 9404 26280 9432
rect 26471 9404 26516 9432
rect 26510 9392 26516 9404
rect 26568 9392 26574 9444
rect 27157 9435 27215 9441
rect 27157 9401 27169 9435
rect 27203 9432 27215 9435
rect 27908 9432 27936 9463
rect 27982 9460 27988 9512
rect 28040 9500 28046 9512
rect 28169 9503 28227 9509
rect 28169 9500 28181 9503
rect 28040 9472 28181 9500
rect 28040 9460 28046 9472
rect 28169 9469 28181 9472
rect 28215 9500 28227 9503
rect 28994 9500 29000 9512
rect 28215 9472 29000 9500
rect 28215 9469 28227 9472
rect 28169 9463 28227 9469
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 29178 9460 29184 9512
rect 29236 9500 29242 9512
rect 29273 9503 29331 9509
rect 29273 9500 29285 9503
rect 29236 9472 29285 9500
rect 29236 9460 29242 9472
rect 29273 9469 29285 9472
rect 29319 9469 29331 9503
rect 29273 9463 29331 9469
rect 29362 9460 29368 9512
rect 29420 9500 29426 9512
rect 29748 9509 29776 9608
rect 31021 9605 31033 9608
rect 31067 9605 31079 9639
rect 31021 9599 31079 9605
rect 35161 9639 35219 9645
rect 35161 9605 35173 9639
rect 35207 9636 35219 9639
rect 35250 9636 35256 9648
rect 35207 9608 35256 9636
rect 35207 9605 35219 9608
rect 35161 9599 35219 9605
rect 35250 9596 35256 9608
rect 35308 9596 35314 9648
rect 35710 9636 35716 9648
rect 35671 9608 35716 9636
rect 35710 9596 35716 9608
rect 35768 9596 35774 9648
rect 40126 9636 40132 9648
rect 40087 9608 40132 9636
rect 40126 9596 40132 9608
rect 40184 9596 40190 9648
rect 43070 9636 43076 9648
rect 43031 9608 43076 9636
rect 43070 9596 43076 9608
rect 43128 9596 43134 9648
rect 45557 9639 45615 9645
rect 45557 9605 45569 9639
rect 45603 9636 45615 9639
rect 46014 9636 46020 9648
rect 45603 9608 46020 9636
rect 45603 9605 45615 9608
rect 45557 9599 45615 9605
rect 46014 9596 46020 9608
rect 46072 9596 46078 9648
rect 35618 9528 35624 9580
rect 35676 9568 35682 9580
rect 35805 9571 35863 9577
rect 35805 9568 35817 9571
rect 35676 9540 35817 9568
rect 35676 9528 35682 9540
rect 35805 9537 35817 9540
rect 35851 9537 35863 9571
rect 35805 9531 35863 9537
rect 36998 9528 37004 9580
rect 37056 9568 37062 9580
rect 39393 9571 39451 9577
rect 39393 9568 39405 9571
rect 37056 9540 39405 9568
rect 37056 9528 37062 9540
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29420 9472 29745 9500
rect 29420 9460 29426 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 30190 9460 30196 9512
rect 30248 9500 30254 9512
rect 30837 9503 30895 9509
rect 30837 9500 30849 9503
rect 30248 9472 30849 9500
rect 30248 9460 30254 9472
rect 30837 9469 30849 9472
rect 30883 9500 30895 9503
rect 31297 9503 31355 9509
rect 31297 9500 31309 9503
rect 30883 9472 31309 9500
rect 30883 9469 30895 9472
rect 30837 9463 30895 9469
rect 31297 9469 31309 9472
rect 31343 9469 31355 9503
rect 31297 9463 31355 9469
rect 31849 9503 31907 9509
rect 31849 9469 31861 9503
rect 31895 9500 31907 9503
rect 32398 9500 32404 9512
rect 31895 9472 32404 9500
rect 31895 9469 31907 9472
rect 31849 9463 31907 9469
rect 32398 9460 32404 9472
rect 32456 9460 32462 9512
rect 32674 9460 32680 9512
rect 32732 9500 32738 9512
rect 32861 9503 32919 9509
rect 32861 9500 32873 9503
rect 32732 9472 32873 9500
rect 32732 9460 32738 9472
rect 32861 9469 32873 9472
rect 32907 9469 32919 9503
rect 32861 9463 32919 9469
rect 34422 9460 34428 9512
rect 34480 9500 34486 9512
rect 38615 9509 38643 9540
rect 39393 9537 39405 9540
rect 39439 9537 39451 9571
rect 42518 9568 42524 9580
rect 42479 9540 42524 9568
rect 39393 9531 39451 9537
rect 42518 9528 42524 9540
rect 42576 9528 42582 9580
rect 43254 9528 43260 9580
rect 43312 9568 43318 9580
rect 43898 9568 43904 9580
rect 43312 9540 43904 9568
rect 43312 9528 43318 9540
rect 43898 9528 43904 9540
rect 43956 9568 43962 9580
rect 44361 9571 44419 9577
rect 44361 9568 44373 9571
rect 43956 9540 44373 9568
rect 43956 9528 43962 9540
rect 44361 9537 44373 9540
rect 44407 9568 44419 9571
rect 45005 9571 45063 9577
rect 45005 9568 45017 9571
rect 44407 9540 45017 9568
rect 44407 9537 44419 9540
rect 44361 9531 44419 9537
rect 45005 9537 45017 9540
rect 45051 9537 45063 9571
rect 45005 9531 45063 9537
rect 46201 9571 46259 9577
rect 46201 9537 46213 9571
rect 46247 9568 46259 9571
rect 46382 9568 46388 9580
rect 46247 9540 46388 9568
rect 46247 9537 46259 9540
rect 46201 9531 46259 9537
rect 46382 9528 46388 9540
rect 46440 9568 46446 9580
rect 47121 9571 47179 9577
rect 47121 9568 47133 9571
rect 46440 9540 47133 9568
rect 46440 9528 46446 9540
rect 47121 9537 47133 9540
rect 47167 9537 47179 9571
rect 47121 9531 47179 9537
rect 37553 9503 37611 9509
rect 37553 9500 37565 9503
rect 34480 9472 37565 9500
rect 34480 9460 34486 9472
rect 37553 9469 37565 9472
rect 37599 9500 37611 9503
rect 38013 9503 38071 9509
rect 38013 9500 38025 9503
rect 37599 9472 38025 9500
rect 37599 9469 37611 9472
rect 37553 9463 37611 9469
rect 38013 9469 38025 9472
rect 38059 9469 38071 9503
rect 38013 9463 38071 9469
rect 38600 9503 38658 9509
rect 38600 9469 38612 9503
rect 38646 9469 38658 9503
rect 38600 9463 38658 9469
rect 38746 9460 38752 9512
rect 38804 9500 38810 9512
rect 40532 9503 40590 9509
rect 40532 9500 40544 9503
rect 38804 9472 40544 9500
rect 38804 9460 38810 9472
rect 40532 9469 40544 9472
rect 40578 9500 40590 9503
rect 41325 9503 41383 9509
rect 41325 9500 41337 9503
rect 40578 9472 41337 9500
rect 40578 9469 40590 9472
rect 40532 9463 40590 9469
rect 41325 9469 41337 9472
rect 41371 9469 41383 9503
rect 41325 9463 41383 9469
rect 30006 9432 30012 9444
rect 27203 9404 30012 9432
rect 27203 9401 27215 9404
rect 27157 9395 27215 9401
rect 30006 9392 30012 9404
rect 30064 9392 30070 9444
rect 30374 9392 30380 9444
rect 30432 9432 30438 9444
rect 30432 9404 33088 9432
rect 30432 9392 30438 9404
rect 33060 9376 33088 9404
rect 35710 9392 35716 9444
rect 35768 9432 35774 9444
rect 36126 9435 36184 9441
rect 36126 9432 36138 9435
rect 35768 9404 36138 9432
rect 35768 9392 35774 9404
rect 36126 9401 36138 9404
rect 36172 9401 36184 9435
rect 42613 9435 42671 9441
rect 42613 9432 42625 9435
rect 36126 9395 36184 9401
rect 42260 9404 42625 9432
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 19978 9364 19984 9376
rect 19843 9336 19984 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 21450 9324 21456 9376
rect 21508 9364 21514 9376
rect 21545 9367 21603 9373
rect 21545 9364 21557 9367
rect 21508 9336 21557 9364
rect 21508 9324 21514 9336
rect 21545 9333 21557 9336
rect 21591 9333 21603 9367
rect 21545 9327 21603 9333
rect 22695 9367 22753 9373
rect 22695 9333 22707 9367
rect 22741 9364 22753 9367
rect 22922 9364 22928 9376
rect 22741 9336 22928 9364
rect 22741 9333 22753 9336
rect 22695 9327 22753 9333
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 23106 9364 23112 9376
rect 23067 9336 23112 9364
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 23842 9364 23848 9376
rect 23803 9336 23848 9364
rect 23842 9324 23848 9336
rect 23900 9324 23906 9376
rect 24854 9364 24860 9376
rect 24815 9336 24860 9364
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 27062 9324 27068 9376
rect 27120 9364 27126 9376
rect 27433 9367 27491 9373
rect 27433 9364 27445 9367
rect 27120 9336 27445 9364
rect 27120 9324 27126 9336
rect 27433 9333 27445 9336
rect 27479 9333 27491 9367
rect 27433 9327 27491 9333
rect 27522 9324 27528 9376
rect 27580 9364 27586 9376
rect 27709 9367 27767 9373
rect 27709 9364 27721 9367
rect 27580 9336 27721 9364
rect 27580 9324 27586 9336
rect 27709 9333 27721 9336
rect 27755 9333 27767 9367
rect 27709 9327 27767 9333
rect 29549 9367 29607 9373
rect 29549 9333 29561 9367
rect 29595 9364 29607 9367
rect 29638 9364 29644 9376
rect 29595 9336 29644 9364
rect 29595 9333 29607 9336
rect 29549 9327 29607 9333
rect 29638 9324 29644 9336
rect 29696 9324 29702 9376
rect 32033 9367 32091 9373
rect 32033 9333 32045 9367
rect 32079 9364 32091 9367
rect 32582 9364 32588 9376
rect 32079 9336 32588 9364
rect 32079 9333 32091 9336
rect 32033 9327 32091 9333
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 33042 9364 33048 9376
rect 32955 9336 33048 9364
rect 33042 9324 33048 9336
rect 33100 9324 33106 9376
rect 36725 9367 36783 9373
rect 36725 9333 36737 9367
rect 36771 9364 36783 9367
rect 36906 9364 36912 9376
rect 36771 9336 36912 9364
rect 36771 9333 36783 9336
rect 36725 9327 36783 9333
rect 36906 9324 36912 9336
rect 36964 9324 36970 9376
rect 37734 9364 37740 9376
rect 37695 9336 37740 9364
rect 37734 9324 37740 9336
rect 37792 9324 37798 9376
rect 42150 9324 42156 9376
rect 42208 9364 42214 9376
rect 42260 9373 42288 9404
rect 42613 9401 42625 9404
rect 42659 9432 42671 9435
rect 43809 9435 43867 9441
rect 43809 9432 43821 9435
rect 42659 9404 42794 9432
rect 42659 9401 42671 9404
rect 42613 9395 42671 9401
rect 42245 9367 42303 9373
rect 42245 9364 42257 9367
rect 42208 9336 42257 9364
rect 42208 9324 42214 9336
rect 42245 9333 42257 9336
rect 42291 9333 42303 9367
rect 42766 9364 42794 9404
rect 43364 9404 43821 9432
rect 43364 9364 43392 9404
rect 43809 9401 43821 9404
rect 43855 9401 43867 9435
rect 44082 9432 44088 9444
rect 44043 9404 44088 9432
rect 43809 9395 43867 9401
rect 42766 9336 43392 9364
rect 43824 9364 43852 9395
rect 44082 9392 44088 9404
rect 44140 9392 44146 9444
rect 44177 9435 44235 9441
rect 44177 9401 44189 9435
rect 44223 9401 44235 9435
rect 44177 9395 44235 9401
rect 46293 9435 46351 9441
rect 46293 9401 46305 9435
rect 46339 9401 46351 9435
rect 46842 9432 46848 9444
rect 46803 9404 46848 9432
rect 46293 9395 46351 9401
rect 44192 9364 44220 9395
rect 43824 9336 44220 9364
rect 42245 9327 42303 9333
rect 45922 9324 45928 9376
rect 45980 9364 45986 9376
rect 46308 9364 46336 9395
rect 46842 9392 46848 9404
rect 46900 9392 46906 9444
rect 45980 9336 46336 9364
rect 45980 9324 45986 9336
rect 1104 9274 48852 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 48852 9274
rect 1104 9200 48852 9222
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 17862 9160 17868 9172
rect 17635 9132 17868 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18831 9163 18889 9169
rect 18831 9160 18843 9163
rect 18012 9132 18843 9160
rect 18012 9120 18018 9132
rect 18831 9129 18843 9132
rect 18877 9129 18889 9163
rect 18831 9123 18889 9129
rect 19889 9163 19947 9169
rect 19889 9129 19901 9163
rect 19935 9160 19947 9163
rect 20162 9160 20168 9172
rect 19935 9132 20168 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 24210 9160 24216 9172
rect 24171 9132 24216 9160
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 25682 9120 25688 9172
rect 25740 9160 25746 9172
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 25740 9132 25789 9160
rect 25740 9120 25746 9132
rect 25777 9129 25789 9132
rect 25823 9129 25835 9163
rect 26234 9160 26240 9172
rect 26195 9132 26240 9160
rect 25777 9123 25835 9129
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 27801 9163 27859 9169
rect 27801 9129 27813 9163
rect 27847 9160 27859 9163
rect 27982 9160 27988 9172
rect 27847 9132 27988 9160
rect 27847 9129 27859 9132
rect 27801 9123 27859 9129
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 28166 9160 28172 9172
rect 28127 9132 28172 9160
rect 28166 9120 28172 9132
rect 28224 9120 28230 9172
rect 30607 9163 30665 9169
rect 30607 9129 30619 9163
rect 30653 9160 30665 9163
rect 30834 9160 30840 9172
rect 30653 9132 30840 9160
rect 30653 9129 30665 9132
rect 30607 9123 30665 9129
rect 30834 9120 30840 9132
rect 30892 9120 30898 9172
rect 35526 9160 35532 9172
rect 35487 9132 35532 9160
rect 35526 9120 35532 9132
rect 35584 9120 35590 9172
rect 35618 9120 35624 9172
rect 35676 9160 35682 9172
rect 35805 9163 35863 9169
rect 35805 9160 35817 9163
rect 35676 9132 35817 9160
rect 35676 9120 35682 9132
rect 35805 9129 35817 9132
rect 35851 9129 35863 9163
rect 35805 9123 35863 9129
rect 38010 9120 38016 9172
rect 38068 9160 38074 9172
rect 38105 9163 38163 9169
rect 38105 9160 38117 9163
rect 38068 9132 38117 9160
rect 38068 9120 38074 9132
rect 38105 9129 38117 9132
rect 38151 9129 38163 9163
rect 39850 9160 39856 9172
rect 39811 9132 39856 9160
rect 38105 9123 38163 9129
rect 39850 9120 39856 9132
rect 39908 9120 39914 9172
rect 41601 9163 41659 9169
rect 41601 9129 41613 9163
rect 41647 9160 41659 9163
rect 41782 9160 41788 9172
rect 41647 9132 41788 9160
rect 41647 9129 41659 9132
rect 41601 9123 41659 9129
rect 41782 9120 41788 9132
rect 41840 9120 41846 9172
rect 42518 9120 42524 9172
rect 42576 9160 42582 9172
rect 42705 9163 42763 9169
rect 42705 9160 42717 9163
rect 42576 9132 42717 9160
rect 42576 9120 42582 9132
rect 42705 9129 42717 9132
rect 42751 9129 42763 9163
rect 42705 9123 42763 9129
rect 44082 9120 44088 9172
rect 44140 9160 44146 9172
rect 44453 9163 44511 9169
rect 44453 9160 44465 9163
rect 44140 9132 44465 9160
rect 44140 9120 44146 9132
rect 44453 9129 44465 9132
rect 44499 9160 44511 9163
rect 47351 9163 47409 9169
rect 47351 9160 47363 9163
rect 44499 9132 47363 9160
rect 44499 9129 44511 9132
rect 44453 9123 44511 9129
rect 47351 9129 47363 9132
rect 47397 9129 47409 9163
rect 47351 9123 47409 9129
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 26875 9095 26933 9101
rect 18656 9064 21036 9092
rect 18656 9052 18662 9064
rect 18690 9024 18696 9036
rect 18651 8996 18696 9024
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 18840 8996 19717 9024
rect 18840 8984 18846 8996
rect 19705 8993 19717 8996
rect 19751 9024 19763 9027
rect 20070 9024 20076 9036
rect 19751 8996 20076 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 21008 9033 21036 9064
rect 26875 9061 26887 9095
rect 26921 9092 26933 9095
rect 27062 9092 27068 9104
rect 26921 9064 27068 9092
rect 26921 9061 26933 9064
rect 26875 9055 26933 9061
rect 27062 9052 27068 9064
rect 27120 9052 27126 9104
rect 20993 9027 21051 9033
rect 20993 8993 21005 9027
rect 21039 9024 21051 9027
rect 21634 9024 21640 9036
rect 21039 8996 21640 9024
rect 21039 8993 21051 8996
rect 20993 8987 21051 8993
rect 21634 8984 21640 8996
rect 21692 8984 21698 9036
rect 22738 8984 22744 9036
rect 22796 9024 22802 9036
rect 23201 9027 23259 9033
rect 23201 9024 23213 9027
rect 22796 8996 23213 9024
rect 22796 8984 22802 8996
rect 23201 8993 23213 8996
rect 23247 8993 23259 9027
rect 23201 8987 23259 8993
rect 24026 8984 24032 9036
rect 24084 9024 24090 9036
rect 24708 9027 24766 9033
rect 24708 9024 24720 9027
rect 24084 8996 24720 9024
rect 24084 8984 24090 8996
rect 24708 8993 24720 8996
rect 24754 9024 24766 9027
rect 24946 9024 24952 9036
rect 24754 8996 24952 9024
rect 24754 8993 24766 8996
rect 24708 8987 24766 8993
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 28810 8984 28816 9036
rect 28868 9024 28874 9036
rect 28905 9027 28963 9033
rect 28905 9024 28917 9027
rect 28868 8996 28917 9024
rect 28868 8984 28874 8996
rect 28905 8993 28917 8996
rect 28951 8993 28963 9027
rect 28905 8987 28963 8993
rect 29270 8984 29276 9036
rect 29328 9024 29334 9036
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 29328 8996 29377 9024
rect 29328 8984 29334 8996
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 29365 8987 29423 8993
rect 30536 9027 30594 9033
rect 30536 8993 30548 9027
rect 30582 9024 30594 9027
rect 30834 9024 30840 9036
rect 30582 8996 30840 9024
rect 30582 8993 30594 8996
rect 30536 8987 30594 8993
rect 30834 8984 30840 8996
rect 30892 9024 30898 9036
rect 32122 9024 32128 9036
rect 30892 8996 32128 9024
rect 30892 8984 30898 8996
rect 32122 8984 32128 8996
rect 32180 8984 32186 9036
rect 32582 9024 32588 9036
rect 32543 8996 32588 9024
rect 32582 8984 32588 8996
rect 32640 8984 32646 9036
rect 32950 8984 32956 9036
rect 33008 9024 33014 9036
rect 33045 9027 33103 9033
rect 33045 9024 33057 9027
rect 33008 8996 33057 9024
rect 33008 8984 33014 8996
rect 33045 8993 33057 8996
rect 33091 8993 33103 9027
rect 33045 8987 33103 8993
rect 33410 8984 33416 9036
rect 33468 9024 33474 9036
rect 34422 9024 34428 9036
rect 33468 8996 34428 9024
rect 33468 8984 33474 8996
rect 34422 8984 34428 8996
rect 34480 8984 34486 9036
rect 34977 9027 35035 9033
rect 34977 8993 34989 9027
rect 35023 9024 35035 9027
rect 35544 9024 35572 9120
rect 41874 9092 41880 9104
rect 41835 9064 41880 9092
rect 41874 9052 41880 9064
rect 41932 9052 41938 9104
rect 42429 9095 42487 9101
rect 42429 9061 42441 9095
rect 42475 9092 42487 9095
rect 43254 9092 43260 9104
rect 42475 9064 43260 9092
rect 42475 9061 42487 9064
rect 42429 9055 42487 9061
rect 43254 9052 43260 9064
rect 43312 9052 43318 9104
rect 43530 9092 43536 9104
rect 43491 9064 43536 9092
rect 43530 9052 43536 9064
rect 43588 9052 43594 9104
rect 45833 9095 45891 9101
rect 45833 9061 45845 9095
rect 45879 9092 45891 9095
rect 46106 9092 46112 9104
rect 45879 9064 46112 9092
rect 45879 9061 45891 9064
rect 45833 9055 45891 9061
rect 46106 9052 46112 9064
rect 46164 9052 46170 9104
rect 36078 9024 36084 9036
rect 35023 8996 35572 9024
rect 36039 8996 36084 9024
rect 35023 8993 35035 8996
rect 34977 8987 35035 8993
rect 36078 8984 36084 8996
rect 36136 8984 36142 9036
rect 36354 8984 36360 9036
rect 36412 9024 36418 9036
rect 36541 9027 36599 9033
rect 36541 9024 36553 9027
rect 36412 8996 36553 9024
rect 36412 8984 36418 8996
rect 36541 8993 36553 8996
rect 36587 8993 36599 9027
rect 47210 9024 47216 9036
rect 47171 8996 47216 9024
rect 36541 8987 36599 8993
rect 47210 8984 47216 8996
rect 47268 8984 47274 9036
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 25038 8956 25044 8968
rect 23891 8928 25044 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 26510 8956 26516 8968
rect 26471 8928 26516 8956
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 29546 8916 29552 8968
rect 29604 8956 29610 8968
rect 29641 8959 29699 8965
rect 29641 8956 29653 8959
rect 29604 8928 29653 8956
rect 29604 8916 29610 8928
rect 29641 8925 29653 8928
rect 29687 8956 29699 8959
rect 29917 8959 29975 8965
rect 29917 8956 29929 8959
rect 29687 8928 29929 8956
rect 29687 8925 29699 8928
rect 29641 8919 29699 8925
rect 29917 8925 29929 8928
rect 29963 8925 29975 8959
rect 29917 8919 29975 8925
rect 33321 8959 33379 8965
rect 33321 8925 33333 8959
rect 33367 8956 33379 8959
rect 34790 8956 34796 8968
rect 33367 8928 34796 8956
rect 33367 8925 33379 8928
rect 33321 8919 33379 8925
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 35161 8959 35219 8965
rect 35161 8925 35173 8959
rect 35207 8956 35219 8959
rect 36722 8956 36728 8968
rect 35207 8928 36728 8956
rect 35207 8925 35219 8928
rect 35161 8919 35219 8925
rect 36722 8916 36728 8928
rect 36780 8916 36786 8968
rect 36817 8959 36875 8965
rect 36817 8925 36829 8959
rect 36863 8956 36875 8959
rect 37737 8959 37795 8965
rect 37737 8956 37749 8959
rect 36863 8928 37749 8956
rect 36863 8925 36875 8928
rect 36817 8919 36875 8925
rect 37737 8925 37749 8928
rect 37783 8956 37795 8959
rect 38102 8956 38108 8968
rect 37783 8928 38108 8956
rect 37783 8925 37795 8928
rect 37737 8919 37795 8925
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 39482 8956 39488 8968
rect 39443 8928 39488 8956
rect 39482 8916 39488 8928
rect 39540 8916 39546 8968
rect 41782 8956 41788 8968
rect 41743 8928 41788 8956
rect 41782 8916 41788 8928
rect 41840 8956 41846 8968
rect 43438 8956 43444 8968
rect 41840 8928 42794 8956
rect 43399 8928 43444 8956
rect 41840 8916 41846 8928
rect 40405 8891 40463 8897
rect 40405 8857 40417 8891
rect 40451 8888 40463 8891
rect 42766 8888 42794 8928
rect 43438 8916 43444 8928
rect 43496 8916 43502 8968
rect 43714 8956 43720 8968
rect 43675 8928 43720 8956
rect 43714 8916 43720 8928
rect 43772 8916 43778 8968
rect 45738 8956 45744 8968
rect 45699 8928 45744 8956
rect 45738 8916 45744 8928
rect 45796 8916 45802 8968
rect 46014 8956 46020 8968
rect 45975 8928 46020 8956
rect 46014 8916 46020 8928
rect 46072 8956 46078 8968
rect 46842 8956 46848 8968
rect 46072 8928 46848 8956
rect 46072 8916 46078 8928
rect 46842 8916 46848 8928
rect 46900 8916 46906 8968
rect 47486 8888 47492 8900
rect 40451 8860 42355 8888
rect 42766 8860 47492 8888
rect 40451 8857 40463 8860
rect 40405 8851 40463 8857
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24811 8823 24869 8829
rect 24811 8820 24823 8823
rect 23992 8792 24823 8820
rect 23992 8780 23998 8792
rect 24811 8789 24823 8792
rect 24857 8789 24869 8823
rect 24811 8783 24869 8789
rect 27433 8823 27491 8829
rect 27433 8789 27445 8823
rect 27479 8820 27491 8823
rect 27614 8820 27620 8832
rect 27479 8792 27620 8820
rect 27479 8789 27491 8792
rect 27433 8783 27491 8789
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 33686 8820 33692 8832
rect 33647 8792 33692 8820
rect 33686 8780 33692 8792
rect 33744 8780 33750 8832
rect 38654 8820 38660 8832
rect 38615 8792 38660 8820
rect 38654 8780 38660 8792
rect 38712 8780 38718 8832
rect 42327 8820 42355 8860
rect 47486 8848 47492 8860
rect 47544 8848 47550 8900
rect 45922 8820 45928 8832
rect 42327 8792 45928 8820
rect 45922 8780 45928 8792
rect 45980 8780 45986 8832
rect 1104 8730 48852 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 48852 8730
rect 1104 8656 48852 8678
rect 20070 8616 20076 8628
rect 20031 8588 20076 8616
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 21634 8616 21640 8628
rect 21595 8588 21640 8616
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 22465 8619 22523 8625
rect 22465 8585 22477 8619
rect 22511 8616 22523 8619
rect 22738 8616 22744 8628
rect 22511 8588 22744 8616
rect 22511 8585 22523 8588
rect 22465 8579 22523 8585
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 24673 8619 24731 8625
rect 24673 8616 24685 8619
rect 23164 8588 24685 8616
rect 23164 8576 23170 8588
rect 24673 8585 24685 8588
rect 24719 8585 24731 8619
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24673 8579 24731 8585
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27341 8579 27399 8585
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 27663 8619 27721 8625
rect 27663 8616 27675 8619
rect 27488 8588 27675 8616
rect 27488 8576 27494 8588
rect 27663 8585 27675 8588
rect 27709 8585 27721 8619
rect 27663 8579 27721 8585
rect 28721 8619 28779 8625
rect 28721 8585 28733 8619
rect 28767 8616 28779 8619
rect 28810 8616 28816 8628
rect 28767 8588 28816 8616
rect 28767 8585 28779 8588
rect 28721 8579 28779 8585
rect 28810 8576 28816 8588
rect 28868 8576 28874 8628
rect 30834 8616 30840 8628
rect 30795 8588 30840 8616
rect 30834 8576 30840 8588
rect 30892 8576 30898 8628
rect 32582 8616 32588 8628
rect 32543 8588 32588 8616
rect 32582 8576 32588 8588
rect 32640 8576 32646 8628
rect 33042 8616 33048 8628
rect 33003 8588 33048 8616
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 34422 8616 34428 8628
rect 34383 8588 34428 8616
rect 34422 8576 34428 8588
rect 34480 8576 34486 8628
rect 38102 8616 38108 8628
rect 38063 8588 38108 8616
rect 38102 8576 38108 8588
rect 38160 8576 38166 8628
rect 40957 8619 41015 8625
rect 40957 8585 40969 8619
rect 41003 8616 41015 8619
rect 41782 8616 41788 8628
rect 41003 8588 41788 8616
rect 41003 8585 41015 8588
rect 40957 8579 41015 8585
rect 41782 8576 41788 8588
rect 41840 8576 41846 8628
rect 41874 8576 41880 8628
rect 41932 8616 41938 8628
rect 42429 8619 42487 8625
rect 42429 8616 42441 8619
rect 41932 8588 42441 8616
rect 41932 8576 41938 8588
rect 42429 8585 42441 8588
rect 42475 8616 42487 8619
rect 43530 8616 43536 8628
rect 42475 8588 43536 8616
rect 42475 8585 42487 8588
rect 42429 8579 42487 8585
rect 43530 8576 43536 8588
rect 43588 8616 43594 8628
rect 43625 8619 43683 8625
rect 43625 8616 43637 8619
rect 43588 8588 43637 8616
rect 43588 8576 43594 8588
rect 43625 8585 43637 8588
rect 43671 8585 43683 8619
rect 43625 8579 43683 8585
rect 45373 8619 45431 8625
rect 45373 8585 45385 8619
rect 45419 8616 45431 8619
rect 45738 8616 45744 8628
rect 45419 8588 45744 8616
rect 45419 8585 45431 8588
rect 45373 8579 45431 8585
rect 45738 8576 45744 8588
rect 45796 8576 45802 8628
rect 23017 8551 23075 8557
rect 23017 8517 23029 8551
rect 23063 8548 23075 8551
rect 24026 8548 24032 8560
rect 23063 8520 24032 8548
rect 23063 8517 23075 8520
rect 23017 8511 23075 8517
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18690 8480 18696 8492
rect 18647 8452 18696 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18690 8440 18696 8452
rect 18748 8480 18754 8492
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 18748 8452 19809 8480
rect 18748 8440 18754 8452
rect 19797 8449 19809 8452
rect 19843 8480 19855 8483
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 19843 8452 21005 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 22557 8415 22615 8421
rect 22557 8381 22569 8415
rect 22603 8412 22615 8415
rect 23032 8412 23060 8511
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 25682 8508 25688 8560
rect 25740 8548 25746 8560
rect 28261 8551 28319 8557
rect 28261 8548 28273 8551
rect 25740 8520 28273 8548
rect 25740 8508 25746 8520
rect 28261 8517 28273 8520
rect 28307 8548 28319 8551
rect 28442 8548 28448 8560
rect 28307 8520 28448 8548
rect 28307 8517 28319 8520
rect 28261 8511 28319 8517
rect 28442 8508 28448 8520
rect 28500 8548 28506 8560
rect 29270 8548 29276 8560
rect 28500 8520 29276 8548
rect 28500 8508 28506 8520
rect 29270 8508 29276 8520
rect 29328 8508 29334 8560
rect 31205 8551 31263 8557
rect 31205 8517 31217 8551
rect 31251 8548 31263 8551
rect 31570 8548 31576 8560
rect 31251 8520 31576 8548
rect 31251 8517 31263 8520
rect 31205 8511 31263 8517
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 23842 8480 23848 8492
rect 23799 8452 23848 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 23842 8440 23848 8452
rect 23900 8440 23906 8492
rect 29546 8480 29552 8492
rect 29507 8452 29552 8480
rect 29546 8440 29552 8452
rect 29604 8440 29610 8492
rect 22603 8384 23060 8412
rect 27592 8415 27650 8421
rect 22603 8381 22615 8384
rect 22557 8375 22615 8381
rect 27592 8381 27604 8415
rect 27638 8412 27650 8415
rect 28350 8412 28356 8424
rect 27638 8384 28356 8412
rect 27638 8381 27650 8384
rect 27592 8375 27650 8381
rect 28350 8372 28356 8384
rect 28408 8372 28414 8424
rect 28994 8412 29000 8424
rect 28966 8372 29000 8412
rect 29052 8412 29058 8424
rect 31220 8412 31248 8511
rect 31570 8508 31576 8520
rect 31628 8508 31634 8560
rect 39758 8508 39764 8560
rect 39816 8548 39822 8560
rect 42245 8551 42303 8557
rect 42245 8548 42257 8551
rect 39816 8520 42257 8548
rect 39816 8508 39822 8520
rect 42245 8517 42257 8520
rect 42291 8517 42303 8551
rect 42245 8511 42303 8517
rect 43073 8551 43131 8557
rect 43073 8517 43085 8551
rect 43119 8548 43131 8551
rect 43438 8548 43444 8560
rect 43119 8520 43444 8548
rect 43119 8517 43131 8520
rect 43073 8511 43131 8517
rect 43438 8508 43444 8520
rect 43496 8548 43502 8560
rect 46290 8548 46296 8560
rect 43496 8520 46296 8548
rect 43496 8508 43502 8520
rect 46290 8508 46296 8520
rect 46348 8508 46354 8560
rect 31386 8480 31392 8492
rect 31347 8452 31392 8480
rect 31386 8440 31392 8452
rect 31444 8440 31450 8492
rect 31478 8440 31484 8492
rect 31536 8480 31542 8492
rect 31665 8483 31723 8489
rect 31665 8480 31677 8483
rect 31536 8452 31677 8480
rect 31536 8440 31542 8452
rect 31665 8449 31677 8452
rect 31711 8449 31723 8483
rect 31665 8443 31723 8449
rect 33686 8440 33692 8492
rect 33744 8480 33750 8492
rect 35621 8483 35679 8489
rect 33744 8452 35480 8480
rect 33744 8440 33750 8452
rect 29052 8384 31248 8412
rect 29052 8372 29058 8384
rect 33042 8372 33048 8424
rect 33100 8412 33106 8424
rect 33796 8421 33824 8452
rect 33229 8415 33287 8421
rect 33229 8412 33241 8415
rect 33100 8384 33241 8412
rect 33100 8372 33106 8384
rect 33229 8381 33241 8384
rect 33275 8381 33287 8415
rect 33229 8375 33287 8381
rect 33781 8415 33839 8421
rect 33781 8381 33793 8415
rect 33827 8381 33839 8415
rect 33781 8375 33839 8381
rect 34330 8372 34336 8424
rect 34388 8412 34394 8424
rect 34882 8412 34888 8424
rect 34388 8384 34888 8412
rect 34388 8372 34394 8384
rect 34882 8372 34888 8384
rect 34940 8372 34946 8424
rect 35452 8421 35480 8452
rect 35621 8449 35633 8483
rect 35667 8480 35679 8483
rect 39482 8480 39488 8492
rect 35667 8452 39488 8480
rect 35667 8449 35679 8452
rect 35621 8443 35679 8449
rect 39482 8440 39488 8452
rect 39540 8480 39546 8492
rect 40221 8483 40279 8489
rect 40221 8480 40233 8483
rect 39540 8452 40233 8480
rect 39540 8440 39546 8452
rect 40221 8449 40233 8452
rect 40267 8449 40279 8483
rect 40221 8443 40279 8449
rect 42153 8483 42211 8489
rect 42153 8449 42165 8483
rect 42199 8480 42211 8483
rect 43714 8480 43720 8492
rect 42199 8452 43720 8480
rect 42199 8449 42211 8452
rect 42153 8443 42211 8449
rect 43714 8440 43720 8452
rect 43772 8440 43778 8492
rect 45741 8483 45799 8489
rect 45741 8449 45753 8483
rect 45787 8480 45799 8483
rect 46106 8480 46112 8492
rect 45787 8452 46112 8480
rect 45787 8449 45799 8452
rect 45741 8443 45799 8449
rect 46106 8440 46112 8452
rect 46164 8440 46170 8492
rect 35437 8415 35495 8421
rect 35437 8381 35449 8415
rect 35483 8412 35495 8415
rect 35526 8412 35532 8424
rect 35483 8384 35532 8412
rect 35483 8381 35495 8384
rect 35437 8375 35495 8381
rect 35526 8372 35532 8384
rect 35584 8372 35590 8424
rect 36630 8372 36636 8424
rect 36688 8412 36694 8424
rect 36725 8415 36783 8421
rect 36725 8412 36737 8415
rect 36688 8384 36737 8412
rect 36688 8372 36694 8384
rect 36725 8381 36737 8384
rect 36771 8381 36783 8415
rect 36725 8375 36783 8381
rect 36814 8372 36820 8424
rect 36872 8412 36878 8424
rect 37185 8415 37243 8421
rect 37185 8412 37197 8415
rect 36872 8384 37197 8412
rect 36872 8372 36878 8384
rect 37185 8381 37197 8384
rect 37231 8381 37243 8415
rect 37185 8375 37243 8381
rect 38657 8415 38715 8421
rect 38657 8381 38669 8415
rect 38703 8381 38715 8415
rect 38657 8375 38715 8381
rect 19150 8344 19156 8356
rect 19111 8316 19156 8344
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8344 19303 8347
rect 19426 8344 19432 8356
rect 19291 8316 19432 8344
rect 19291 8313 19303 8316
rect 19245 8307 19303 8313
rect 18969 8279 19027 8285
rect 18969 8245 18981 8279
rect 19015 8276 19027 8279
rect 19260 8276 19288 8307
rect 19426 8304 19432 8316
rect 19484 8304 19490 8356
rect 20714 8344 20720 8356
rect 20675 8316 20720 8344
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 20809 8347 20867 8353
rect 20809 8313 20821 8347
rect 20855 8344 20867 8347
rect 20898 8344 20904 8356
rect 20855 8316 20904 8344
rect 20855 8313 20867 8316
rect 20809 8307 20867 8313
rect 19015 8248 19288 8276
rect 20533 8279 20591 8285
rect 19015 8245 19027 8248
rect 18969 8239 19027 8245
rect 20533 8245 20545 8279
rect 20579 8276 20591 8279
rect 20824 8276 20852 8307
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 23385 8347 23443 8353
rect 23385 8313 23397 8347
rect 23431 8344 23443 8347
rect 23566 8344 23572 8356
rect 23431 8316 23572 8344
rect 23431 8313 23443 8316
rect 23385 8307 23443 8313
rect 23566 8304 23572 8316
rect 23624 8344 23630 8356
rect 24074 8347 24132 8353
rect 24074 8344 24086 8347
rect 23624 8316 24086 8344
rect 23624 8304 23630 8316
rect 24074 8313 24086 8316
rect 24120 8313 24132 8347
rect 26050 8344 26056 8356
rect 26011 8316 26056 8344
rect 24074 8307 24132 8313
rect 26050 8304 26056 8316
rect 26108 8304 26114 8356
rect 26145 8347 26203 8353
rect 26145 8313 26157 8347
rect 26191 8313 26203 8347
rect 26694 8344 26700 8356
rect 26655 8316 26700 8344
rect 26145 8307 26203 8313
rect 20579 8248 20852 8276
rect 20579 8245 20591 8248
rect 20533 8239 20591 8245
rect 23658 8236 23664 8288
rect 23716 8276 23722 8288
rect 25869 8279 25927 8285
rect 25869 8276 25881 8279
rect 23716 8248 25881 8276
rect 23716 8236 23722 8248
rect 25869 8245 25881 8248
rect 25915 8276 25927 8279
rect 26160 8276 26188 8307
rect 26694 8304 26700 8316
rect 26752 8304 26758 8356
rect 28966 8344 28994 8372
rect 26804 8316 28994 8344
rect 29089 8347 29147 8353
rect 26804 8276 26832 8316
rect 29089 8313 29101 8347
rect 29135 8344 29147 8347
rect 29911 8347 29969 8353
rect 29911 8344 29923 8347
rect 29135 8316 29923 8344
rect 29135 8313 29147 8316
rect 29089 8307 29147 8313
rect 29911 8313 29923 8316
rect 29957 8344 29969 8347
rect 30282 8344 30288 8356
rect 29957 8316 30288 8344
rect 29957 8313 29969 8316
rect 29911 8307 29969 8313
rect 27062 8276 27068 8288
rect 25915 8248 26832 8276
rect 26975 8248 27068 8276
rect 25915 8245 25927 8248
rect 25869 8239 25927 8245
rect 27062 8236 27068 8248
rect 27120 8276 27126 8288
rect 29104 8276 29132 8307
rect 30282 8304 30288 8316
rect 30340 8304 30346 8356
rect 31481 8347 31539 8353
rect 31481 8313 31493 8347
rect 31527 8344 31539 8347
rect 31570 8344 31576 8356
rect 31527 8316 31576 8344
rect 31527 8313 31539 8316
rect 31481 8307 31539 8313
rect 31570 8304 31576 8316
rect 31628 8304 31634 8356
rect 33965 8347 34023 8353
rect 33965 8313 33977 8347
rect 34011 8344 34023 8347
rect 38672 8344 38700 8375
rect 39114 8372 39120 8424
rect 39172 8412 39178 8424
rect 41233 8415 41291 8421
rect 41233 8412 41245 8415
rect 39172 8384 41245 8412
rect 39172 8372 39178 8384
rect 41233 8381 41245 8384
rect 41279 8381 41291 8415
rect 41233 8375 41291 8381
rect 42245 8415 42303 8421
rect 42245 8381 42257 8415
rect 42291 8412 42303 8415
rect 43200 8415 43258 8421
rect 43200 8412 43212 8415
rect 42291 8384 43212 8412
rect 42291 8381 42303 8384
rect 42245 8375 42303 8381
rect 43200 8381 43212 8384
rect 43246 8381 43258 8415
rect 43200 8375 43258 8381
rect 43303 8415 43361 8421
rect 43303 8381 43315 8415
rect 43349 8412 43361 8415
rect 44266 8412 44272 8424
rect 43349 8384 44272 8412
rect 43349 8381 43361 8384
rect 43303 8375 43361 8381
rect 38746 8344 38752 8356
rect 34011 8316 38752 8344
rect 34011 8313 34023 8316
rect 33965 8307 34023 8313
rect 38746 8304 38752 8316
rect 38804 8304 38810 8356
rect 39019 8347 39077 8353
rect 39019 8344 39031 8347
rect 38856 8316 39031 8344
rect 30466 8276 30472 8288
rect 27120 8248 29132 8276
rect 30427 8248 30472 8276
rect 27120 8236 27126 8248
rect 30466 8236 30472 8248
rect 30524 8236 30530 8288
rect 36078 8276 36084 8288
rect 36039 8248 36084 8276
rect 36078 8236 36084 8248
rect 36136 8276 36142 8288
rect 36541 8279 36599 8285
rect 36541 8276 36553 8279
rect 36136 8248 36553 8276
rect 36136 8236 36142 8248
rect 36541 8245 36553 8248
rect 36587 8276 36599 8279
rect 36630 8276 36636 8288
rect 36587 8248 36636 8276
rect 36587 8245 36599 8248
rect 36541 8239 36599 8245
rect 36630 8236 36636 8248
rect 36688 8236 36694 8288
rect 36998 8276 37004 8288
rect 36959 8248 37004 8276
rect 36998 8236 37004 8248
rect 37056 8236 37062 8288
rect 37829 8279 37887 8285
rect 37829 8245 37841 8279
rect 37875 8276 37887 8279
rect 38010 8276 38016 8288
rect 37875 8248 38016 8276
rect 37875 8245 37887 8248
rect 37829 8239 37887 8245
rect 38010 8236 38016 8248
rect 38068 8276 38074 8288
rect 38565 8279 38623 8285
rect 38565 8276 38577 8279
rect 38068 8248 38577 8276
rect 38068 8236 38074 8248
rect 38565 8245 38577 8248
rect 38611 8276 38623 8279
rect 38856 8276 38884 8316
rect 39019 8313 39031 8316
rect 39065 8344 39077 8347
rect 39065 8316 39896 8344
rect 39065 8313 39077 8316
rect 39019 8307 39077 8313
rect 39868 8288 39896 8316
rect 39574 8276 39580 8288
rect 38611 8248 38884 8276
rect 39535 8248 39580 8276
rect 38611 8245 38623 8248
rect 38565 8239 38623 8245
rect 39574 8236 39580 8248
rect 39632 8236 39638 8288
rect 39850 8276 39856 8288
rect 39811 8248 39856 8276
rect 39850 8236 39856 8248
rect 39908 8236 39914 8288
rect 41248 8276 41276 8375
rect 41506 8344 41512 8356
rect 41467 8316 41512 8344
rect 41506 8304 41512 8316
rect 41564 8304 41570 8356
rect 41601 8347 41659 8353
rect 41601 8313 41613 8347
rect 41647 8344 41659 8347
rect 42150 8344 42156 8356
rect 41647 8316 42156 8344
rect 41647 8313 41659 8316
rect 41601 8307 41659 8313
rect 41616 8276 41644 8307
rect 42150 8304 42156 8316
rect 42208 8304 42214 8356
rect 43215 8344 43243 8375
rect 44266 8372 44272 8384
rect 44324 8372 44330 8424
rect 46198 8412 46204 8424
rect 46159 8384 46204 8412
rect 46198 8372 46204 8384
rect 46256 8372 46262 8424
rect 43806 8344 43812 8356
rect 43215 8316 43812 8344
rect 43806 8304 43812 8316
rect 43864 8344 43870 8356
rect 43993 8347 44051 8353
rect 43993 8344 44005 8347
rect 43864 8316 44005 8344
rect 43864 8304 43870 8316
rect 43993 8313 44005 8316
rect 44039 8313 44051 8347
rect 46106 8344 46112 8356
rect 46067 8316 46112 8344
rect 43993 8307 44051 8313
rect 46106 8304 46112 8316
rect 46164 8304 46170 8356
rect 41248 8248 41644 8276
rect 44358 8236 44364 8288
rect 44416 8276 44422 8288
rect 44453 8279 44511 8285
rect 44453 8276 44465 8279
rect 44416 8248 44465 8276
rect 44416 8236 44422 8248
rect 44453 8245 44465 8248
rect 44499 8245 44511 8279
rect 47210 8276 47216 8288
rect 47171 8248 47216 8276
rect 44453 8239 44511 8245
rect 47210 8236 47216 8248
rect 47268 8236 47274 8288
rect 1104 8186 48852 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 48852 8186
rect 1104 8112 48852 8134
rect 23658 8072 23664 8084
rect 23619 8044 23664 8072
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 23842 8032 23848 8084
rect 23900 8072 23906 8084
rect 24213 8075 24271 8081
rect 24213 8072 24225 8075
rect 23900 8044 24225 8072
rect 23900 8032 23906 8044
rect 24213 8041 24225 8044
rect 24259 8041 24271 8075
rect 24213 8035 24271 8041
rect 27617 8075 27675 8081
rect 27617 8041 27629 8075
rect 27663 8072 27675 8075
rect 28350 8072 28356 8084
rect 27663 8044 28356 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 32861 8075 32919 8081
rect 32861 8041 32873 8075
rect 32907 8072 32919 8075
rect 32950 8072 32956 8084
rect 32907 8044 32956 8072
rect 32907 8041 32919 8044
rect 32861 8035 32919 8041
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 34882 8072 34888 8084
rect 34843 8044 34888 8072
rect 34882 8032 34888 8044
rect 34940 8032 34946 8084
rect 36354 8072 36360 8084
rect 36315 8044 36360 8072
rect 36354 8032 36360 8044
rect 36412 8032 36418 8084
rect 36814 8072 36820 8084
rect 36775 8044 36820 8072
rect 36814 8032 36820 8044
rect 36872 8032 36878 8084
rect 38746 8072 38752 8084
rect 38707 8044 38752 8072
rect 38746 8032 38752 8044
rect 38804 8032 38810 8084
rect 44266 8072 44272 8084
rect 44227 8044 44272 8072
rect 44266 8032 44272 8044
rect 44324 8032 44330 8084
rect 46290 8032 46296 8084
rect 46348 8072 46354 8084
rect 46523 8075 46581 8081
rect 46523 8072 46535 8075
rect 46348 8044 46535 8072
rect 46348 8032 46354 8044
rect 46523 8041 46535 8044
rect 46569 8041 46581 8075
rect 46523 8035 46581 8041
rect 21082 8004 21088 8016
rect 21043 7976 21088 8004
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 22922 7964 22928 8016
rect 22980 8004 22986 8016
rect 24946 8004 24952 8016
rect 22980 7976 24952 8004
rect 22980 7964 22986 7976
rect 24946 7964 24952 7976
rect 25004 7964 25010 8016
rect 25038 7964 25044 8016
rect 25096 8004 25102 8016
rect 25593 8007 25651 8013
rect 25096 7976 25141 8004
rect 25096 7964 25102 7976
rect 25593 7973 25605 8007
rect 25639 8004 25651 8007
rect 26602 8004 26608 8016
rect 25639 7976 26608 8004
rect 25639 7973 25651 7976
rect 25593 7967 25651 7973
rect 26602 7964 26608 7976
rect 26660 7964 26666 8016
rect 26697 8007 26755 8013
rect 26697 7973 26709 8007
rect 26743 8004 26755 8007
rect 26786 8004 26792 8016
rect 26743 7976 26792 8004
rect 26743 7973 26755 7976
rect 26697 7967 26755 7973
rect 26786 7964 26792 7976
rect 26844 7964 26850 8016
rect 28166 7964 28172 8016
rect 28224 8004 28230 8016
rect 28261 8007 28319 8013
rect 28261 8004 28273 8007
rect 28224 7976 28273 8004
rect 28224 7964 28230 7976
rect 28261 7973 28273 7976
rect 28307 7973 28319 8007
rect 28261 7967 28319 7973
rect 30003 8007 30061 8013
rect 30003 7973 30015 8007
rect 30049 8004 30061 8007
rect 30282 8004 30288 8016
rect 30049 7976 30288 8004
rect 30049 7973 30061 7976
rect 30003 7967 30061 7973
rect 30282 7964 30288 7976
rect 30340 7964 30346 8016
rect 33683 8007 33741 8013
rect 33683 7973 33695 8007
rect 33729 8004 33741 8007
rect 33778 8004 33784 8016
rect 33729 7976 33784 8004
rect 33729 7973 33741 7976
rect 33683 7967 33741 7973
rect 33778 7964 33784 7976
rect 33836 7964 33842 8016
rect 35431 8007 35489 8013
rect 35431 7973 35443 8007
rect 35477 8004 35489 8007
rect 35710 8004 35716 8016
rect 35477 7976 35716 8004
rect 35477 7973 35489 7976
rect 35431 7967 35489 7973
rect 35710 7964 35716 7976
rect 35768 7964 35774 8016
rect 39755 8007 39813 8013
rect 39755 7973 39767 8007
rect 39801 8004 39813 8007
rect 39850 8004 39856 8016
rect 39801 7976 39856 8004
rect 39801 7973 39813 7976
rect 39755 7967 39813 7973
rect 39850 7964 39856 7976
rect 39908 7964 39914 8016
rect 45002 8004 45008 8016
rect 44963 7976 45008 8004
rect 45002 7964 45008 7976
rect 45060 7964 45066 8016
rect 45557 8007 45615 8013
rect 45557 7973 45569 8007
rect 45603 8004 45615 8007
rect 45738 8004 45744 8016
rect 45603 7976 45744 8004
rect 45603 7973 45615 7976
rect 45557 7967 45615 7973
rect 45738 7964 45744 7976
rect 45796 7964 45802 8016
rect 46198 8004 46204 8016
rect 46159 7976 46204 8004
rect 46198 7964 46204 7976
rect 46256 7964 46262 8016
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 19426 7936 19432 7948
rect 19484 7945 19490 7948
rect 19484 7939 19522 7945
rect 18932 7908 19432 7936
rect 18932 7896 18938 7908
rect 19426 7896 19432 7908
rect 19510 7905 19522 7939
rect 19484 7899 19522 7905
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 23934 7936 23940 7948
rect 23891 7908 23940 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 19484 7896 19490 7899
rect 23934 7896 23940 7908
rect 23992 7896 23998 7948
rect 29638 7936 29644 7948
rect 29599 7908 29644 7936
rect 29638 7896 29644 7908
rect 29696 7896 29702 7948
rect 32214 7896 32220 7948
rect 32272 7936 32278 7948
rect 32376 7939 32434 7945
rect 32376 7936 32388 7939
rect 32272 7908 32388 7936
rect 32272 7896 32278 7908
rect 32376 7905 32388 7908
rect 32422 7936 32434 7939
rect 34241 7939 34299 7945
rect 34241 7936 34253 7939
rect 32422 7908 34253 7936
rect 32422 7905 32434 7908
rect 32376 7899 32434 7905
rect 34241 7905 34253 7908
rect 34287 7905 34299 7939
rect 34241 7899 34299 7905
rect 34790 7896 34796 7948
rect 34848 7936 34854 7948
rect 35069 7939 35127 7945
rect 35069 7936 35081 7939
rect 34848 7908 35081 7936
rect 34848 7896 34854 7908
rect 35069 7905 35081 7908
rect 35115 7905 35127 7939
rect 35069 7899 35127 7905
rect 38356 7939 38414 7945
rect 38356 7905 38368 7939
rect 38402 7936 38414 7939
rect 38470 7936 38476 7948
rect 38402 7908 38476 7936
rect 38402 7905 38414 7908
rect 38356 7899 38414 7905
rect 38470 7896 38476 7908
rect 38528 7896 38534 7948
rect 41690 7936 41696 7948
rect 41651 7908 41696 7936
rect 41690 7896 41696 7908
rect 41748 7896 41754 7948
rect 42334 7936 42340 7948
rect 42295 7908 42340 7936
rect 42334 7896 42340 7908
rect 42392 7896 42398 7948
rect 43806 7936 43812 7948
rect 43767 7908 43812 7936
rect 43806 7896 43812 7908
rect 43864 7896 43870 7948
rect 45922 7896 45928 7948
rect 45980 7936 45986 7948
rect 46420 7939 46478 7945
rect 46420 7936 46432 7939
rect 45980 7908 46432 7936
rect 45980 7896 45986 7908
rect 46420 7905 46432 7908
rect 46466 7936 46478 7939
rect 47118 7936 47124 7948
rect 46466 7908 47124 7936
rect 46466 7905 46478 7908
rect 46420 7899 46478 7905
rect 47118 7896 47124 7908
rect 47176 7896 47182 7948
rect 47394 7936 47400 7948
rect 47355 7908 47400 7936
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 22646 7868 22652 7880
rect 21039 7840 22652 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 22646 7828 22652 7840
rect 22704 7868 22710 7880
rect 26605 7871 26663 7877
rect 22704 7840 23474 7868
rect 22704 7828 22710 7840
rect 19150 7800 19156 7812
rect 19063 7772 19156 7800
rect 19150 7760 19156 7772
rect 19208 7800 19214 7812
rect 20714 7800 20720 7812
rect 19208 7772 20576 7800
rect 20627 7772 20720 7800
rect 19208 7760 19214 7772
rect 19567 7735 19625 7741
rect 19567 7701 19579 7735
rect 19613 7732 19625 7735
rect 19794 7732 19800 7744
rect 19613 7704 19800 7732
rect 19613 7701 19625 7704
rect 19567 7695 19625 7701
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 20548 7732 20576 7772
rect 20714 7760 20720 7772
rect 20772 7800 20778 7812
rect 21545 7803 21603 7809
rect 21545 7800 21557 7803
rect 20772 7772 21557 7800
rect 20772 7760 20778 7772
rect 21545 7769 21557 7772
rect 21591 7800 21603 7803
rect 21634 7800 21640 7812
rect 21591 7772 21640 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 21634 7760 21640 7772
rect 21692 7760 21698 7812
rect 23446 7800 23474 7840
rect 25424 7840 26464 7868
rect 25424 7800 25452 7840
rect 23446 7772 25452 7800
rect 26436 7800 26464 7840
rect 26605 7837 26617 7871
rect 26651 7868 26663 7871
rect 26694 7868 26700 7880
rect 26651 7840 26700 7868
rect 26651 7837 26663 7840
rect 26605 7831 26663 7837
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 26881 7871 26939 7877
rect 26881 7837 26893 7871
rect 26927 7837 26939 7871
rect 26881 7831 26939 7837
rect 28169 7871 28227 7877
rect 28169 7837 28181 7871
rect 28215 7868 28227 7871
rect 28258 7868 28264 7880
rect 28215 7840 28264 7868
rect 28215 7837 28227 7840
rect 28169 7831 28227 7837
rect 26896 7800 26924 7831
rect 28258 7828 28264 7840
rect 28316 7828 28322 7880
rect 28445 7871 28503 7877
rect 28445 7837 28457 7871
rect 28491 7837 28503 7871
rect 33318 7868 33324 7880
rect 33279 7840 33324 7868
rect 28445 7831 28503 7837
rect 28460 7800 28488 7831
rect 33318 7828 33324 7840
rect 33376 7828 33382 7880
rect 34609 7871 34667 7877
rect 34609 7837 34621 7871
rect 34655 7868 34667 7871
rect 35526 7868 35532 7880
rect 34655 7840 35532 7868
rect 34655 7837 34667 7840
rect 34609 7831 34667 7837
rect 35526 7828 35532 7840
rect 35584 7828 35590 7880
rect 36722 7828 36728 7880
rect 36780 7868 36786 7880
rect 39114 7868 39120 7880
rect 36780 7840 39120 7868
rect 36780 7828 36786 7840
rect 39114 7828 39120 7840
rect 39172 7868 39178 7880
rect 39393 7871 39451 7877
rect 39393 7868 39405 7871
rect 39172 7840 39405 7868
rect 39172 7828 39178 7840
rect 39393 7837 39405 7840
rect 39439 7837 39451 7871
rect 41506 7868 41512 7880
rect 41419 7840 41512 7868
rect 39393 7831 39451 7837
rect 41506 7828 41512 7840
rect 41564 7868 41570 7880
rect 42610 7868 42616 7880
rect 41564 7840 42616 7868
rect 41564 7828 41570 7840
rect 42610 7828 42616 7840
rect 42668 7828 42674 7880
rect 44450 7828 44456 7880
rect 44508 7868 44514 7880
rect 44913 7871 44971 7877
rect 44913 7868 44925 7871
rect 44508 7840 44925 7868
rect 44508 7828 44514 7840
rect 44913 7837 44925 7840
rect 44959 7837 44971 7871
rect 44913 7831 44971 7837
rect 47486 7828 47492 7880
rect 47544 7868 47550 7880
rect 47544 7828 47578 7868
rect 26436 7772 28488 7800
rect 32447 7803 32505 7809
rect 32447 7769 32459 7803
rect 32493 7800 32505 7803
rect 35434 7800 35440 7812
rect 32493 7772 35440 7800
rect 32493 7769 32505 7772
rect 32447 7763 32505 7769
rect 35434 7760 35440 7772
rect 35492 7760 35498 7812
rect 38427 7803 38485 7809
rect 38427 7769 38439 7803
rect 38473 7800 38485 7803
rect 40218 7800 40224 7812
rect 38473 7772 40224 7800
rect 38473 7769 38485 7772
rect 38427 7763 38485 7769
rect 40218 7760 40224 7772
rect 40276 7760 40282 7812
rect 40313 7803 40371 7809
rect 40313 7769 40325 7803
rect 40359 7800 40371 7803
rect 43898 7800 43904 7812
rect 40359 7772 43904 7800
rect 40359 7769 40371 7772
rect 40313 7763 40371 7769
rect 43898 7760 43904 7772
rect 43956 7760 43962 7812
rect 43993 7803 44051 7809
rect 43993 7769 44005 7803
rect 44039 7800 44051 7803
rect 46198 7800 46204 7812
rect 44039 7772 46204 7800
rect 44039 7769 44051 7772
rect 43993 7763 44051 7769
rect 46198 7760 46204 7772
rect 46256 7760 46262 7812
rect 21726 7732 21732 7744
rect 20548 7704 21732 7732
rect 21726 7692 21732 7704
rect 21784 7692 21790 7744
rect 26050 7732 26056 7744
rect 26011 7704 26056 7732
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 30561 7735 30619 7741
rect 30561 7701 30573 7735
rect 30607 7732 30619 7735
rect 30650 7732 30656 7744
rect 30607 7704 30656 7732
rect 30607 7701 30619 7704
rect 30561 7695 30619 7701
rect 30650 7692 30656 7704
rect 30708 7692 30714 7744
rect 30834 7732 30840 7744
rect 30795 7704 30840 7732
rect 30834 7692 30840 7704
rect 30892 7692 30898 7744
rect 31294 7732 31300 7744
rect 31255 7704 31300 7732
rect 31294 7692 31300 7704
rect 31352 7692 31358 7744
rect 35986 7732 35992 7744
rect 35947 7704 35992 7732
rect 35986 7692 35992 7704
rect 36044 7692 36050 7744
rect 44450 7692 44456 7744
rect 44508 7732 44514 7744
rect 47550 7741 47578 7828
rect 44637 7735 44695 7741
rect 44637 7732 44649 7735
rect 44508 7704 44649 7732
rect 44508 7692 44514 7704
rect 44637 7701 44649 7704
rect 44683 7701 44695 7735
rect 44637 7695 44695 7701
rect 47535 7735 47593 7741
rect 47535 7701 47547 7735
rect 47581 7701 47593 7735
rect 47535 7695 47593 7701
rect 1104 7642 48852 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 48852 7642
rect 1104 7568 48852 7590
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 22646 7528 22652 7540
rect 22607 7500 22652 7528
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23934 7528 23940 7540
rect 23339 7500 23940 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 23934 7488 23940 7500
rect 23992 7488 23998 7540
rect 24118 7528 24124 7540
rect 24079 7500 24124 7528
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25225 7531 25283 7537
rect 25225 7528 25237 7531
rect 25004 7500 25237 7528
rect 25004 7488 25010 7500
rect 25225 7497 25237 7500
rect 25271 7497 25283 7531
rect 25225 7491 25283 7497
rect 26050 7488 26056 7540
rect 26108 7528 26114 7540
rect 27847 7531 27905 7537
rect 27847 7528 27859 7531
rect 26108 7500 27859 7528
rect 26108 7488 26114 7500
rect 27847 7497 27859 7500
rect 27893 7497 27905 7531
rect 28166 7528 28172 7540
rect 28127 7500 28172 7528
rect 27847 7491 27905 7497
rect 28166 7488 28172 7500
rect 28224 7488 28230 7540
rect 29641 7531 29699 7537
rect 29641 7497 29653 7531
rect 29687 7528 29699 7531
rect 30466 7528 30472 7540
rect 29687 7500 30472 7528
rect 29687 7497 29699 7500
rect 29641 7491 29699 7497
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20487 7364 20729 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 20717 7361 20729 7364
rect 20763 7392 20775 7395
rect 21082 7392 21088 7404
rect 20763 7364 21088 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21407 7364 22416 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 19794 7324 19800 7336
rect 19755 7296 19800 7324
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 21100 7188 21128 7352
rect 21453 7259 21511 7265
rect 21453 7225 21465 7259
rect 21499 7225 21511 7259
rect 21453 7219 21511 7225
rect 21468 7188 21496 7219
rect 21726 7216 21732 7268
rect 21784 7256 21790 7268
rect 22005 7259 22063 7265
rect 22005 7256 22017 7259
rect 21784 7228 22017 7256
rect 21784 7216 21790 7228
rect 22005 7225 22017 7228
rect 22051 7225 22063 7259
rect 22005 7219 22063 7225
rect 22388 7197 22416 7364
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 24949 7395 25007 7401
rect 24949 7392 24961 7395
rect 24452 7364 24961 7392
rect 24452 7352 24458 7364
rect 24949 7361 24961 7364
rect 24995 7392 25007 7395
rect 25038 7392 25044 7404
rect 24995 7364 25044 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 24118 7284 24124 7336
rect 24176 7324 24182 7336
rect 24305 7327 24363 7333
rect 24305 7324 24317 7327
rect 24176 7296 24317 7324
rect 24176 7284 24182 7296
rect 24305 7293 24317 7296
rect 24351 7293 24363 7327
rect 26237 7327 26295 7333
rect 26237 7324 26249 7327
rect 24305 7287 24363 7293
rect 25976 7296 26249 7324
rect 25976 7200 26004 7296
rect 26237 7293 26249 7296
rect 26283 7293 26295 7327
rect 26237 7287 26295 7293
rect 27614 7284 27620 7336
rect 27672 7324 27678 7336
rect 29783 7333 29811 7500
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 32214 7528 32220 7540
rect 32175 7500 32220 7528
rect 32214 7488 32220 7500
rect 32272 7488 32278 7540
rect 32582 7528 32588 7540
rect 32543 7500 32588 7528
rect 32582 7488 32588 7500
rect 32640 7488 32646 7540
rect 33778 7528 33784 7540
rect 33691 7500 33784 7528
rect 33778 7488 33784 7500
rect 33836 7528 33842 7540
rect 35161 7531 35219 7537
rect 35161 7528 35173 7531
rect 33836 7500 35173 7528
rect 33836 7488 33842 7500
rect 35161 7497 35173 7500
rect 35207 7528 35219 7531
rect 35710 7528 35716 7540
rect 35207 7500 35716 7528
rect 35207 7497 35219 7500
rect 35161 7491 35219 7497
rect 35710 7488 35716 7500
rect 35768 7488 35774 7540
rect 36998 7528 37004 7540
rect 36959 7500 37004 7528
rect 36998 7488 37004 7500
rect 37056 7488 37062 7540
rect 38470 7528 38476 7540
rect 38431 7500 38476 7528
rect 38470 7488 38476 7500
rect 38528 7528 38534 7540
rect 38749 7531 38807 7537
rect 38749 7528 38761 7531
rect 38528 7500 38761 7528
rect 38528 7488 38534 7500
rect 38749 7497 38761 7500
rect 38795 7497 38807 7531
rect 39114 7528 39120 7540
rect 39075 7500 39120 7528
rect 38749 7491 38807 7497
rect 39114 7488 39120 7500
rect 39172 7488 39178 7540
rect 42334 7488 42340 7540
rect 42392 7528 42398 7540
rect 42521 7531 42579 7537
rect 42521 7528 42533 7531
rect 42392 7500 42533 7528
rect 42392 7488 42398 7500
rect 42521 7497 42533 7500
rect 42567 7497 42579 7531
rect 42521 7491 42579 7497
rect 42610 7488 42616 7540
rect 42668 7528 42674 7540
rect 43211 7531 43269 7537
rect 43211 7528 43223 7531
rect 42668 7500 43223 7528
rect 42668 7488 42674 7500
rect 43211 7497 43223 7500
rect 43257 7497 43269 7531
rect 43806 7528 43812 7540
rect 43767 7500 43812 7528
rect 43211 7491 43269 7497
rect 43806 7488 43812 7500
rect 43864 7488 43870 7540
rect 44358 7528 44364 7540
rect 44319 7500 44364 7528
rect 44358 7488 44364 7500
rect 44416 7488 44422 7540
rect 45002 7488 45008 7540
rect 45060 7528 45066 7540
rect 45557 7531 45615 7537
rect 45557 7528 45569 7531
rect 45060 7500 45569 7528
rect 45060 7488 45066 7500
rect 45557 7497 45569 7500
rect 45603 7528 45615 7531
rect 45925 7531 45983 7537
rect 45925 7528 45937 7531
rect 45603 7500 45937 7528
rect 45603 7497 45615 7500
rect 45557 7491 45615 7497
rect 45925 7497 45937 7500
rect 45971 7528 45983 7531
rect 46106 7528 46112 7540
rect 45971 7500 46112 7528
rect 45971 7497 45983 7500
rect 45925 7491 45983 7497
rect 46106 7488 46112 7500
rect 46164 7488 46170 7540
rect 47118 7528 47124 7540
rect 47079 7500 47124 7528
rect 47118 7488 47124 7500
rect 47176 7488 47182 7540
rect 30282 7460 30288 7472
rect 30195 7432 30288 7460
rect 30282 7420 30288 7432
rect 30340 7460 30346 7472
rect 33796 7460 33824 7488
rect 30340 7432 33824 7460
rect 30340 7420 30346 7432
rect 29871 7395 29929 7401
rect 29871 7361 29883 7395
rect 29917 7392 29929 7395
rect 30834 7392 30840 7404
rect 29917 7364 30840 7392
rect 29917 7361 29929 7364
rect 29871 7355 29929 7361
rect 30834 7352 30840 7364
rect 30892 7352 30898 7404
rect 31478 7392 31484 7404
rect 31439 7364 31484 7392
rect 31478 7352 31484 7364
rect 31536 7352 31542 7404
rect 33318 7352 33324 7404
rect 33376 7392 33382 7404
rect 33413 7395 33471 7401
rect 33413 7392 33425 7395
rect 33376 7364 33425 7392
rect 33376 7352 33382 7364
rect 33413 7361 33425 7364
rect 33459 7392 33471 7395
rect 34057 7395 34115 7401
rect 34057 7392 34069 7395
rect 33459 7364 34069 7392
rect 33459 7361 33471 7364
rect 33413 7355 33471 7361
rect 34057 7361 34069 7364
rect 34103 7361 34115 7395
rect 35618 7392 35624 7404
rect 35531 7364 35624 7392
rect 34057 7355 34115 7361
rect 35618 7352 35624 7364
rect 35676 7392 35682 7404
rect 36541 7395 36599 7401
rect 36541 7392 36553 7395
rect 35676 7364 36553 7392
rect 35676 7352 35682 7364
rect 36541 7361 36553 7364
rect 36587 7361 36599 7395
rect 37016 7392 37044 7488
rect 39574 7420 39580 7472
rect 39632 7460 39638 7472
rect 42889 7463 42947 7469
rect 42889 7460 42901 7463
rect 39632 7432 42901 7460
rect 39632 7420 39638 7432
rect 42889 7429 42901 7432
rect 42935 7429 42947 7463
rect 42889 7423 42947 7429
rect 37553 7395 37611 7401
rect 37553 7392 37565 7395
rect 37016 7364 37565 7392
rect 36541 7355 36599 7361
rect 37553 7361 37565 7364
rect 37599 7361 37611 7395
rect 37553 7355 37611 7361
rect 40678 7352 40684 7404
rect 40736 7392 40742 7404
rect 41509 7395 41567 7401
rect 41509 7392 41521 7395
rect 40736 7364 41521 7392
rect 40736 7352 40742 7364
rect 41509 7361 41521 7364
rect 41555 7361 41567 7395
rect 41509 7355 41567 7361
rect 27744 7327 27802 7333
rect 27744 7324 27756 7327
rect 27672 7296 27756 7324
rect 27672 7284 27678 7296
rect 27744 7293 27756 7296
rect 27790 7324 27802 7327
rect 28537 7327 28595 7333
rect 28537 7324 28549 7327
rect 27790 7296 28549 7324
rect 27790 7293 27802 7296
rect 27744 7287 27802 7293
rect 28537 7293 28549 7296
rect 28583 7293 28595 7327
rect 28537 7287 28595 7293
rect 29768 7327 29826 7333
rect 29768 7293 29780 7327
rect 29814 7293 29826 7327
rect 29768 7287 29826 7293
rect 32582 7284 32588 7336
rect 32640 7324 32646 7336
rect 32677 7327 32735 7333
rect 32677 7324 32689 7327
rect 32640 7296 32689 7324
rect 32640 7284 32646 7296
rect 32677 7293 32689 7296
rect 32723 7293 32735 7327
rect 32677 7287 32735 7293
rect 32766 7284 32772 7336
rect 32824 7324 32830 7336
rect 33137 7327 33195 7333
rect 33137 7324 33149 7327
rect 32824 7296 33149 7324
rect 32824 7284 32830 7296
rect 33137 7293 33149 7296
rect 33183 7293 33195 7327
rect 33137 7287 33195 7293
rect 38654 7284 38660 7336
rect 38712 7324 38718 7336
rect 39336 7327 39394 7333
rect 39336 7324 39348 7327
rect 38712 7296 39348 7324
rect 38712 7284 38718 7296
rect 39336 7293 39348 7296
rect 39382 7324 39394 7327
rect 40129 7327 40187 7333
rect 40129 7324 40141 7327
rect 39382 7296 40141 7324
rect 39382 7293 39394 7296
rect 39336 7287 39394 7293
rect 40129 7293 40141 7296
rect 40175 7293 40187 7327
rect 40129 7287 40187 7293
rect 40564 7327 40622 7333
rect 40564 7293 40576 7327
rect 40610 7324 40622 7327
rect 41417 7327 41475 7333
rect 40610 7296 41092 7324
rect 40610 7293 40622 7296
rect 40564 7287 40622 7293
rect 28258 7216 28264 7268
rect 28316 7256 28322 7268
rect 28997 7259 29055 7265
rect 28997 7256 29009 7259
rect 28316 7228 29009 7256
rect 28316 7216 28322 7228
rect 28997 7225 29009 7228
rect 29043 7256 29055 7259
rect 30926 7256 30932 7268
rect 29043 7228 30696 7256
rect 30887 7228 30932 7256
rect 29043 7225 29055 7228
rect 28997 7219 29055 7225
rect 21100 7160 21496 7188
rect 22373 7191 22431 7197
rect 22373 7157 22385 7191
rect 22419 7188 22431 7191
rect 22462 7188 22468 7200
rect 22419 7160 22468 7188
rect 22419 7157 22431 7160
rect 22373 7151 22431 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24578 7188 24584 7200
rect 24535 7160 24584 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24578 7148 24584 7160
rect 24636 7148 24642 7200
rect 25958 7188 25964 7200
rect 25919 7160 25964 7188
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 26418 7188 26424 7200
rect 26379 7160 26424 7188
rect 26418 7148 26424 7160
rect 26476 7188 26482 7200
rect 26786 7188 26792 7200
rect 26476 7160 26792 7188
rect 26476 7148 26482 7160
rect 26786 7148 26792 7160
rect 26844 7188 26850 7200
rect 27157 7191 27215 7197
rect 27157 7188 27169 7191
rect 26844 7160 27169 7188
rect 26844 7148 26850 7160
rect 27157 7157 27169 7160
rect 27203 7157 27215 7191
rect 30558 7188 30564 7200
rect 30519 7160 30564 7188
rect 27157 7151 27215 7157
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 30668 7188 30696 7228
rect 30926 7216 30932 7228
rect 30984 7216 30990 7268
rect 34701 7259 34759 7265
rect 34701 7225 34713 7259
rect 34747 7256 34759 7259
rect 35710 7256 35716 7268
rect 34747 7228 35716 7256
rect 34747 7225 34759 7228
rect 34701 7219 34759 7225
rect 35710 7216 35716 7228
rect 35768 7216 35774 7268
rect 36262 7256 36268 7268
rect 36223 7228 36268 7256
rect 36262 7216 36268 7228
rect 36320 7216 36326 7268
rect 37461 7259 37519 7265
rect 37461 7225 37473 7259
rect 37507 7256 37519 7259
rect 37915 7259 37973 7265
rect 37915 7256 37927 7259
rect 37507 7228 37927 7256
rect 37507 7225 37519 7228
rect 37461 7219 37519 7225
rect 37915 7225 37927 7228
rect 37961 7256 37973 7259
rect 38010 7256 38016 7268
rect 37961 7228 38016 7256
rect 37961 7225 37973 7228
rect 37915 7219 37973 7225
rect 38010 7216 38016 7228
rect 38068 7216 38074 7268
rect 39022 7216 39028 7268
rect 39080 7256 39086 7268
rect 39439 7259 39497 7265
rect 39439 7256 39451 7259
rect 39080 7228 39451 7256
rect 39080 7216 39086 7228
rect 39439 7225 39451 7228
rect 39485 7225 39497 7259
rect 39439 7219 39497 7225
rect 31478 7188 31484 7200
rect 30668 7160 31484 7188
rect 31478 7148 31484 7160
rect 31536 7148 31542 7200
rect 39761 7191 39819 7197
rect 39761 7157 39773 7191
rect 39807 7188 39819 7191
rect 39850 7188 39856 7200
rect 39807 7160 39856 7188
rect 39807 7157 39819 7160
rect 39761 7151 39819 7157
rect 39850 7148 39856 7160
rect 39908 7148 39914 7200
rect 40635 7191 40693 7197
rect 40635 7157 40647 7191
rect 40681 7188 40693 7191
rect 40862 7188 40868 7200
rect 40681 7160 40868 7188
rect 40681 7157 40693 7160
rect 40635 7151 40693 7157
rect 40862 7148 40868 7160
rect 40920 7148 40926 7200
rect 41064 7197 41092 7296
rect 41417 7293 41429 7327
rect 41463 7324 41475 7327
rect 42150 7324 42156 7336
rect 41463 7296 42156 7324
rect 41463 7293 41475 7296
rect 41417 7287 41475 7293
rect 42150 7284 42156 7296
rect 42208 7284 42214 7336
rect 42904 7324 42932 7423
rect 43898 7420 43904 7472
rect 43956 7460 43962 7472
rect 47394 7460 47400 7472
rect 43956 7432 47400 7460
rect 43956 7420 43962 7432
rect 47394 7420 47400 7432
rect 47452 7460 47458 7472
rect 47489 7463 47547 7469
rect 47489 7460 47501 7463
rect 47452 7432 47501 7460
rect 47452 7420 47458 7432
rect 47489 7429 47501 7432
rect 47535 7429 47547 7463
rect 47489 7423 47547 7429
rect 45189 7395 45247 7401
rect 45189 7361 45201 7395
rect 45235 7392 45247 7395
rect 45738 7392 45744 7404
rect 45235 7364 45744 7392
rect 45235 7361 45247 7364
rect 45189 7355 45247 7361
rect 45738 7352 45744 7364
rect 45796 7352 45802 7404
rect 46382 7352 46388 7404
rect 46440 7392 46446 7404
rect 46477 7395 46535 7401
rect 46477 7392 46489 7395
rect 46440 7364 46489 7392
rect 46440 7352 46446 7364
rect 46477 7361 46489 7364
rect 46523 7361 46535 7395
rect 46477 7355 46535 7361
rect 43108 7327 43166 7333
rect 43108 7324 43120 7327
rect 42904 7296 43120 7324
rect 43108 7293 43120 7296
rect 43154 7293 43166 7327
rect 43108 7287 43166 7293
rect 44542 7256 44548 7268
rect 44503 7228 44548 7256
rect 44542 7216 44548 7228
rect 44600 7216 44606 7268
rect 44637 7259 44695 7265
rect 44637 7225 44649 7259
rect 44683 7225 44695 7259
rect 46198 7256 46204 7268
rect 46159 7228 46204 7256
rect 44637 7219 44695 7225
rect 41049 7191 41107 7197
rect 41049 7157 41061 7191
rect 41095 7188 41107 7191
rect 41138 7188 41144 7200
rect 41095 7160 41144 7188
rect 41095 7157 41107 7160
rect 41049 7151 41107 7157
rect 41138 7148 41144 7160
rect 41196 7148 41202 7200
rect 44358 7148 44364 7200
rect 44416 7188 44422 7200
rect 44652 7188 44680 7219
rect 46198 7216 46204 7228
rect 46256 7216 46262 7268
rect 46293 7259 46351 7265
rect 46293 7225 46305 7259
rect 46339 7225 46351 7259
rect 46293 7219 46351 7225
rect 44416 7160 44680 7188
rect 44416 7148 44422 7160
rect 46106 7148 46112 7200
rect 46164 7188 46170 7200
rect 46308 7188 46336 7219
rect 46164 7160 46336 7188
rect 46164 7148 46170 7160
rect 1104 7098 48852 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 48852 7098
rect 1104 7024 48852 7046
rect 26694 6984 26700 6996
rect 26655 6956 26700 6984
rect 26694 6944 26700 6956
rect 26752 6944 26758 6996
rect 29638 6944 29644 6996
rect 29696 6984 29702 6996
rect 29825 6987 29883 6993
rect 29825 6984 29837 6987
rect 29696 6956 29837 6984
rect 29696 6944 29702 6956
rect 29825 6953 29837 6956
rect 29871 6953 29883 6987
rect 32677 6987 32735 6993
rect 32677 6984 32689 6987
rect 29825 6947 29883 6953
rect 30018 6956 32689 6984
rect 19797 6919 19855 6925
rect 19797 6885 19809 6919
rect 19843 6916 19855 6919
rect 19886 6916 19892 6928
rect 19843 6888 19892 6916
rect 19843 6885 19855 6888
rect 19797 6879 19855 6885
rect 19886 6876 19892 6888
rect 19944 6876 19950 6928
rect 21082 6916 21088 6928
rect 21043 6888 21088 6916
rect 21082 6876 21088 6888
rect 21140 6876 21146 6928
rect 21634 6916 21640 6928
rect 21595 6888 21640 6916
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 22827 6919 22885 6925
rect 22827 6885 22839 6919
rect 22873 6916 22885 6919
rect 23106 6916 23112 6928
rect 22873 6888 23112 6916
rect 22873 6885 22885 6888
rect 22827 6879 22885 6885
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 27433 6919 27491 6925
rect 27433 6885 27445 6919
rect 27479 6916 27491 6919
rect 28166 6916 28172 6928
rect 27479 6888 28172 6916
rect 27479 6885 27491 6888
rect 27433 6879 27491 6885
rect 28166 6876 28172 6888
rect 28224 6876 28230 6928
rect 28994 6876 29000 6928
rect 29052 6916 29058 6928
rect 29052 6888 29097 6916
rect 29052 6876 29058 6888
rect 29178 6876 29184 6928
rect 29236 6916 29242 6928
rect 30018 6916 30046 6956
rect 32677 6953 32689 6956
rect 32723 6984 32735 6987
rect 32766 6984 32772 6996
rect 32723 6956 32772 6984
rect 32723 6953 32735 6956
rect 32677 6947 32735 6953
rect 32766 6944 32772 6956
rect 32824 6944 32830 6996
rect 35069 6987 35127 6993
rect 35069 6953 35081 6987
rect 35115 6984 35127 6987
rect 35250 6984 35256 6996
rect 35115 6956 35256 6984
rect 35115 6953 35127 6956
rect 35069 6947 35127 6953
rect 35250 6944 35256 6956
rect 35308 6984 35314 6996
rect 35986 6984 35992 6996
rect 35308 6956 35992 6984
rect 35308 6944 35314 6956
rect 35986 6944 35992 6956
rect 36044 6944 36050 6996
rect 42150 6944 42156 6996
rect 42208 6984 42214 6996
rect 42245 6987 42303 6993
rect 42245 6984 42257 6987
rect 42208 6956 42257 6984
rect 42208 6944 42214 6956
rect 42245 6953 42257 6956
rect 42291 6953 42303 6987
rect 42245 6947 42303 6953
rect 42334 6944 42340 6996
rect 42392 6984 42398 6996
rect 46615 6987 46673 6993
rect 46615 6984 46627 6987
rect 42392 6956 46627 6984
rect 42392 6944 42398 6956
rect 46615 6953 46627 6956
rect 46661 6953 46673 6987
rect 46615 6947 46673 6953
rect 29236 6888 30046 6916
rect 29236 6876 29242 6888
rect 30098 6876 30104 6928
rect 30156 6916 30162 6928
rect 30558 6916 30564 6928
rect 30156 6888 30564 6916
rect 30156 6876 30162 6888
rect 30558 6876 30564 6888
rect 30616 6916 30622 6928
rect 30653 6919 30711 6925
rect 30653 6916 30665 6919
rect 30616 6888 30665 6916
rect 30616 6876 30622 6888
rect 30653 6885 30665 6888
rect 30699 6916 30711 6919
rect 30926 6916 30932 6928
rect 30699 6888 30932 6916
rect 30699 6885 30711 6888
rect 30653 6879 30711 6885
rect 30926 6876 30932 6888
rect 30984 6876 30990 6928
rect 34790 6876 34796 6928
rect 34848 6916 34854 6928
rect 35345 6919 35403 6925
rect 35345 6916 35357 6919
rect 34848 6888 35357 6916
rect 34848 6876 34854 6888
rect 35345 6885 35357 6888
rect 35391 6885 35403 6919
rect 35345 6879 35403 6885
rect 35434 6876 35440 6928
rect 35492 6916 35498 6928
rect 35621 6919 35679 6925
rect 35621 6916 35633 6919
rect 35492 6888 35633 6916
rect 35492 6876 35498 6888
rect 35621 6885 35633 6888
rect 35667 6885 35679 6919
rect 35621 6879 35679 6885
rect 35713 6919 35771 6925
rect 35713 6885 35725 6919
rect 35759 6916 35771 6919
rect 35802 6916 35808 6928
rect 35759 6888 35808 6916
rect 35759 6885 35771 6888
rect 35713 6879 35771 6885
rect 35802 6876 35808 6888
rect 35860 6876 35866 6928
rect 39022 6916 39028 6928
rect 38983 6888 39028 6916
rect 39022 6876 39028 6888
rect 39080 6876 39086 6928
rect 39114 6876 39120 6928
rect 39172 6916 39178 6928
rect 39172 6888 39217 6916
rect 39172 6876 39178 6888
rect 40218 6876 40224 6928
rect 40276 6916 40282 6928
rect 40589 6919 40647 6925
rect 40589 6916 40601 6919
rect 40276 6888 40601 6916
rect 40276 6876 40282 6888
rect 40589 6885 40601 6888
rect 40635 6885 40647 6919
rect 40589 6879 40647 6885
rect 40678 6876 40684 6928
rect 40736 6916 40742 6928
rect 43530 6916 43536 6928
rect 40736 6888 40781 6916
rect 43491 6888 43536 6916
rect 40736 6876 40742 6888
rect 43530 6876 43536 6888
rect 43588 6876 43594 6928
rect 44358 6876 44364 6928
rect 44416 6916 44422 6928
rect 45097 6919 45155 6925
rect 45097 6916 45109 6919
rect 44416 6888 45109 6916
rect 44416 6876 44422 6888
rect 45097 6885 45109 6888
rect 45143 6916 45155 6919
rect 45186 6916 45192 6928
rect 45143 6888 45192 6916
rect 45143 6885 45155 6888
rect 45097 6879 45155 6885
rect 45186 6876 45192 6888
rect 45244 6876 45250 6928
rect 45649 6919 45707 6925
rect 45649 6885 45661 6919
rect 45695 6916 45707 6919
rect 46382 6916 46388 6928
rect 45695 6888 46388 6916
rect 45695 6885 45707 6888
rect 45649 6879 45707 6885
rect 46382 6876 46388 6888
rect 46440 6876 46446 6928
rect 19153 6851 19211 6857
rect 19153 6817 19165 6851
rect 19199 6848 19211 6851
rect 19426 6848 19432 6860
rect 19199 6820 19432 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 24280 6851 24338 6857
rect 24280 6817 24292 6851
rect 24326 6848 24338 6851
rect 24670 6848 24676 6860
rect 24326 6820 24676 6848
rect 24326 6817 24338 6820
rect 24280 6811 24338 6817
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 32582 6808 32588 6860
rect 32640 6848 32646 6860
rect 32950 6848 32956 6860
rect 32640 6820 32956 6848
rect 32640 6808 32646 6820
rect 32950 6808 32956 6820
rect 33008 6808 33014 6860
rect 33410 6808 33416 6860
rect 33468 6848 33474 6860
rect 33965 6851 34023 6857
rect 33965 6848 33977 6851
rect 33468 6820 33977 6848
rect 33468 6808 33474 6820
rect 33965 6817 33977 6820
rect 34011 6817 34023 6851
rect 33965 6811 34023 6817
rect 34517 6851 34575 6857
rect 34517 6817 34529 6851
rect 34563 6848 34575 6851
rect 34606 6848 34612 6860
rect 34563 6820 34612 6848
rect 34563 6817 34575 6820
rect 34517 6811 34575 6817
rect 34606 6808 34612 6820
rect 34664 6848 34670 6860
rect 35158 6848 35164 6860
rect 34664 6820 35164 6848
rect 34664 6808 34670 6820
rect 35158 6808 35164 6820
rect 35216 6808 35222 6860
rect 37734 6848 37740 6860
rect 37695 6820 37740 6848
rect 37734 6808 37740 6820
rect 37792 6808 37798 6860
rect 42061 6851 42119 6857
rect 42061 6817 42073 6851
rect 42107 6848 42119 6851
rect 42150 6848 42156 6860
rect 42107 6820 42156 6848
rect 42107 6817 42119 6820
rect 42061 6811 42119 6817
rect 42150 6808 42156 6820
rect 42208 6848 42214 6860
rect 42702 6848 42708 6860
rect 42208 6820 42708 6848
rect 42208 6808 42214 6820
rect 42702 6808 42708 6820
rect 42760 6808 42766 6860
rect 46198 6848 46204 6860
rect 46159 6820 46204 6848
rect 46198 6808 46204 6820
rect 46256 6808 46262 6860
rect 46290 6808 46296 6860
rect 46348 6848 46354 6860
rect 46512 6851 46570 6857
rect 46512 6848 46524 6851
rect 46348 6820 46524 6848
rect 46348 6808 46354 6820
rect 46512 6817 46524 6820
rect 46558 6817 46570 6851
rect 46512 6811 46570 6817
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21358 6780 21364 6792
rect 21039 6752 21364 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22388 6752 22477 6780
rect 22388 6656 22416 6752
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6780 27399 6783
rect 27982 6780 27988 6792
rect 27387 6752 27988 6780
rect 27387 6749 27399 6752
rect 27341 6743 27399 6749
rect 27982 6740 27988 6752
rect 28040 6740 28046 6792
rect 28905 6783 28963 6789
rect 28905 6780 28917 6783
rect 28736 6752 28917 6780
rect 27246 6672 27252 6724
rect 27304 6712 27310 6724
rect 27893 6715 27951 6721
rect 27893 6712 27905 6715
rect 27304 6684 27905 6712
rect 27304 6672 27310 6684
rect 27893 6681 27905 6684
rect 27939 6681 27951 6715
rect 27893 6675 27951 6681
rect 19334 6644 19340 6656
rect 19295 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 22370 6644 22376 6656
rect 22331 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 23382 6644 23388 6656
rect 23343 6616 23388 6644
rect 23382 6604 23388 6616
rect 23440 6604 23446 6656
rect 23750 6644 23756 6656
rect 23663 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6644 23814 6656
rect 24351 6647 24409 6653
rect 24351 6644 24363 6647
rect 23808 6616 24363 6644
rect 23808 6604 23814 6616
rect 24351 6613 24363 6616
rect 24397 6613 24409 6647
rect 25314 6644 25320 6656
rect 25275 6616 25320 6644
rect 24351 6607 24409 6613
rect 25314 6604 25320 6616
rect 25372 6604 25378 6656
rect 25590 6644 25596 6656
rect 25551 6616 25596 6644
rect 25590 6604 25596 6616
rect 25648 6604 25654 6656
rect 27154 6644 27160 6656
rect 27115 6616 27160 6644
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 28626 6644 28632 6656
rect 28587 6616 28632 6644
rect 28626 6604 28632 6616
rect 28684 6644 28690 6656
rect 28736 6644 28764 6752
rect 28905 6749 28917 6752
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 30561 6783 30619 6789
rect 30561 6749 30573 6783
rect 30607 6780 30619 6783
rect 31754 6780 31760 6792
rect 30607 6752 31760 6780
rect 30607 6749 30619 6752
rect 30561 6743 30619 6749
rect 31754 6740 31760 6752
rect 31812 6740 31818 6792
rect 34698 6780 34704 6792
rect 34659 6752 34704 6780
rect 34698 6740 34704 6752
rect 34756 6740 34762 6792
rect 36262 6780 36268 6792
rect 36223 6752 36268 6780
rect 36262 6740 36268 6752
rect 36320 6740 36326 6792
rect 40865 6783 40923 6789
rect 40865 6749 40877 6783
rect 40911 6749 40923 6783
rect 43438 6780 43444 6792
rect 43399 6752 43444 6780
rect 40865 6743 40923 6749
rect 28810 6672 28816 6724
rect 28868 6712 28874 6724
rect 29457 6715 29515 6721
rect 29457 6712 29469 6715
rect 28868 6684 29469 6712
rect 28868 6672 28874 6684
rect 29457 6681 29469 6684
rect 29503 6712 29515 6715
rect 31113 6715 31171 6721
rect 31113 6712 31125 6715
rect 29503 6684 31125 6712
rect 29503 6681 29515 6684
rect 29457 6675 29515 6681
rect 31113 6681 31125 6684
rect 31159 6681 31171 6715
rect 31113 6675 31171 6681
rect 39577 6715 39635 6721
rect 39577 6681 39589 6715
rect 39623 6712 39635 6715
rect 40880 6712 40908 6743
rect 43438 6740 43444 6752
rect 43496 6740 43502 6792
rect 43898 6740 43904 6792
rect 43956 6780 43962 6792
rect 44085 6783 44143 6789
rect 44085 6780 44097 6783
rect 43956 6752 44097 6780
rect 43956 6740 43962 6752
rect 44085 6749 44097 6752
rect 44131 6780 44143 6783
rect 45005 6783 45063 6789
rect 45005 6780 45017 6783
rect 44131 6752 45017 6780
rect 44131 6749 44143 6752
rect 44085 6743 44143 6749
rect 45005 6749 45017 6752
rect 45051 6749 45063 6783
rect 45005 6743 45063 6749
rect 42610 6712 42616 6724
rect 39623 6684 42616 6712
rect 39623 6681 39635 6684
rect 39577 6675 39635 6681
rect 42610 6672 42616 6684
rect 42668 6672 42674 6724
rect 28684 6616 28764 6644
rect 33137 6647 33195 6653
rect 28684 6604 28690 6616
rect 33137 6613 33149 6647
rect 33183 6644 33195 6647
rect 33410 6644 33416 6656
rect 33183 6616 33416 6644
rect 33183 6613 33195 6616
rect 33137 6607 33195 6613
rect 33410 6604 33416 6616
rect 33468 6604 33474 6656
rect 36262 6604 36268 6656
rect 36320 6644 36326 6656
rect 36541 6647 36599 6653
rect 36541 6644 36553 6647
rect 36320 6616 36553 6644
rect 36320 6604 36326 6616
rect 36541 6613 36553 6616
rect 36587 6613 36599 6647
rect 36541 6607 36599 6613
rect 37921 6647 37979 6653
rect 37921 6613 37933 6647
rect 37967 6644 37979 6647
rect 38286 6644 38292 6656
rect 37967 6616 38292 6644
rect 37967 6613 37979 6616
rect 37921 6607 37979 6613
rect 38286 6604 38292 6616
rect 38344 6604 38350 6656
rect 38470 6644 38476 6656
rect 38431 6616 38476 6644
rect 38470 6604 38476 6616
rect 38528 6604 38534 6656
rect 41046 6604 41052 6656
rect 41104 6644 41110 6656
rect 41601 6647 41659 6653
rect 41601 6644 41613 6647
rect 41104 6616 41613 6644
rect 41104 6604 41110 6616
rect 41601 6613 41613 6616
rect 41647 6644 41659 6647
rect 42334 6644 42340 6656
rect 41647 6616 42340 6644
rect 41647 6613 41659 6616
rect 41601 6607 41659 6613
rect 42334 6604 42340 6616
rect 42392 6604 42398 6656
rect 44082 6604 44088 6656
rect 44140 6644 44146 6656
rect 44453 6647 44511 6653
rect 44453 6644 44465 6647
rect 44140 6616 44465 6644
rect 44140 6604 44146 6616
rect 44453 6613 44465 6616
rect 44499 6644 44511 6647
rect 44542 6644 44548 6656
rect 44499 6616 44548 6644
rect 44499 6613 44511 6616
rect 44453 6607 44511 6613
rect 44542 6604 44548 6616
rect 44600 6604 44606 6656
rect 1104 6554 48852 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 48852 6554
rect 1104 6480 48852 6502
rect 19245 6443 19303 6449
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19426 6440 19432 6452
rect 19291 6412 19432 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 20346 6440 20352 6452
rect 20211 6412 20352 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 20346 6400 20352 6412
rect 20404 6440 20410 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20404 6412 21005 6440
rect 20404 6400 20410 6412
rect 20993 6409 21005 6412
rect 21039 6440 21051 6443
rect 21082 6440 21088 6452
rect 21039 6412 21088 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 25406 6400 25412 6452
rect 25464 6440 25470 6452
rect 26237 6443 26295 6449
rect 26237 6440 26249 6443
rect 25464 6412 26249 6440
rect 25464 6400 25470 6412
rect 26237 6409 26249 6412
rect 26283 6409 26295 6443
rect 26237 6403 26295 6409
rect 27893 6443 27951 6449
rect 27893 6409 27905 6443
rect 27939 6440 27951 6443
rect 28166 6440 28172 6452
rect 27939 6412 28172 6440
rect 27939 6409 27951 6412
rect 27893 6403 27951 6409
rect 28166 6400 28172 6412
rect 28224 6400 28230 6452
rect 28442 6440 28448 6452
rect 28403 6412 28448 6440
rect 28442 6400 28448 6412
rect 28500 6400 28506 6452
rect 28905 6443 28963 6449
rect 28905 6409 28917 6443
rect 28951 6440 28963 6443
rect 28994 6440 29000 6452
rect 28951 6412 29000 6440
rect 28951 6409 28963 6412
rect 28905 6403 28963 6409
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 30282 6400 30288 6452
rect 30340 6440 30346 6452
rect 30377 6443 30435 6449
rect 30377 6440 30389 6443
rect 30340 6412 30389 6440
rect 30340 6400 30346 6412
rect 30377 6409 30389 6412
rect 30423 6409 30435 6443
rect 31754 6440 31760 6452
rect 31715 6412 31760 6440
rect 30377 6403 30435 6409
rect 31754 6400 31760 6412
rect 31812 6400 31818 6452
rect 32950 6440 32956 6452
rect 32911 6412 32956 6440
rect 32950 6400 32956 6412
rect 33008 6440 33014 6452
rect 34606 6440 34612 6452
rect 33008 6412 33134 6440
rect 34567 6412 34612 6440
rect 33008 6400 33014 6412
rect 22462 6332 22468 6384
rect 22520 6372 22526 6384
rect 27338 6372 27344 6384
rect 22520 6344 27344 6372
rect 22520 6332 22526 6344
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 22557 6307 22615 6313
rect 22557 6304 22569 6307
rect 22428 6276 22569 6304
rect 22428 6264 22434 6276
rect 22557 6273 22569 6276
rect 22603 6273 22615 6307
rect 23750 6304 23756 6316
rect 23711 6276 23756 6304
rect 22557 6267 22615 6273
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6304 24455 6307
rect 24854 6304 24860 6316
rect 24443 6276 24860 6304
rect 24443 6273 24455 6276
rect 24397 6267 24455 6273
rect 24854 6264 24860 6276
rect 24912 6304 24918 6316
rect 25314 6304 25320 6316
rect 24912 6276 25320 6304
rect 24912 6264 24918 6276
rect 25314 6264 25320 6276
rect 25372 6264 25378 6316
rect 25608 6313 25636 6344
rect 27338 6332 27344 6344
rect 27396 6332 27402 6384
rect 27982 6332 27988 6384
rect 28040 6372 28046 6384
rect 28810 6372 28816 6384
rect 28040 6344 28816 6372
rect 28040 6332 28046 6344
rect 28810 6332 28816 6344
rect 28868 6332 28874 6384
rect 33106 6372 33134 6412
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 35023 6443 35081 6449
rect 35023 6409 35035 6443
rect 35069 6440 35081 6443
rect 35618 6440 35624 6452
rect 35069 6412 35624 6440
rect 35069 6409 35081 6412
rect 35023 6403 35081 6409
rect 35618 6400 35624 6412
rect 35676 6400 35682 6452
rect 38286 6440 38292 6452
rect 38247 6412 38292 6440
rect 38286 6400 38292 6412
rect 38344 6400 38350 6452
rect 42150 6440 42156 6452
rect 42111 6412 42156 6440
rect 42150 6400 42156 6412
rect 42208 6400 42214 6452
rect 42610 6440 42616 6452
rect 42571 6412 42616 6440
rect 42610 6400 42616 6412
rect 42668 6440 42674 6452
rect 42668 6412 42794 6440
rect 42668 6400 42674 6412
rect 36078 6372 36084 6384
rect 33106 6344 36084 6372
rect 36078 6332 36084 6344
rect 36136 6372 36142 6384
rect 37734 6372 37740 6384
rect 36136 6344 37740 6372
rect 36136 6332 36142 6344
rect 37734 6332 37740 6344
rect 37792 6332 37798 6384
rect 25593 6307 25651 6313
rect 25593 6273 25605 6307
rect 25639 6273 25651 6307
rect 25593 6267 25651 6273
rect 26881 6307 26939 6313
rect 26881 6273 26893 6307
rect 26927 6304 26939 6307
rect 27154 6304 27160 6316
rect 26927 6276 27160 6304
rect 26927 6273 26939 6276
rect 26881 6267 26939 6273
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27304 6276 27349 6304
rect 27304 6264 27310 6276
rect 30466 6264 30472 6316
rect 30524 6304 30530 6316
rect 32677 6307 32735 6313
rect 32677 6304 32689 6307
rect 30524 6276 32689 6304
rect 30524 6264 30530 6276
rect 32677 6273 32689 6276
rect 32723 6304 32735 6307
rect 33318 6304 33324 6316
rect 32723 6276 33324 6304
rect 32723 6273 32735 6276
rect 32677 6267 32735 6273
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19392 6208 19625 6236
rect 19392 6196 19398 6208
rect 19613 6205 19625 6208
rect 19659 6236 19671 6239
rect 19797 6239 19855 6245
rect 19797 6236 19809 6239
rect 19659 6208 19809 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 19797 6205 19809 6208
rect 19843 6205 19855 6239
rect 19797 6199 19855 6205
rect 21913 6239 21971 6245
rect 21913 6205 21925 6239
rect 21959 6236 21971 6239
rect 22094 6236 22100 6248
rect 21959 6208 22100 6236
rect 21959 6205 21971 6208
rect 21913 6199 21971 6205
rect 22094 6196 22100 6208
rect 22152 6236 22158 6248
rect 22278 6236 22284 6248
rect 22152 6208 22284 6236
rect 22152 6196 22158 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22462 6236 22468 6248
rect 22423 6208 22468 6236
rect 22462 6196 22468 6208
rect 22520 6196 22526 6248
rect 28442 6196 28448 6248
rect 28500 6236 28506 6248
rect 29273 6239 29331 6245
rect 29273 6236 29285 6239
rect 28500 6208 29285 6236
rect 28500 6196 28506 6208
rect 29273 6205 29285 6208
rect 29319 6205 29331 6239
rect 30558 6236 30564 6248
rect 30471 6208 30564 6236
rect 29273 6199 29331 6205
rect 30558 6196 30564 6208
rect 30616 6236 30622 6248
rect 32125 6239 32183 6245
rect 32125 6236 32137 6239
rect 30616 6208 32137 6236
rect 30616 6196 30622 6208
rect 32125 6205 32137 6208
rect 32171 6205 32183 6239
rect 32125 6199 32183 6205
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 23845 6171 23903 6177
rect 23845 6168 23857 6171
rect 23523 6140 23857 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23845 6137 23857 6140
rect 23891 6168 23903 6171
rect 23934 6168 23940 6180
rect 23891 6140 23940 6168
rect 23891 6137 23903 6140
rect 23845 6131 23903 6137
rect 23934 6128 23940 6140
rect 23992 6128 23998 6180
rect 25409 6171 25467 6177
rect 25409 6137 25421 6171
rect 25455 6168 25467 6171
rect 26418 6168 26424 6180
rect 25455 6140 26424 6168
rect 25455 6137 25467 6140
rect 25409 6131 25467 6137
rect 21358 6100 21364 6112
rect 21319 6072 21364 6100
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 23106 6100 23112 6112
rect 23067 6072 23112 6100
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 24670 6100 24676 6112
rect 24631 6072 24676 6100
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 25130 6100 25136 6112
rect 25091 6072 25136 6100
rect 25130 6060 25136 6072
rect 25188 6100 25194 6112
rect 25424 6100 25452 6131
rect 26418 6128 26424 6140
rect 26476 6168 26482 6180
rect 26605 6171 26663 6177
rect 26605 6168 26617 6171
rect 26476 6140 26617 6168
rect 26476 6128 26482 6140
rect 26605 6137 26617 6140
rect 26651 6168 26663 6171
rect 26973 6171 27031 6177
rect 26973 6168 26985 6171
rect 26651 6140 26985 6168
rect 26651 6137 26663 6140
rect 26605 6131 26663 6137
rect 26973 6137 26985 6140
rect 27019 6137 27031 6171
rect 26973 6131 27031 6137
rect 30282 6128 30288 6180
rect 30340 6168 30346 6180
rect 30882 6171 30940 6177
rect 30882 6168 30894 6171
rect 30340 6140 30894 6168
rect 30340 6128 30346 6140
rect 30882 6137 30894 6140
rect 30928 6137 30940 6171
rect 33244 6168 33272 6276
rect 33318 6264 33324 6276
rect 33376 6264 33382 6316
rect 41046 6304 41052 6316
rect 41007 6276 41052 6304
rect 41046 6264 41052 6276
rect 41104 6264 41110 6316
rect 41506 6304 41512 6316
rect 41467 6276 41512 6304
rect 41506 6264 41512 6276
rect 41564 6264 41570 6316
rect 42766 6304 42794 6412
rect 43438 6400 43444 6452
rect 43496 6440 43502 6452
rect 44545 6443 44603 6449
rect 44545 6440 44557 6443
rect 43496 6412 44557 6440
rect 43496 6400 43502 6412
rect 44545 6409 44557 6412
rect 44591 6409 44603 6443
rect 45186 6440 45192 6452
rect 45147 6412 45192 6440
rect 44545 6403 44603 6409
rect 45186 6400 45192 6412
rect 45244 6400 45250 6452
rect 46290 6400 46296 6452
rect 46348 6440 46354 6452
rect 47121 6443 47179 6449
rect 47121 6440 47133 6443
rect 46348 6412 47133 6440
rect 46348 6400 46354 6412
rect 47121 6409 47133 6412
rect 47167 6409 47179 6443
rect 47121 6403 47179 6409
rect 44913 6375 44971 6381
rect 44913 6341 44925 6375
rect 44959 6341 44971 6375
rect 44913 6335 44971 6341
rect 43257 6307 43315 6313
rect 43257 6304 43269 6307
rect 42766 6276 43269 6304
rect 43257 6273 43269 6276
rect 43303 6273 43315 6307
rect 43898 6304 43904 6316
rect 43859 6276 43904 6304
rect 43257 6267 43315 6273
rect 43898 6264 43904 6276
rect 43956 6264 43962 6316
rect 33410 6236 33416 6248
rect 33371 6208 33416 6236
rect 33410 6196 33416 6208
rect 33468 6196 33474 6248
rect 33689 6239 33747 6245
rect 33689 6205 33701 6239
rect 33735 6205 33747 6239
rect 33689 6199 33747 6205
rect 34952 6239 35010 6245
rect 34952 6205 34964 6239
rect 34998 6236 35010 6239
rect 35250 6236 35256 6248
rect 34998 6208 35256 6236
rect 34998 6205 35010 6208
rect 34952 6199 35010 6205
rect 33704 6168 33732 6199
rect 35250 6196 35256 6208
rect 35308 6196 35314 6248
rect 38286 6196 38292 6248
rect 38344 6236 38350 6248
rect 38473 6239 38531 6245
rect 38473 6236 38485 6239
rect 38344 6208 38485 6236
rect 38344 6196 38350 6208
rect 38473 6205 38485 6208
rect 38519 6205 38531 6239
rect 38473 6199 38531 6205
rect 38562 6196 38568 6248
rect 38620 6236 38626 6248
rect 38933 6239 38991 6245
rect 38933 6236 38945 6239
rect 38620 6208 38945 6236
rect 38620 6196 38626 6208
rect 38933 6205 38945 6208
rect 38979 6205 38991 6239
rect 38933 6199 38991 6205
rect 39114 6196 39120 6248
rect 39172 6236 39178 6248
rect 39577 6239 39635 6245
rect 39577 6236 39589 6239
rect 39172 6208 39589 6236
rect 39172 6196 39178 6208
rect 39577 6205 39589 6208
rect 39623 6236 39635 6239
rect 44726 6236 44732 6248
rect 39623 6208 40908 6236
rect 44687 6208 44732 6236
rect 39623 6205 39635 6208
rect 39577 6199 39635 6205
rect 33962 6168 33968 6180
rect 33244 6140 33732 6168
rect 33923 6140 33968 6168
rect 30882 6131 30940 6137
rect 33962 6128 33968 6140
rect 34020 6128 34026 6180
rect 36170 6168 36176 6180
rect 36131 6140 36176 6168
rect 36170 6128 36176 6140
rect 36228 6128 36234 6180
rect 36265 6171 36323 6177
rect 36265 6137 36277 6171
rect 36311 6168 36323 6171
rect 36446 6168 36452 6180
rect 36311 6140 36452 6168
rect 36311 6137 36323 6140
rect 36265 6131 36323 6137
rect 25188 6072 25452 6100
rect 29457 6103 29515 6109
rect 25188 6060 25194 6072
rect 29457 6069 29469 6103
rect 29503 6100 29515 6103
rect 29822 6100 29828 6112
rect 29503 6072 29828 6100
rect 29503 6069 29515 6072
rect 29457 6063 29515 6069
rect 29822 6060 29828 6072
rect 29880 6060 29886 6112
rect 30098 6100 30104 6112
rect 30059 6072 30104 6100
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 31478 6100 31484 6112
rect 31439 6072 31484 6100
rect 31478 6060 31484 6072
rect 31536 6060 31542 6112
rect 33410 6060 33416 6112
rect 33468 6100 33474 6112
rect 34241 6103 34299 6109
rect 34241 6100 34253 6103
rect 33468 6072 34253 6100
rect 33468 6060 33474 6072
rect 34241 6069 34253 6072
rect 34287 6069 34299 6103
rect 34241 6063 34299 6069
rect 35621 6103 35679 6109
rect 35621 6069 35633 6103
rect 35667 6100 35679 6103
rect 35802 6100 35808 6112
rect 35667 6072 35808 6100
rect 35667 6069 35679 6072
rect 35621 6063 35679 6069
rect 35802 6060 35808 6072
rect 35860 6100 35866 6112
rect 35989 6103 36047 6109
rect 35989 6100 36001 6103
rect 35860 6072 36001 6100
rect 35860 6060 35866 6072
rect 35989 6069 36001 6072
rect 36035 6100 36047 6103
rect 36280 6100 36308 6131
rect 36446 6128 36452 6140
rect 36504 6128 36510 6180
rect 36817 6171 36875 6177
rect 36817 6137 36829 6171
rect 36863 6168 36875 6171
rect 36906 6168 36912 6180
rect 36863 6140 36912 6168
rect 36863 6137 36875 6140
rect 36817 6131 36875 6137
rect 36906 6128 36912 6140
rect 36964 6128 36970 6180
rect 39209 6171 39267 6177
rect 39209 6137 39221 6171
rect 39255 6168 39267 6171
rect 40126 6168 40132 6180
rect 39255 6140 40132 6168
rect 39255 6137 39267 6140
rect 39209 6131 39267 6137
rect 40126 6128 40132 6140
rect 40184 6128 40190 6180
rect 40880 6177 40908 6208
rect 44726 6196 44732 6208
rect 44784 6196 44790 6248
rect 44928 6236 44956 6335
rect 46106 6236 46112 6248
rect 44928 6208 46112 6236
rect 46106 6196 46112 6208
rect 46164 6236 46170 6248
rect 46201 6239 46259 6245
rect 46201 6236 46213 6239
rect 46164 6208 46213 6236
rect 46164 6196 46170 6208
rect 46201 6205 46213 6208
rect 46247 6205 46259 6239
rect 46201 6199 46259 6205
rect 40865 6171 40923 6177
rect 40865 6137 40877 6171
rect 40911 6168 40923 6171
rect 41141 6171 41199 6177
rect 41141 6168 41153 6171
rect 40911 6140 41153 6168
rect 40911 6137 40923 6140
rect 40865 6131 40923 6137
rect 41141 6137 41153 6140
rect 41187 6168 41199 6171
rect 41690 6168 41696 6180
rect 41187 6140 41696 6168
rect 41187 6137 41199 6140
rect 41141 6131 41199 6137
rect 41690 6128 41696 6140
rect 41748 6168 41754 6180
rect 41966 6168 41972 6180
rect 41748 6140 41972 6168
rect 41748 6128 41754 6140
rect 41966 6128 41972 6140
rect 42024 6128 42030 6180
rect 43073 6171 43131 6177
rect 43073 6137 43085 6171
rect 43119 6168 43131 6171
rect 43349 6171 43407 6177
rect 43349 6168 43361 6171
rect 43119 6140 43361 6168
rect 43119 6137 43131 6140
rect 43073 6131 43131 6137
rect 43349 6137 43361 6140
rect 43395 6168 43407 6171
rect 43438 6168 43444 6180
rect 43395 6140 43444 6168
rect 43395 6137 43407 6140
rect 43349 6131 43407 6137
rect 43438 6128 43444 6140
rect 43496 6128 43502 6180
rect 43530 6128 43536 6180
rect 43588 6168 43594 6180
rect 44269 6171 44327 6177
rect 44269 6168 44281 6171
rect 43588 6140 44281 6168
rect 43588 6128 43594 6140
rect 44269 6137 44281 6140
rect 44315 6168 44327 6171
rect 44315 6140 45876 6168
rect 44315 6137 44327 6140
rect 44269 6131 44327 6137
rect 36035 6072 36308 6100
rect 36035 6069 36047 6072
rect 35989 6063 36047 6069
rect 39758 6060 39764 6112
rect 39816 6100 39822 6112
rect 40221 6103 40279 6109
rect 40221 6100 40233 6103
rect 39816 6072 40233 6100
rect 39816 6060 39822 6072
rect 40221 6069 40233 6072
rect 40267 6100 40279 6103
rect 40678 6100 40684 6112
rect 40267 6072 40684 6100
rect 40267 6069 40279 6072
rect 40221 6063 40279 6069
rect 40678 6060 40684 6072
rect 40736 6060 40742 6112
rect 44726 6060 44732 6112
rect 44784 6100 44790 6112
rect 45370 6100 45376 6112
rect 44784 6072 45376 6100
rect 44784 6060 44790 6072
rect 45370 6060 45376 6072
rect 45428 6100 45434 6112
rect 45557 6103 45615 6109
rect 45557 6100 45569 6103
rect 45428 6072 45569 6100
rect 45428 6060 45434 6072
rect 45557 6069 45569 6072
rect 45603 6069 45615 6103
rect 45848 6100 45876 6140
rect 46385 6103 46443 6109
rect 46385 6100 46397 6103
rect 45848 6072 46397 6100
rect 45557 6063 45615 6069
rect 46385 6069 46397 6072
rect 46431 6069 46443 6103
rect 46385 6063 46443 6069
rect 1104 6010 48852 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 48852 6010
rect 1104 5936 48852 5958
rect 23293 5899 23351 5905
rect 23293 5865 23305 5899
rect 23339 5896 23351 5899
rect 24670 5896 24676 5908
rect 23339 5868 24676 5896
rect 23339 5865 23351 5868
rect 23293 5859 23351 5865
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 27982 5896 27988 5908
rect 27943 5868 27988 5896
rect 27982 5856 27988 5868
rect 28040 5856 28046 5908
rect 30558 5896 30564 5908
rect 30519 5868 30564 5896
rect 30558 5856 30564 5868
rect 30616 5856 30622 5908
rect 31018 5856 31024 5908
rect 31076 5896 31082 5908
rect 31389 5899 31447 5905
rect 31389 5896 31401 5899
rect 31076 5868 31401 5896
rect 31076 5856 31082 5868
rect 31389 5865 31401 5868
rect 31435 5896 31447 5899
rect 32217 5899 32275 5905
rect 32217 5896 32229 5899
rect 31435 5868 32229 5896
rect 31435 5865 31447 5868
rect 31389 5859 31447 5865
rect 32217 5865 32229 5868
rect 32263 5865 32275 5899
rect 34790 5896 34796 5908
rect 34751 5868 34796 5896
rect 32217 5859 32275 5865
rect 34790 5856 34796 5868
rect 34848 5856 34854 5908
rect 35434 5856 35440 5908
rect 35492 5896 35498 5908
rect 35621 5899 35679 5905
rect 35621 5896 35633 5899
rect 35492 5868 35633 5896
rect 35492 5856 35498 5868
rect 35621 5865 35633 5868
rect 35667 5865 35679 5899
rect 35621 5859 35679 5865
rect 39022 5856 39028 5908
rect 39080 5896 39086 5908
rect 39117 5899 39175 5905
rect 39117 5896 39129 5899
rect 39080 5868 39129 5896
rect 39080 5856 39086 5868
rect 39117 5865 39129 5868
rect 39163 5865 39175 5899
rect 39117 5859 39175 5865
rect 39574 5856 39580 5908
rect 39632 5896 39638 5908
rect 39669 5899 39727 5905
rect 39669 5896 39681 5899
rect 39632 5868 39681 5896
rect 39632 5856 39638 5868
rect 39669 5865 39681 5868
rect 39715 5865 39727 5899
rect 39669 5859 39727 5865
rect 22735 5831 22793 5837
rect 22735 5797 22747 5831
rect 22781 5828 22793 5831
rect 23106 5828 23112 5840
rect 22781 5800 23112 5828
rect 22781 5797 22793 5800
rect 22735 5791 22793 5797
rect 23106 5788 23112 5800
rect 23164 5788 23170 5840
rect 24305 5831 24363 5837
rect 24305 5797 24317 5831
rect 24351 5828 24363 5831
rect 24394 5828 24400 5840
rect 24351 5800 24400 5828
rect 24351 5797 24363 5800
rect 24305 5791 24363 5797
rect 24394 5788 24400 5800
rect 24452 5788 24458 5840
rect 24854 5828 24860 5840
rect 24815 5800 24860 5828
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 27062 5788 27068 5840
rect 27120 5828 27126 5840
rect 27157 5831 27215 5837
rect 27157 5828 27169 5831
rect 27120 5800 27169 5828
rect 27120 5788 27126 5800
rect 27157 5797 27169 5800
rect 27203 5828 27215 5831
rect 28166 5828 28172 5840
rect 27203 5800 28172 5828
rect 27203 5797 27215 5800
rect 27157 5791 27215 5797
rect 28166 5788 28172 5800
rect 28224 5788 28230 5840
rect 28534 5788 28540 5840
rect 28592 5828 28598 5840
rect 28899 5831 28957 5837
rect 28899 5828 28911 5831
rect 28592 5800 28911 5828
rect 28592 5788 28598 5800
rect 28899 5797 28911 5800
rect 28945 5828 28957 5831
rect 30282 5828 30288 5840
rect 28945 5800 30288 5828
rect 28945 5797 28957 5800
rect 28899 5791 28957 5797
rect 30282 5788 30288 5800
rect 30340 5788 30346 5840
rect 33042 5828 33048 5840
rect 32416 5800 33048 5828
rect 21428 5763 21486 5769
rect 21428 5729 21440 5763
rect 21474 5760 21486 5763
rect 21542 5760 21548 5772
rect 21474 5732 21548 5760
rect 21474 5729 21486 5732
rect 21428 5723 21486 5729
rect 21542 5720 21548 5732
rect 21600 5760 21606 5772
rect 23382 5760 23388 5772
rect 21600 5732 23388 5760
rect 21600 5720 21606 5732
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 30466 5760 30472 5772
rect 30427 5732 30472 5760
rect 30466 5720 30472 5732
rect 30524 5720 30530 5772
rect 30834 5760 30840 5772
rect 30795 5732 30840 5760
rect 30834 5720 30840 5732
rect 30892 5720 30898 5772
rect 32306 5720 32312 5772
rect 32364 5760 32370 5772
rect 32416 5769 32444 5800
rect 33042 5788 33048 5800
rect 33100 5788 33106 5840
rect 37921 5831 37979 5837
rect 37921 5797 37933 5831
rect 37967 5828 37979 5831
rect 38010 5828 38016 5840
rect 37967 5800 38016 5828
rect 37967 5797 37979 5800
rect 37921 5791 37979 5797
rect 38010 5788 38016 5800
rect 38068 5828 38074 5840
rect 38930 5828 38936 5840
rect 38068 5800 38936 5828
rect 38068 5788 38074 5800
rect 38930 5788 38936 5800
rect 38988 5788 38994 5840
rect 39684 5828 39712 5859
rect 40218 5856 40224 5908
rect 40276 5896 40282 5908
rect 40497 5899 40555 5905
rect 40497 5896 40509 5899
rect 40276 5868 40509 5896
rect 40276 5856 40282 5868
rect 40497 5865 40509 5868
rect 40543 5865 40555 5899
rect 40862 5896 40868 5908
rect 40823 5868 40868 5896
rect 40497 5859 40555 5865
rect 40862 5856 40868 5868
rect 40920 5856 40926 5908
rect 41138 5856 41144 5908
rect 41196 5896 41202 5908
rect 41969 5899 42027 5905
rect 41969 5896 41981 5899
rect 41196 5868 41981 5896
rect 41196 5856 41202 5868
rect 41969 5865 41981 5868
rect 42015 5865 42027 5899
rect 41969 5859 42027 5865
rect 43898 5856 43904 5908
rect 43956 5896 43962 5908
rect 44729 5899 44787 5905
rect 44729 5896 44741 5899
rect 43956 5868 44741 5896
rect 43956 5856 43962 5868
rect 44729 5865 44741 5868
rect 44775 5865 44787 5899
rect 46106 5896 46112 5908
rect 46067 5868 46112 5896
rect 44729 5859 44787 5865
rect 46106 5856 46112 5868
rect 46164 5856 46170 5908
rect 41411 5831 41469 5837
rect 41411 5828 41423 5831
rect 39684 5800 41423 5828
rect 41411 5797 41423 5800
rect 41457 5828 41469 5831
rect 41874 5828 41880 5840
rect 41457 5800 41880 5828
rect 41457 5797 41469 5800
rect 41411 5791 41469 5797
rect 41874 5788 41880 5800
rect 41932 5788 41938 5840
rect 43438 5788 43444 5840
rect 43496 5828 43502 5840
rect 43533 5831 43591 5837
rect 43533 5828 43545 5831
rect 43496 5800 43545 5828
rect 43496 5788 43502 5800
rect 43533 5797 43545 5800
rect 43579 5828 43591 5831
rect 44913 5831 44971 5837
rect 44913 5828 44925 5831
rect 43579 5800 44925 5828
rect 43579 5797 43591 5800
rect 43533 5791 43591 5797
rect 44913 5797 44925 5800
rect 44959 5797 44971 5831
rect 44913 5791 44971 5797
rect 32401 5763 32459 5769
rect 32401 5760 32413 5763
rect 32364 5732 32413 5760
rect 32364 5720 32370 5732
rect 32401 5729 32413 5732
rect 32447 5729 32459 5763
rect 32674 5760 32680 5772
rect 32635 5732 32680 5760
rect 32401 5723 32459 5729
rect 32674 5720 32680 5732
rect 32732 5720 32738 5772
rect 33962 5720 33968 5772
rect 34020 5760 34026 5772
rect 34425 5763 34483 5769
rect 34425 5760 34437 5763
rect 34020 5732 34437 5760
rect 34020 5720 34026 5732
rect 34425 5729 34437 5732
rect 34471 5729 34483 5763
rect 34425 5723 34483 5729
rect 35345 5763 35403 5769
rect 35345 5729 35357 5763
rect 35391 5760 35403 5763
rect 36208 5763 36266 5769
rect 36208 5760 36220 5763
rect 35391 5732 36220 5760
rect 35391 5729 35403 5732
rect 35345 5723 35403 5729
rect 36208 5729 36220 5732
rect 36254 5760 36266 5763
rect 36354 5760 36360 5772
rect 36254 5732 36360 5760
rect 36254 5729 36266 5732
rect 36208 5723 36266 5729
rect 36354 5720 36360 5732
rect 36412 5720 36418 5772
rect 45002 5760 45008 5772
rect 44963 5732 45008 5760
rect 45002 5720 45008 5732
rect 45060 5720 45066 5772
rect 22370 5692 22376 5704
rect 22331 5664 22376 5692
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 24210 5692 24216 5704
rect 23446 5664 24216 5692
rect 21499 5627 21557 5633
rect 21499 5593 21511 5627
rect 21545 5624 21557 5627
rect 23446 5624 23474 5664
rect 24210 5652 24216 5664
rect 24268 5652 24274 5704
rect 27065 5695 27123 5701
rect 27065 5661 27077 5695
rect 27111 5661 27123 5695
rect 27338 5692 27344 5704
rect 27299 5664 27344 5692
rect 27065 5655 27123 5661
rect 21545 5596 23474 5624
rect 21545 5593 21557 5596
rect 21499 5587 21557 5593
rect 26326 5584 26332 5636
rect 26384 5624 26390 5636
rect 27080 5624 27108 5655
rect 27338 5652 27344 5664
rect 27396 5652 27402 5704
rect 28442 5652 28448 5704
rect 28500 5692 28506 5704
rect 28537 5695 28595 5701
rect 28537 5692 28549 5695
rect 28500 5664 28549 5692
rect 28500 5652 28506 5664
rect 28537 5661 28549 5664
rect 28583 5661 28595 5695
rect 28537 5655 28595 5661
rect 37458 5652 37464 5704
rect 37516 5692 37522 5704
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 37516 5664 37841 5692
rect 37516 5652 37522 5664
rect 37829 5661 37841 5664
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 38473 5695 38531 5701
rect 38473 5661 38485 5695
rect 38519 5692 38531 5695
rect 39114 5692 39120 5704
rect 38519 5664 39120 5692
rect 38519 5661 38531 5664
rect 38473 5655 38531 5661
rect 39114 5652 39120 5664
rect 39172 5652 39178 5704
rect 39298 5692 39304 5704
rect 39259 5664 39304 5692
rect 39298 5652 39304 5664
rect 39356 5652 39362 5704
rect 40126 5652 40132 5704
rect 40184 5692 40190 5704
rect 41049 5695 41107 5701
rect 41049 5692 41061 5695
rect 40184 5664 41061 5692
rect 40184 5652 40190 5664
rect 41049 5661 41061 5664
rect 41095 5661 41107 5695
rect 41049 5655 41107 5661
rect 41506 5652 41512 5704
rect 41564 5692 41570 5704
rect 43070 5692 43076 5704
rect 41564 5664 43076 5692
rect 41564 5652 41570 5664
rect 43070 5652 43076 5664
rect 43128 5692 43134 5704
rect 43441 5695 43499 5701
rect 43441 5692 43453 5695
rect 43128 5664 43453 5692
rect 43128 5652 43134 5664
rect 43441 5661 43453 5664
rect 43487 5661 43499 5695
rect 44082 5692 44088 5704
rect 44043 5664 44088 5692
rect 43441 5655 43499 5661
rect 44082 5652 44088 5664
rect 44140 5652 44146 5704
rect 29638 5624 29644 5636
rect 26384 5596 29644 5624
rect 26384 5584 26390 5596
rect 29638 5584 29644 5596
rect 29696 5584 29702 5636
rect 38841 5627 38899 5633
rect 38841 5593 38853 5627
rect 38887 5624 38899 5627
rect 39022 5624 39028 5636
rect 38887 5596 39028 5624
rect 38887 5593 38899 5596
rect 38841 5587 38899 5593
rect 39022 5584 39028 5596
rect 39080 5624 39086 5636
rect 39666 5624 39672 5636
rect 39080 5596 39672 5624
rect 39080 5584 39086 5596
rect 39666 5584 39672 5596
rect 39724 5584 39730 5636
rect 22097 5559 22155 5565
rect 22097 5525 22109 5559
rect 22143 5556 22155 5559
rect 22462 5556 22468 5568
rect 22143 5528 22468 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 23750 5556 23756 5568
rect 23711 5528 23756 5556
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 25314 5556 25320 5568
rect 25275 5528 25320 5556
rect 25314 5516 25320 5528
rect 25372 5516 25378 5568
rect 26878 5556 26884 5568
rect 26839 5528 26884 5556
rect 26878 5516 26884 5528
rect 26936 5516 26942 5568
rect 29454 5556 29460 5568
rect 29415 5528 29460 5556
rect 29454 5516 29460 5528
rect 29512 5516 29518 5568
rect 33321 5559 33379 5565
rect 33321 5525 33333 5559
rect 33367 5556 33379 5559
rect 33410 5556 33416 5568
rect 33367 5528 33416 5556
rect 33367 5525 33379 5528
rect 33321 5519 33379 5525
rect 33410 5516 33416 5528
rect 33468 5516 33474 5568
rect 36311 5559 36369 5565
rect 36311 5525 36323 5559
rect 36357 5556 36369 5559
rect 36814 5556 36820 5568
rect 36357 5528 36820 5556
rect 36357 5525 36369 5528
rect 36311 5519 36369 5525
rect 36814 5516 36820 5528
rect 36872 5516 36878 5568
rect 36998 5556 37004 5568
rect 36959 5528 37004 5556
rect 36998 5516 37004 5528
rect 37056 5516 37062 5568
rect 40218 5556 40224 5568
rect 40179 5528 40224 5556
rect 40218 5516 40224 5528
rect 40276 5516 40282 5568
rect 43806 5516 43812 5568
rect 43864 5556 43870 5568
rect 44361 5559 44419 5565
rect 44361 5556 44373 5559
rect 43864 5528 44373 5556
rect 43864 5516 43870 5528
rect 44361 5525 44373 5528
rect 44407 5525 44419 5559
rect 44361 5519 44419 5525
rect 1104 5466 48852 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 48852 5466
rect 1104 5392 48852 5414
rect 20346 5352 20352 5364
rect 20307 5324 20352 5352
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 21542 5352 21548 5364
rect 21503 5324 21548 5352
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 21910 5352 21916 5364
rect 21871 5324 21916 5352
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23842 5352 23848 5364
rect 23523 5324 23848 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23842 5312 23848 5324
rect 23900 5352 23906 5364
rect 24394 5352 24400 5364
rect 23900 5324 24400 5352
rect 23900 5312 23906 5324
rect 24394 5312 24400 5324
rect 24452 5352 24458 5364
rect 24670 5352 24676 5364
rect 24452 5324 24676 5352
rect 24452 5312 24458 5324
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 27893 5355 27951 5361
rect 27893 5321 27905 5355
rect 27939 5352 27951 5355
rect 28166 5352 28172 5364
rect 27939 5324 28172 5352
rect 27939 5321 27951 5324
rect 27893 5315 27951 5321
rect 28166 5312 28172 5324
rect 28224 5312 28230 5364
rect 28534 5352 28540 5364
rect 28495 5324 28540 5352
rect 28534 5312 28540 5324
rect 28592 5312 28598 5364
rect 30377 5355 30435 5361
rect 30377 5321 30389 5355
rect 30423 5352 30435 5355
rect 30466 5352 30472 5364
rect 30423 5324 30472 5352
rect 30423 5321 30435 5324
rect 30377 5315 30435 5321
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 32306 5352 32312 5364
rect 32267 5324 32312 5352
rect 32306 5312 32312 5324
rect 32364 5312 32370 5364
rect 33962 5312 33968 5364
rect 34020 5352 34026 5364
rect 34057 5355 34115 5361
rect 34057 5352 34069 5355
rect 34020 5324 34069 5352
rect 34020 5312 34026 5324
rect 34057 5321 34069 5324
rect 34103 5321 34115 5355
rect 36354 5352 36360 5364
rect 36315 5324 36360 5352
rect 34057 5315 34115 5321
rect 36354 5312 36360 5324
rect 36412 5312 36418 5364
rect 36446 5312 36452 5364
rect 36504 5352 36510 5364
rect 36817 5355 36875 5361
rect 36817 5352 36829 5355
rect 36504 5324 36829 5352
rect 36504 5312 36510 5324
rect 36817 5321 36829 5324
rect 36863 5352 36875 5355
rect 37090 5352 37096 5364
rect 36863 5324 37096 5352
rect 36863 5321 36875 5324
rect 36817 5315 36875 5321
rect 37090 5312 37096 5324
rect 37148 5352 37154 5364
rect 38010 5352 38016 5364
rect 37148 5324 38016 5352
rect 37148 5312 37154 5324
rect 38010 5312 38016 5324
rect 38068 5312 38074 5364
rect 38286 5352 38292 5364
rect 38247 5324 38292 5352
rect 38286 5312 38292 5324
rect 38344 5312 38350 5364
rect 39574 5352 39580 5364
rect 39535 5324 39580 5352
rect 39574 5312 39580 5324
rect 39632 5312 39638 5364
rect 40218 5312 40224 5364
rect 40276 5352 40282 5364
rect 42245 5355 42303 5361
rect 42245 5352 42257 5355
rect 40276 5324 42257 5352
rect 40276 5312 40282 5324
rect 42245 5321 42257 5324
rect 42291 5321 42303 5355
rect 42245 5315 42303 5321
rect 21358 5244 21364 5296
rect 21416 5284 21422 5296
rect 34606 5284 34612 5296
rect 21416 5256 27200 5284
rect 21416 5244 21422 5256
rect 20530 5216 20536 5228
rect 20491 5188 20536 5216
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21726 5216 21732 5228
rect 21223 5188 21732 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 22370 5176 22376 5228
rect 22428 5216 22434 5228
rect 22557 5219 22615 5225
rect 22557 5216 22569 5219
rect 22428 5188 22569 5216
rect 22428 5176 22434 5188
rect 22557 5185 22569 5188
rect 22603 5185 22615 5219
rect 23750 5216 23756 5228
rect 23711 5188 23756 5216
rect 22557 5179 22615 5185
rect 23750 5176 23756 5188
rect 23808 5176 23814 5228
rect 24394 5216 24400 5228
rect 24307 5188 24400 5216
rect 24394 5176 24400 5188
rect 24452 5216 24458 5228
rect 25314 5216 25320 5228
rect 24452 5188 25320 5216
rect 24452 5176 24458 5188
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 25608 5225 25636 5256
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5185 25651 5219
rect 26878 5216 26884 5228
rect 26839 5188 26884 5216
rect 25593 5179 25651 5185
rect 26878 5176 26884 5188
rect 26936 5176 26942 5228
rect 27172 5225 27200 5256
rect 29564 5256 34612 5284
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 22005 5151 22063 5157
rect 22005 5148 22017 5151
rect 21968 5120 22017 5148
rect 21968 5108 21974 5120
rect 22005 5117 22017 5120
rect 22051 5148 22063 5151
rect 22094 5148 22100 5160
rect 22051 5120 22100 5148
rect 22051 5117 22063 5120
rect 22005 5111 22063 5117
rect 22094 5108 22100 5120
rect 22152 5108 22158 5160
rect 22462 5148 22468 5160
rect 22423 5120 22468 5148
rect 22462 5108 22468 5120
rect 22520 5148 22526 5160
rect 29564 5157 29592 5256
rect 34606 5244 34612 5256
rect 34664 5244 34670 5296
rect 40678 5284 40684 5296
rect 40639 5256 40684 5284
rect 40678 5244 40684 5256
rect 40736 5244 40742 5296
rect 40862 5244 40868 5296
rect 40920 5284 40926 5296
rect 41506 5284 41512 5296
rect 40920 5256 41000 5284
rect 41467 5256 41512 5284
rect 40920 5244 40926 5256
rect 31018 5216 31024 5228
rect 30979 5188 31024 5216
rect 31018 5176 31024 5188
rect 31076 5176 31082 5228
rect 33410 5216 33416 5228
rect 33244 5188 33416 5216
rect 29089 5151 29147 5157
rect 22520 5120 23474 5148
rect 22520 5108 22526 5120
rect 20625 5083 20683 5089
rect 20625 5049 20637 5083
rect 20671 5049 20683 5083
rect 23446 5080 23474 5120
rect 29089 5117 29101 5151
rect 29135 5148 29147 5151
rect 29549 5151 29607 5157
rect 29549 5148 29561 5151
rect 29135 5120 29561 5148
rect 29135 5117 29147 5120
rect 29089 5111 29147 5117
rect 29549 5117 29561 5120
rect 29595 5117 29607 5151
rect 29822 5148 29828 5160
rect 29735 5120 29828 5148
rect 29549 5111 29607 5117
rect 29822 5108 29828 5120
rect 29880 5148 29886 5160
rect 30834 5148 30840 5160
rect 29880 5120 30840 5148
rect 29880 5108 29886 5120
rect 30834 5108 30840 5120
rect 30892 5108 30898 5160
rect 33244 5157 33272 5188
rect 33410 5176 33416 5188
rect 33468 5176 33474 5228
rect 33594 5216 33600 5228
rect 33555 5188 33600 5216
rect 33594 5176 33600 5188
rect 33652 5176 33658 5228
rect 34698 5176 34704 5228
rect 34756 5216 34762 5228
rect 35161 5219 35219 5225
rect 35161 5216 35173 5219
rect 34756 5188 35173 5216
rect 34756 5176 34762 5188
rect 35161 5185 35173 5188
rect 35207 5216 35219 5219
rect 35526 5216 35532 5228
rect 35207 5188 35532 5216
rect 35207 5185 35219 5188
rect 35161 5179 35219 5185
rect 35526 5176 35532 5188
rect 35584 5176 35590 5228
rect 36998 5216 37004 5228
rect 36959 5188 37004 5216
rect 36998 5176 37004 5188
rect 37056 5176 37062 5228
rect 39209 5219 39267 5225
rect 39209 5185 39221 5219
rect 39255 5216 39267 5219
rect 39298 5216 39304 5228
rect 39255 5188 39304 5216
rect 39255 5185 39267 5188
rect 39209 5179 39267 5185
rect 39298 5176 39304 5188
rect 39356 5216 39362 5228
rect 39853 5219 39911 5225
rect 39853 5216 39865 5219
rect 39356 5188 39865 5216
rect 39356 5176 39362 5188
rect 39853 5185 39865 5188
rect 39899 5185 39911 5219
rect 39853 5179 39911 5185
rect 40126 5176 40132 5228
rect 40184 5216 40190 5228
rect 40972 5225 41000 5256
rect 41506 5244 41512 5256
rect 41564 5244 41570 5296
rect 41874 5284 41880 5296
rect 41835 5256 41880 5284
rect 41874 5244 41880 5256
rect 41932 5244 41938 5296
rect 40221 5219 40279 5225
rect 40221 5216 40233 5219
rect 40184 5188 40233 5216
rect 40184 5176 40190 5188
rect 40221 5185 40233 5188
rect 40267 5185 40279 5219
rect 40221 5179 40279 5185
rect 40957 5219 41015 5225
rect 40957 5185 40969 5219
rect 41003 5185 41015 5219
rect 40957 5179 41015 5185
rect 33229 5151 33287 5157
rect 33229 5117 33241 5151
rect 33275 5117 33287 5151
rect 33505 5151 33563 5157
rect 33505 5148 33517 5151
rect 33229 5111 33287 5117
rect 33336 5120 33517 5148
rect 23446 5052 23796 5080
rect 20625 5043 20683 5049
rect 20346 4972 20352 5024
rect 20404 5012 20410 5024
rect 20640 5012 20668 5043
rect 23106 5012 23112 5024
rect 20404 4984 20668 5012
rect 23067 4984 23112 5012
rect 20404 4972 20410 4984
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 23768 5012 23796 5052
rect 23842 5040 23848 5092
rect 23900 5080 23906 5092
rect 25130 5080 25136 5092
rect 23900 5052 23945 5080
rect 25043 5052 25136 5080
rect 23900 5040 23906 5052
rect 25130 5040 25136 5052
rect 25188 5080 25194 5092
rect 25409 5083 25467 5089
rect 25409 5080 25421 5083
rect 25188 5052 25421 5080
rect 25188 5040 25194 5052
rect 25409 5049 25421 5052
rect 25455 5049 25467 5083
rect 25409 5043 25467 5049
rect 26697 5083 26755 5089
rect 26697 5049 26709 5083
rect 26743 5080 26755 5083
rect 26973 5083 27031 5089
rect 26973 5080 26985 5083
rect 26743 5052 26985 5080
rect 26743 5049 26755 5052
rect 26697 5043 26755 5049
rect 26973 5049 26985 5052
rect 27019 5080 27031 5083
rect 27062 5080 27068 5092
rect 27019 5052 27068 5080
rect 27019 5049 27031 5052
rect 26973 5043 27031 5049
rect 27062 5040 27068 5052
rect 27120 5040 27126 5092
rect 28261 5083 28319 5089
rect 28261 5049 28273 5083
rect 28307 5080 28319 5083
rect 28442 5080 28448 5092
rect 28307 5052 28448 5080
rect 28307 5049 28319 5052
rect 28261 5043 28319 5049
rect 28442 5040 28448 5052
rect 28500 5080 28506 5092
rect 30929 5083 30987 5089
rect 28500 5052 29408 5080
rect 28500 5040 28506 5052
rect 24578 5012 24584 5024
rect 23768 4984 24584 5012
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 29380 5021 29408 5052
rect 30929 5049 30941 5083
rect 30975 5080 30987 5083
rect 31018 5080 31024 5092
rect 30975 5052 31024 5080
rect 30975 5049 30987 5052
rect 30929 5043 30987 5049
rect 31018 5040 31024 5052
rect 31076 5080 31082 5092
rect 31342 5083 31400 5089
rect 31342 5080 31354 5083
rect 31076 5052 31354 5080
rect 31076 5040 31082 5052
rect 31342 5049 31354 5052
rect 31388 5049 31400 5083
rect 31342 5043 31400 5049
rect 33042 5040 33048 5092
rect 33100 5080 33106 5092
rect 33336 5080 33364 5120
rect 33505 5117 33517 5120
rect 33551 5117 33563 5151
rect 33505 5111 33563 5117
rect 38286 5108 38292 5160
rect 38344 5148 38350 5160
rect 38473 5151 38531 5157
rect 38473 5148 38485 5151
rect 38344 5120 38485 5148
rect 38344 5108 38350 5120
rect 38473 5117 38485 5120
rect 38519 5117 38531 5151
rect 39022 5148 39028 5160
rect 38983 5120 39028 5148
rect 38473 5111 38531 5117
rect 39022 5108 39028 5120
rect 39080 5108 39086 5160
rect 42260 5148 42288 5315
rect 42334 5312 42340 5364
rect 42392 5352 42398 5364
rect 42567 5355 42625 5361
rect 42567 5352 42579 5355
rect 42392 5324 42579 5352
rect 42392 5312 42398 5324
rect 42567 5321 42579 5324
rect 42613 5321 42625 5355
rect 43438 5352 43444 5364
rect 43399 5324 43444 5352
rect 42567 5315 42625 5321
rect 43438 5312 43444 5324
rect 43496 5312 43502 5364
rect 45002 5352 45008 5364
rect 44963 5324 45008 5352
rect 45002 5312 45008 5324
rect 45060 5312 45066 5364
rect 43806 5216 43812 5228
rect 43767 5188 43812 5216
rect 43806 5176 43812 5188
rect 43864 5176 43870 5228
rect 42464 5151 42522 5157
rect 42464 5148 42476 5151
rect 42260 5120 42476 5148
rect 42464 5117 42476 5120
rect 42510 5117 42522 5151
rect 42464 5111 42522 5117
rect 34790 5080 34796 5092
rect 33100 5052 33364 5080
rect 34440 5052 34796 5080
rect 33100 5040 33106 5052
rect 29365 5015 29423 5021
rect 29365 4981 29377 5015
rect 29411 4981 29423 5015
rect 31938 5012 31944 5024
rect 31899 4984 31944 5012
rect 29365 4975 29423 4981
rect 31938 4972 31944 4984
rect 31996 4972 32002 5024
rect 32953 5015 33011 5021
rect 32953 4981 32965 5015
rect 32999 5012 33011 5015
rect 33410 5012 33416 5024
rect 32999 4984 33416 5012
rect 32999 4981 33011 4984
rect 32953 4975 33011 4981
rect 33410 4972 33416 4984
rect 33468 4972 33474 5024
rect 33686 4972 33692 5024
rect 33744 5012 33750 5024
rect 34440 5021 34468 5052
rect 34790 5040 34796 5052
rect 34848 5080 34854 5092
rect 35482 5083 35540 5089
rect 35482 5080 35494 5083
rect 34848 5052 35494 5080
rect 34848 5040 34854 5052
rect 35482 5049 35494 5052
rect 35528 5049 35540 5083
rect 37090 5080 37096 5092
rect 37051 5052 37096 5080
rect 35482 5043 35540 5049
rect 37090 5040 37096 5052
rect 37148 5040 37154 5092
rect 37642 5080 37648 5092
rect 37603 5052 37648 5080
rect 37642 5040 37648 5052
rect 37700 5040 37706 5092
rect 37734 5040 37740 5092
rect 37792 5080 37798 5092
rect 39040 5080 39068 5108
rect 37792 5052 39068 5080
rect 37792 5040 37798 5052
rect 40678 5040 40684 5092
rect 40736 5080 40742 5092
rect 41049 5083 41107 5089
rect 41049 5080 41061 5083
rect 40736 5052 41061 5080
rect 40736 5040 40742 5052
rect 41049 5049 41061 5052
rect 41095 5080 41107 5083
rect 41598 5080 41604 5092
rect 41095 5052 41604 5080
rect 41095 5049 41107 5052
rect 41049 5043 41107 5049
rect 41598 5040 41604 5052
rect 41656 5040 41662 5092
rect 43073 5083 43131 5089
rect 43073 5049 43085 5083
rect 43119 5080 43131 5083
rect 43530 5080 43536 5092
rect 43119 5052 43536 5080
rect 43119 5049 43131 5052
rect 43073 5043 43131 5049
rect 43530 5040 43536 5052
rect 43588 5080 43594 5092
rect 43901 5083 43959 5089
rect 43901 5080 43913 5083
rect 43588 5052 43913 5080
rect 43588 5040 43594 5052
rect 43901 5049 43913 5052
rect 43947 5049 43959 5083
rect 44450 5080 44456 5092
rect 44411 5052 44456 5080
rect 43901 5043 43959 5049
rect 44450 5040 44456 5052
rect 44508 5040 44514 5092
rect 34425 5015 34483 5021
rect 34425 5012 34437 5015
rect 33744 4984 34437 5012
rect 33744 4972 33750 4984
rect 34425 4981 34437 4984
rect 34471 4981 34483 5015
rect 36078 5012 36084 5024
rect 36039 4984 36084 5012
rect 34425 4975 34483 4981
rect 36078 4972 36084 4984
rect 36136 4972 36142 5024
rect 1104 4922 48852 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 48852 4922
rect 1104 4848 48852 4870
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 22370 4808 22376 4820
rect 22331 4780 22376 4808
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 22695 4811 22753 4817
rect 22695 4777 22707 4811
rect 22741 4808 22753 4811
rect 23658 4808 23664 4820
rect 22741 4780 23664 4808
rect 22741 4777 22753 4780
rect 22695 4771 22753 4777
rect 23658 4768 23664 4780
rect 23716 4768 23722 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 24949 4811 25007 4817
rect 24949 4808 24961 4811
rect 24268 4780 24961 4808
rect 24268 4768 24274 4780
rect 24949 4777 24961 4780
rect 24995 4777 25007 4811
rect 24949 4771 25007 4777
rect 25547 4811 25605 4817
rect 25547 4777 25559 4811
rect 25593 4808 25605 4811
rect 25958 4808 25964 4820
rect 25593 4780 25964 4808
rect 25593 4777 25605 4780
rect 25547 4771 25605 4777
rect 25958 4768 25964 4780
rect 26016 4768 26022 4820
rect 26973 4811 27031 4817
rect 26973 4777 26985 4811
rect 27019 4808 27031 4811
rect 27062 4808 27068 4820
rect 27019 4780 27068 4808
rect 27019 4777 27031 4780
rect 26973 4771 27031 4777
rect 27062 4768 27068 4780
rect 27120 4768 27126 4820
rect 28258 4808 28264 4820
rect 28171 4780 28264 4808
rect 28258 4768 28264 4780
rect 28316 4808 28322 4820
rect 29454 4808 29460 4820
rect 28316 4780 29460 4808
rect 28316 4768 28322 4780
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 29641 4811 29699 4817
rect 29641 4777 29653 4811
rect 29687 4808 29699 4811
rect 29822 4808 29828 4820
rect 29687 4780 29828 4808
rect 29687 4777 29699 4780
rect 29641 4771 29699 4777
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 30515 4811 30573 4817
rect 30515 4777 30527 4811
rect 30561 4808 30573 4811
rect 31294 4808 31300 4820
rect 30561 4780 31300 4808
rect 30561 4777 30573 4780
rect 30515 4771 30573 4777
rect 31294 4768 31300 4780
rect 31352 4768 31358 4820
rect 31754 4768 31760 4820
rect 31812 4808 31818 4820
rect 32263 4811 32321 4817
rect 32263 4808 32275 4811
rect 31812 4780 32275 4808
rect 31812 4768 31818 4780
rect 32263 4777 32275 4780
rect 32309 4777 32321 4811
rect 32674 4808 32680 4820
rect 32635 4780 32680 4808
rect 32263 4771 32321 4777
rect 32674 4768 32680 4780
rect 32732 4768 32738 4820
rect 33042 4808 33048 4820
rect 33003 4780 33048 4808
rect 33042 4768 33048 4780
rect 33100 4768 33106 4820
rect 35526 4808 35532 4820
rect 35487 4780 35532 4808
rect 35526 4768 35532 4780
rect 35584 4768 35590 4820
rect 38838 4768 38844 4820
rect 38896 4808 38902 4820
rect 39025 4811 39083 4817
rect 39025 4808 39037 4811
rect 38896 4780 39037 4808
rect 38896 4768 38902 4780
rect 39025 4777 39037 4780
rect 39071 4777 39083 4811
rect 43070 4808 43076 4820
rect 43031 4780 43076 4808
rect 39025 4771 39083 4777
rect 43070 4768 43076 4780
rect 43128 4768 43134 4820
rect 45002 4768 45008 4820
rect 45060 4808 45066 4820
rect 45327 4811 45385 4817
rect 45327 4808 45339 4811
rect 45060 4780 45339 4808
rect 45060 4768 45066 4780
rect 45327 4777 45339 4780
rect 45373 4777 45385 4811
rect 45327 4771 45385 4777
rect 23753 4743 23811 4749
rect 23753 4709 23765 4743
rect 23799 4740 23811 4743
rect 23934 4740 23940 4752
rect 23799 4712 23940 4740
rect 23799 4709 23811 4712
rect 23753 4703 23811 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 24305 4743 24363 4749
rect 24305 4709 24317 4743
rect 24351 4740 24363 4743
rect 24394 4740 24400 4752
rect 24351 4712 24400 4740
rect 24351 4709 24363 4712
rect 24305 4703 24363 4709
rect 24394 4700 24400 4712
rect 24452 4700 24458 4752
rect 24578 4740 24584 4752
rect 24539 4712 24584 4740
rect 24578 4700 24584 4712
rect 24636 4700 24642 4752
rect 28442 4700 28448 4752
rect 28500 4740 28506 4752
rect 28721 4743 28779 4749
rect 28721 4740 28733 4743
rect 28500 4712 28733 4740
rect 28500 4700 28506 4712
rect 28721 4709 28733 4712
rect 28767 4740 28779 4743
rect 30098 4740 30104 4752
rect 28767 4712 30104 4740
rect 28767 4709 28779 4712
rect 28721 4703 28779 4709
rect 30098 4700 30104 4712
rect 30156 4740 30162 4752
rect 32582 4740 32588 4752
rect 30156 4712 32588 4740
rect 30156 4700 30162 4712
rect 32582 4700 32588 4712
rect 32640 4700 32646 4752
rect 33686 4700 33692 4752
rect 33744 4740 33750 4752
rect 33918 4743 33976 4749
rect 33918 4740 33930 4743
rect 33744 4712 33930 4740
rect 33744 4700 33750 4712
rect 33918 4709 33930 4712
rect 33964 4740 33976 4743
rect 35161 4743 35219 4749
rect 35161 4740 35173 4743
rect 33964 4712 35173 4740
rect 33964 4709 33976 4712
rect 33918 4703 33976 4709
rect 35161 4709 35173 4712
rect 35207 4709 35219 4743
rect 35161 4703 35219 4709
rect 35710 4700 35716 4752
rect 35768 4740 35774 4752
rect 36265 4743 36323 4749
rect 36265 4740 36277 4743
rect 35768 4712 36277 4740
rect 35768 4700 35774 4712
rect 36265 4709 36277 4712
rect 36311 4709 36323 4743
rect 36265 4703 36323 4709
rect 36814 4700 36820 4752
rect 36872 4740 36878 4752
rect 39482 4740 39488 4752
rect 36872 4712 39488 4740
rect 36872 4700 36878 4712
rect 39482 4700 39488 4712
rect 39540 4740 39546 4752
rect 39669 4743 39727 4749
rect 39669 4740 39681 4743
rect 39540 4712 39681 4740
rect 39540 4700 39546 4712
rect 39669 4709 39681 4712
rect 39715 4709 39727 4743
rect 39669 4703 39727 4709
rect 39758 4700 39764 4752
rect 39816 4740 39822 4752
rect 39816 4712 39861 4740
rect 39816 4700 39822 4712
rect 43438 4700 43444 4752
rect 43496 4740 43502 4752
rect 43809 4743 43867 4749
rect 43809 4740 43821 4743
rect 43496 4712 43821 4740
rect 43496 4700 43502 4712
rect 43809 4709 43821 4712
rect 43855 4709 43867 4743
rect 43809 4703 43867 4709
rect 44361 4743 44419 4749
rect 44361 4709 44373 4743
rect 44407 4740 44419 4743
rect 44450 4740 44456 4752
rect 44407 4712 44456 4740
rect 44407 4709 44419 4712
rect 44361 4703 44419 4709
rect 44450 4700 44456 4712
rect 44508 4700 44514 4752
rect 22624 4675 22682 4681
rect 22624 4641 22636 4675
rect 22670 4672 22682 4675
rect 22922 4672 22928 4684
rect 22670 4644 22928 4672
rect 22670 4641 22682 4644
rect 22624 4635 22682 4641
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 25406 4672 25412 4684
rect 25367 4644 25412 4672
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 25590 4632 25596 4684
rect 25648 4672 25654 4684
rect 26605 4675 26663 4681
rect 26605 4672 26617 4675
rect 25648 4644 26617 4672
rect 25648 4632 25654 4644
rect 26605 4641 26617 4644
rect 26651 4672 26663 4675
rect 26970 4672 26976 4684
rect 26651 4644 26976 4672
rect 26651 4641 26663 4644
rect 26605 4635 26663 4641
rect 26970 4632 26976 4644
rect 27028 4632 27034 4684
rect 30444 4675 30502 4681
rect 30444 4641 30456 4675
rect 30490 4672 30502 4675
rect 30650 4672 30656 4684
rect 30490 4644 30656 4672
rect 30490 4641 30502 4644
rect 30444 4635 30502 4641
rect 30650 4632 30656 4644
rect 30708 4672 30714 4684
rect 31205 4675 31263 4681
rect 31205 4672 31217 4675
rect 30708 4644 31217 4672
rect 30708 4632 30714 4644
rect 31205 4641 31217 4644
rect 31251 4641 31263 4675
rect 31205 4635 31263 4641
rect 31478 4632 31484 4684
rect 31536 4672 31542 4684
rect 32122 4672 32128 4684
rect 32180 4681 32186 4684
rect 32180 4675 32218 4681
rect 31536 4644 32128 4672
rect 31536 4632 31542 4644
rect 32122 4632 32128 4644
rect 32206 4641 32218 4675
rect 38286 4672 38292 4684
rect 38247 4644 38292 4672
rect 32180 4635 32218 4641
rect 32180 4632 32186 4635
rect 38286 4632 38292 4644
rect 38344 4632 38350 4684
rect 38473 4675 38531 4681
rect 38473 4672 38485 4675
rect 38396 4644 38485 4672
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 23661 4607 23719 4613
rect 23661 4604 23673 4607
rect 23440 4576 23673 4604
rect 23440 4564 23446 4576
rect 23661 4573 23673 4576
rect 23707 4573 23719 4607
rect 23661 4567 23719 4573
rect 28074 4564 28080 4616
rect 28132 4604 28138 4616
rect 28629 4607 28687 4613
rect 28629 4604 28641 4607
rect 28132 4576 28641 4604
rect 28132 4564 28138 4576
rect 28629 4573 28641 4576
rect 28675 4573 28687 4607
rect 28629 4567 28687 4573
rect 29273 4607 29331 4613
rect 29273 4573 29285 4607
rect 29319 4604 29331 4607
rect 29638 4604 29644 4616
rect 29319 4576 29644 4604
rect 29319 4573 29331 4576
rect 29273 4567 29331 4573
rect 29638 4564 29644 4576
rect 29696 4564 29702 4616
rect 30834 4564 30840 4616
rect 30892 4604 30898 4616
rect 30929 4607 30987 4613
rect 30929 4604 30941 4607
rect 30892 4576 30941 4604
rect 30892 4564 30898 4576
rect 30929 4573 30941 4576
rect 30975 4604 30987 4607
rect 32674 4604 32680 4616
rect 30975 4576 32680 4604
rect 30975 4573 30987 4576
rect 30929 4567 30987 4573
rect 32674 4564 32680 4576
rect 32732 4564 32738 4616
rect 33594 4604 33600 4616
rect 33555 4576 33600 4604
rect 33594 4564 33600 4576
rect 33652 4564 33658 4616
rect 35986 4564 35992 4616
rect 36044 4604 36050 4616
rect 36173 4607 36231 4613
rect 36173 4604 36185 4607
rect 36044 4576 36185 4604
rect 36044 4564 36050 4576
rect 36173 4573 36185 4576
rect 36219 4573 36231 4607
rect 36173 4567 36231 4573
rect 36817 4607 36875 4613
rect 36817 4573 36829 4607
rect 36863 4604 36875 4607
rect 37642 4604 37648 4616
rect 36863 4576 37648 4604
rect 36863 4573 36875 4576
rect 36817 4567 36875 4573
rect 37642 4564 37648 4576
rect 37700 4564 37706 4616
rect 37918 4496 37924 4548
rect 37976 4536 37982 4548
rect 38396 4536 38424 4644
rect 38473 4641 38485 4644
rect 38519 4641 38531 4675
rect 38473 4635 38531 4641
rect 41208 4675 41266 4681
rect 41208 4641 41220 4675
rect 41254 4672 41266 4675
rect 41322 4672 41328 4684
rect 41254 4644 41328 4672
rect 41254 4641 41266 4644
rect 41208 4635 41266 4641
rect 41322 4632 41328 4644
rect 41380 4632 41386 4684
rect 42220 4675 42278 4681
rect 42220 4641 42232 4675
rect 42266 4672 42278 4675
rect 42794 4672 42800 4684
rect 42266 4644 42800 4672
rect 42266 4641 42278 4644
rect 42220 4635 42278 4641
rect 42794 4632 42800 4644
rect 42852 4632 42858 4684
rect 45256 4675 45314 4681
rect 45256 4641 45268 4675
rect 45302 4672 45314 4675
rect 45370 4672 45376 4684
rect 45302 4644 45376 4672
rect 45302 4641 45314 4644
rect 45256 4635 45314 4641
rect 45370 4632 45376 4644
rect 45428 4632 45434 4684
rect 38562 4604 38568 4616
rect 38523 4576 38568 4604
rect 38562 4564 38568 4576
rect 38620 4564 38626 4616
rect 39114 4564 39120 4616
rect 39172 4604 39178 4616
rect 39945 4607 40003 4613
rect 39945 4604 39957 4607
rect 39172 4576 39957 4604
rect 39172 4564 39178 4576
rect 39945 4573 39957 4576
rect 39991 4604 40003 4607
rect 43714 4604 43720 4616
rect 39991 4576 42794 4604
rect 43675 4576 43720 4604
rect 39991 4573 40003 4576
rect 39945 4567 40003 4573
rect 37976 4508 38424 4536
rect 37976 4496 37982 4508
rect 41782 4496 41788 4548
rect 41840 4536 41846 4548
rect 42291 4539 42349 4545
rect 42291 4536 42303 4539
rect 41840 4508 42303 4536
rect 41840 4496 41846 4508
rect 42291 4505 42303 4508
rect 42337 4505 42349 4539
rect 42766 4536 42794 4576
rect 43714 4564 43720 4576
rect 43772 4564 43778 4616
rect 43806 4536 43812 4548
rect 42766 4508 43812 4536
rect 42291 4499 42349 4505
rect 43806 4496 43812 4508
rect 43864 4496 43870 4548
rect 22097 4471 22155 4477
rect 22097 4437 22109 4471
rect 22143 4468 22155 4471
rect 22462 4468 22468 4480
rect 22143 4440 22468 4468
rect 22143 4437 22155 4440
rect 22097 4431 22155 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 34514 4468 34520 4480
rect 34475 4440 34520 4468
rect 34514 4428 34520 4440
rect 34572 4428 34578 4480
rect 37458 4468 37464 4480
rect 37419 4440 37464 4468
rect 37458 4428 37464 4440
rect 37516 4428 37522 4480
rect 40770 4468 40776 4480
rect 40731 4440 40776 4468
rect 40770 4428 40776 4440
rect 40828 4428 40834 4480
rect 41279 4471 41337 4477
rect 41279 4437 41291 4471
rect 41325 4468 41337 4471
rect 41690 4468 41696 4480
rect 41325 4440 41696 4468
rect 41325 4437 41337 4440
rect 41279 4431 41337 4437
rect 41690 4428 41696 4440
rect 41748 4428 41754 4480
rect 41874 4468 41880 4480
rect 41835 4440 41880 4468
rect 41874 4428 41880 4440
rect 41932 4428 41938 4480
rect 1104 4378 48852 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 48852 4378
rect 1104 4304 48852 4326
rect 22922 4264 22928 4276
rect 22883 4236 22928 4264
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 25406 4264 25412 4276
rect 25367 4236 25412 4264
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 26970 4264 26976 4276
rect 26931 4236 26976 4264
rect 26970 4224 26976 4236
rect 27028 4224 27034 4276
rect 28307 4267 28365 4273
rect 28307 4233 28319 4267
rect 28353 4264 28365 4267
rect 28626 4264 28632 4276
rect 28353 4236 28632 4264
rect 28353 4233 28365 4236
rect 28307 4227 28365 4233
rect 28626 4224 28632 4236
rect 28684 4224 28690 4276
rect 28994 4264 29000 4276
rect 28736 4236 29000 4264
rect 21726 4196 21732 4208
rect 21687 4168 21732 4196
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 23934 4196 23940 4208
rect 23847 4168 23940 4196
rect 23934 4156 23940 4168
rect 23992 4196 23998 4208
rect 25869 4199 25927 4205
rect 25869 4196 25881 4199
rect 23992 4168 25881 4196
rect 23992 4156 23998 4168
rect 25869 4165 25881 4168
rect 25915 4196 25927 4199
rect 26142 4196 26148 4208
rect 25915 4168 26148 4196
rect 25915 4165 25927 4168
rect 25869 4159 25927 4165
rect 26142 4156 26148 4168
rect 26200 4196 26206 4208
rect 28736 4196 28764 4236
rect 28994 4224 29000 4236
rect 29052 4264 29058 4276
rect 29454 4264 29460 4276
rect 29052 4236 29460 4264
rect 29052 4224 29058 4236
rect 29454 4224 29460 4236
rect 29512 4264 29518 4276
rect 30929 4267 30987 4273
rect 30929 4264 30941 4267
rect 29512 4236 30941 4264
rect 29512 4224 29518 4236
rect 30929 4233 30941 4236
rect 30975 4264 30987 4267
rect 31294 4264 31300 4276
rect 30975 4236 31300 4264
rect 30975 4233 30987 4236
rect 30929 4227 30987 4233
rect 31294 4224 31300 4236
rect 31352 4224 31358 4276
rect 32122 4264 32128 4276
rect 32083 4236 32128 4264
rect 32122 4224 32128 4236
rect 32180 4224 32186 4276
rect 33594 4224 33600 4276
rect 33652 4264 33658 4276
rect 34057 4267 34115 4273
rect 34057 4264 34069 4267
rect 33652 4236 34069 4264
rect 33652 4224 33658 4236
rect 34057 4233 34069 4236
rect 34103 4233 34115 4267
rect 34057 4227 34115 4233
rect 35299 4267 35357 4273
rect 35299 4233 35311 4267
rect 35345 4264 35357 4267
rect 37458 4264 37464 4276
rect 35345 4236 37464 4264
rect 35345 4233 35357 4236
rect 35299 4227 35357 4233
rect 37458 4224 37464 4236
rect 37516 4224 37522 4276
rect 38105 4267 38163 4273
rect 37568 4236 38056 4264
rect 26200 4168 28764 4196
rect 28966 4168 30972 4196
rect 26200 4156 26206 4168
rect 26418 4088 26424 4140
rect 26476 4128 26482 4140
rect 28442 4128 28448 4140
rect 26476 4100 28448 4128
rect 26476 4088 26482 4100
rect 28442 4088 28448 4100
rect 28500 4128 28506 4140
rect 28629 4131 28687 4137
rect 28629 4128 28641 4131
rect 28500 4100 28641 4128
rect 28500 4088 28506 4100
rect 28629 4097 28641 4100
rect 28675 4097 28687 4131
rect 28629 4091 28687 4097
rect 21726 4020 21732 4072
rect 21784 4060 21790 4072
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 21784 4032 21925 4060
rect 21784 4020 21790 4032
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22002 4020 22008 4072
rect 22060 4060 22066 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22060 4032 22385 4060
rect 22060 4020 22066 4032
rect 22373 4029 22385 4032
rect 22419 4060 22431 4063
rect 22462 4060 22468 4072
rect 22419 4032 22468 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4060 24363 4063
rect 24394 4060 24400 4072
rect 24351 4032 24400 4060
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 24394 4020 24400 4032
rect 24452 4020 24458 4072
rect 24486 4020 24492 4072
rect 24544 4060 24550 4072
rect 24854 4060 24860 4072
rect 24544 4032 24860 4060
rect 24544 4020 24550 4032
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 28236 4063 28294 4069
rect 28236 4029 28248 4063
rect 28282 4060 28294 4063
rect 28350 4060 28356 4072
rect 28282 4032 28356 4060
rect 28282 4029 28294 4032
rect 28236 4023 28294 4029
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 22649 3995 22707 4001
rect 22649 3961 22661 3995
rect 22695 3992 22707 3995
rect 22830 3992 22836 4004
rect 22695 3964 22836 3992
rect 22695 3961 22707 3964
rect 22649 3955 22707 3961
rect 22830 3952 22836 3964
rect 22888 3952 22894 4004
rect 25130 3992 25136 4004
rect 25091 3964 25136 3992
rect 25130 3952 25136 3964
rect 25188 3952 25194 4004
rect 26050 3992 26056 4004
rect 26011 3964 26056 3992
rect 26050 3952 26056 3964
rect 26108 3952 26114 4004
rect 26142 3952 26148 4004
rect 26200 3992 26206 4004
rect 26697 3995 26755 4001
rect 26200 3964 26245 3992
rect 26200 3952 26206 3964
rect 26697 3961 26709 3995
rect 26743 3992 26755 3995
rect 26878 3992 26884 4004
rect 26743 3964 26884 3992
rect 26743 3961 26755 3964
rect 26697 3955 26755 3961
rect 26878 3952 26884 3964
rect 26936 3952 26942 4004
rect 27154 3952 27160 4004
rect 27212 3992 27218 4004
rect 28966 3992 28994 4168
rect 29638 4128 29644 4140
rect 29599 4100 29644 4128
rect 29638 4088 29644 4100
rect 29696 4088 29702 4140
rect 30944 4128 30972 4168
rect 31018 4156 31024 4208
rect 31076 4196 31082 4208
rect 33686 4196 33692 4208
rect 31076 4168 33692 4196
rect 31076 4156 31082 4168
rect 33686 4156 33692 4168
rect 33744 4156 33750 4208
rect 35710 4196 35716 4208
rect 35671 4168 35716 4196
rect 35710 4156 35716 4168
rect 35768 4196 35774 4208
rect 35989 4199 36047 4205
rect 35989 4196 36001 4199
rect 35768 4168 36001 4196
rect 35768 4156 35774 4168
rect 35989 4165 36001 4168
rect 36035 4196 36047 4199
rect 36354 4196 36360 4208
rect 36035 4168 36360 4196
rect 36035 4165 36047 4168
rect 35989 4159 36047 4165
rect 36354 4156 36360 4168
rect 36412 4196 36418 4208
rect 37568 4196 37596 4236
rect 36412 4168 37596 4196
rect 37737 4199 37795 4205
rect 36412 4156 36418 4168
rect 37737 4165 37749 4199
rect 37783 4196 37795 4199
rect 37918 4196 37924 4208
rect 37783 4168 37924 4196
rect 37783 4165 37795 4168
rect 37737 4159 37795 4165
rect 37918 4156 37924 4168
rect 37976 4156 37982 4208
rect 38028 4196 38056 4236
rect 38105 4233 38117 4267
rect 38151 4264 38163 4267
rect 38286 4264 38292 4276
rect 38151 4236 38292 4264
rect 38151 4233 38163 4236
rect 38105 4227 38163 4233
rect 38286 4224 38292 4236
rect 38344 4264 38350 4276
rect 38473 4267 38531 4273
rect 38473 4264 38485 4267
rect 38344 4236 38485 4264
rect 38344 4224 38350 4236
rect 38473 4233 38485 4236
rect 38519 4233 38531 4267
rect 38473 4227 38531 4233
rect 39482 4224 39488 4276
rect 39540 4264 39546 4276
rect 40037 4267 40095 4273
rect 40037 4264 40049 4267
rect 39540 4236 40049 4264
rect 39540 4224 39546 4236
rect 40037 4233 40049 4236
rect 40083 4233 40095 4267
rect 41598 4264 41604 4276
rect 41559 4236 41604 4264
rect 40037 4227 40095 4233
rect 41598 4224 41604 4236
rect 41656 4224 41662 4276
rect 43257 4267 43315 4273
rect 43257 4233 43269 4267
rect 43303 4264 43315 4267
rect 43438 4264 43444 4276
rect 43303 4236 43444 4264
rect 43303 4233 43315 4236
rect 43257 4227 43315 4233
rect 43438 4224 43444 4236
rect 43496 4264 43502 4276
rect 44361 4267 44419 4273
rect 44361 4264 44373 4267
rect 43496 4236 44373 4264
rect 43496 4224 43502 4236
rect 44361 4233 44373 4236
rect 44407 4233 44419 4267
rect 46198 4264 46204 4276
rect 44361 4227 44419 4233
rect 44979 4236 46204 4264
rect 39669 4199 39727 4205
rect 39669 4196 39681 4199
rect 38028 4168 39681 4196
rect 39669 4165 39681 4168
rect 39715 4196 39727 4199
rect 39758 4196 39764 4208
rect 39715 4168 39764 4196
rect 39715 4165 39727 4168
rect 39669 4159 39727 4165
rect 39758 4156 39764 4168
rect 39816 4156 39822 4208
rect 43990 4196 43996 4208
rect 43903 4168 43996 4196
rect 43990 4156 43996 4168
rect 44048 4196 44054 4208
rect 44979 4196 45007 4236
rect 46198 4224 46204 4236
rect 46256 4224 46262 4276
rect 45370 4196 45376 4208
rect 44048 4168 45007 4196
rect 45331 4168 45376 4196
rect 44048 4156 44054 4168
rect 45370 4156 45376 4168
rect 45428 4156 45434 4208
rect 31481 4131 31539 4137
rect 31481 4128 31493 4131
rect 30944 4100 31493 4128
rect 31481 4097 31493 4100
rect 31527 4128 31539 4131
rect 33045 4131 33103 4137
rect 33045 4128 33057 4131
rect 31527 4100 33057 4128
rect 31527 4097 31539 4100
rect 31481 4091 31539 4097
rect 33045 4097 33057 4100
rect 33091 4097 33103 4131
rect 33045 4091 33103 4097
rect 42610 4088 42616 4140
rect 42668 4128 42674 4140
rect 43441 4131 43499 4137
rect 43441 4128 43453 4131
rect 42668 4100 43453 4128
rect 42668 4088 42674 4100
rect 43441 4097 43453 4100
rect 43487 4128 43499 4131
rect 44729 4131 44787 4137
rect 44729 4128 44741 4131
rect 43487 4100 44741 4128
rect 43487 4097 43499 4100
rect 43441 4091 43499 4097
rect 44729 4097 44741 4100
rect 44775 4097 44787 4131
rect 44729 4091 44787 4097
rect 34701 4063 34759 4069
rect 34701 4029 34713 4063
rect 34747 4060 34759 4063
rect 35228 4063 35286 4069
rect 35228 4060 35240 4063
rect 34747 4032 35240 4060
rect 34747 4029 34759 4032
rect 34701 4023 34759 4029
rect 35228 4029 35240 4032
rect 35274 4060 35286 4063
rect 36078 4060 36084 4072
rect 35274 4032 36084 4060
rect 35274 4029 35286 4032
rect 35228 4023 35286 4029
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 36906 4020 36912 4072
rect 36964 4060 36970 4072
rect 36964 4032 37009 4060
rect 36964 4020 36970 4032
rect 38286 4020 38292 4072
rect 38344 4060 38350 4072
rect 38657 4063 38715 4069
rect 38657 4060 38669 4063
rect 38344 4032 38669 4060
rect 38344 4020 38350 4032
rect 38657 4029 38669 4032
rect 38703 4029 38715 4063
rect 38657 4023 38715 4029
rect 38838 4020 38844 4072
rect 38896 4060 38902 4072
rect 39117 4063 39175 4069
rect 39117 4060 39129 4063
rect 38896 4032 39129 4060
rect 38896 4020 38902 4032
rect 39117 4029 39129 4032
rect 39163 4029 39175 4063
rect 40770 4060 40776 4072
rect 40731 4032 40776 4060
rect 39117 4023 39175 4029
rect 40770 4020 40776 4032
rect 40828 4020 40834 4072
rect 44964 4063 45022 4069
rect 44964 4029 44976 4063
rect 45010 4060 45022 4063
rect 45738 4060 45744 4072
rect 45010 4032 45744 4060
rect 45010 4029 45022 4032
rect 44964 4023 45022 4029
rect 45738 4020 45744 4032
rect 45796 4020 45802 4072
rect 29362 3992 29368 4004
rect 27212 3964 28994 3992
rect 29323 3964 29368 3992
rect 27212 3952 27218 3964
rect 29362 3952 29368 3964
rect 29420 3952 29426 4004
rect 29454 3952 29460 4004
rect 29512 3992 29518 4004
rect 30653 3995 30711 4001
rect 29512 3964 29557 3992
rect 29512 3952 29518 3964
rect 30653 3961 30665 3995
rect 30699 3992 30711 3995
rect 31202 3992 31208 4004
rect 30699 3964 31208 3992
rect 30699 3961 30711 3964
rect 30653 3955 30711 3961
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 31294 3952 31300 4004
rect 31352 3992 31358 4004
rect 32766 3992 32772 4004
rect 31352 3964 31397 3992
rect 32727 3964 32772 3992
rect 31352 3952 31358 3964
rect 32766 3952 32772 3964
rect 32824 3952 32830 4004
rect 32861 3995 32919 4001
rect 32861 3961 32873 3995
rect 32907 3961 32919 3995
rect 36262 3992 36268 4004
rect 36223 3964 36268 3992
rect 32861 3955 32919 3961
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 23382 3924 23388 3936
rect 22612 3896 23388 3924
rect 22612 3884 22618 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 28074 3924 28080 3936
rect 27987 3896 28080 3924
rect 28074 3884 28080 3896
rect 28132 3924 28138 3936
rect 28442 3924 28448 3936
rect 28132 3896 28448 3924
rect 28132 3884 28138 3896
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 32582 3924 32588 3936
rect 32495 3896 32588 3924
rect 32582 3884 32588 3896
rect 32640 3924 32646 3936
rect 32876 3924 32904 3955
rect 36262 3952 36268 3964
rect 36320 3952 36326 4004
rect 36354 3952 36360 4004
rect 36412 3992 36418 4004
rect 39390 3992 39396 4004
rect 36412 3964 36457 3992
rect 39351 3964 39396 3992
rect 36412 3952 36418 3964
rect 39390 3952 39396 3964
rect 39448 3952 39454 4004
rect 41874 3992 41880 4004
rect 41835 3964 41880 3992
rect 41874 3952 41880 3964
rect 41932 3952 41938 4004
rect 41969 3995 42027 4001
rect 41969 3961 41981 3995
rect 42015 3961 42027 3995
rect 42518 3992 42524 4004
rect 42479 3964 42524 3992
rect 41969 3955 42027 3961
rect 32640 3896 32904 3924
rect 40911 3927 40969 3933
rect 32640 3884 32646 3896
rect 40911 3893 40923 3927
rect 40957 3924 40969 3927
rect 41046 3924 41052 3936
rect 40957 3896 41052 3924
rect 40957 3893 40969 3896
rect 40911 3887 40969 3893
rect 41046 3884 41052 3896
rect 41104 3884 41110 3936
rect 41230 3924 41236 3936
rect 41191 3896 41236 3924
rect 41230 3884 41236 3896
rect 41288 3884 41294 3936
rect 41598 3884 41604 3936
rect 41656 3924 41662 3936
rect 41984 3924 42012 3955
rect 42518 3952 42524 3964
rect 42576 3952 42582 4004
rect 43530 3952 43536 4004
rect 43588 3992 43594 4004
rect 43588 3964 43633 3992
rect 43588 3952 43594 3964
rect 43898 3952 43904 4004
rect 43956 3992 43962 4004
rect 45051 3995 45109 4001
rect 45051 3992 45063 3995
rect 43956 3964 45063 3992
rect 43956 3952 43962 3964
rect 45051 3961 45063 3964
rect 45097 3961 45109 3995
rect 45051 3955 45109 3961
rect 42058 3924 42064 3936
rect 41656 3896 42064 3924
rect 41656 3884 41662 3896
rect 42058 3884 42064 3896
rect 42116 3884 42122 3936
rect 42794 3884 42800 3936
rect 42852 3924 42858 3936
rect 42852 3896 42897 3924
rect 42852 3884 42858 3896
rect 1104 3834 48852 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 48852 3834
rect 1104 3760 48852 3782
rect 22922 3680 22928 3732
rect 22980 3720 22986 3732
rect 23109 3723 23167 3729
rect 23109 3720 23121 3723
rect 22980 3692 23121 3720
rect 22980 3680 22986 3692
rect 23109 3689 23121 3692
rect 23155 3689 23167 3723
rect 23109 3683 23167 3689
rect 32263 3723 32321 3729
rect 32263 3689 32275 3723
rect 32309 3720 32321 3723
rect 32766 3720 32772 3732
rect 32309 3692 32772 3720
rect 32309 3689 32321 3692
rect 32263 3683 32321 3689
rect 32766 3680 32772 3692
rect 32824 3680 32830 3732
rect 36262 3680 36268 3732
rect 36320 3720 36326 3732
rect 36449 3723 36507 3729
rect 36449 3720 36461 3723
rect 36320 3692 36461 3720
rect 36320 3680 36326 3692
rect 36449 3689 36461 3692
rect 36495 3720 36507 3723
rect 36771 3723 36829 3729
rect 36771 3720 36783 3723
rect 36495 3692 36783 3720
rect 36495 3689 36507 3692
rect 36449 3683 36507 3689
rect 36771 3689 36783 3692
rect 36817 3689 36829 3723
rect 36771 3683 36829 3689
rect 37826 3680 37832 3732
rect 37884 3720 37890 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 37884 3692 38117 3720
rect 37884 3680 37890 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 22551 3655 22609 3661
rect 22551 3621 22563 3655
rect 22597 3652 22609 3655
rect 23014 3652 23020 3664
rect 22597 3624 23020 3652
rect 22597 3621 22609 3624
rect 22551 3615 22609 3621
rect 23014 3612 23020 3624
rect 23072 3612 23078 3664
rect 24578 3612 24584 3664
rect 24636 3652 24642 3664
rect 26418 3652 26424 3664
rect 24636 3624 26424 3652
rect 24636 3612 24642 3624
rect 26418 3612 26424 3624
rect 26476 3652 26482 3664
rect 26697 3655 26755 3661
rect 26697 3652 26709 3655
rect 26476 3624 26709 3652
rect 26476 3612 26482 3624
rect 26697 3621 26709 3624
rect 26743 3621 26755 3655
rect 26697 3615 26755 3621
rect 28531 3655 28589 3661
rect 28531 3621 28543 3655
rect 28577 3652 28589 3655
rect 28626 3652 28632 3664
rect 28577 3624 28632 3652
rect 28577 3621 28589 3624
rect 28531 3615 28589 3621
rect 28626 3612 28632 3624
rect 28684 3612 28690 3664
rect 30006 3612 30012 3664
rect 30064 3652 30070 3664
rect 33229 3655 33287 3661
rect 33229 3652 33241 3655
rect 30064 3624 33241 3652
rect 30064 3612 30070 3624
rect 33229 3621 33241 3624
rect 33275 3652 33287 3655
rect 33275 3624 33916 3652
rect 33275 3621 33287 3624
rect 33229 3615 33287 3621
rect 21244 3587 21302 3593
rect 21244 3553 21256 3587
rect 21290 3584 21302 3587
rect 21358 3584 21364 3596
rect 21290 3556 21364 3584
rect 21290 3553 21302 3556
rect 21244 3547 21302 3553
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 24670 3584 24676 3596
rect 24631 3556 24676 3584
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 29362 3584 29368 3596
rect 27448 3556 29368 3584
rect 22189 3519 22247 3525
rect 22189 3485 22201 3519
rect 22235 3516 22247 3519
rect 22830 3516 22836 3528
rect 22235 3488 22836 3516
rect 22235 3485 22247 3488
rect 22189 3479 22247 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 24946 3476 24952 3528
rect 25004 3516 25010 3528
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 25004 3488 25145 3516
rect 25004 3476 25010 3488
rect 25133 3485 25145 3488
rect 25179 3516 25191 3519
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 25179 3488 25421 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 26602 3516 26608 3528
rect 26563 3488 26608 3516
rect 25409 3479 25467 3485
rect 26602 3476 26608 3488
rect 26660 3476 26666 3528
rect 26878 3516 26884 3528
rect 26839 3488 26884 3516
rect 26878 3476 26884 3488
rect 26936 3476 26942 3528
rect 21315 3451 21373 3457
rect 21315 3417 21327 3451
rect 21361 3448 21373 3451
rect 27448 3448 27476 3556
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 30282 3544 30288 3596
rect 30340 3584 30346 3596
rect 30377 3587 30435 3593
rect 30377 3584 30389 3587
rect 30340 3556 30389 3584
rect 30340 3544 30346 3556
rect 30377 3553 30389 3556
rect 30423 3553 30435 3587
rect 30834 3584 30840 3596
rect 30795 3556 30840 3584
rect 30377 3547 30435 3553
rect 30834 3544 30840 3556
rect 30892 3544 30898 3596
rect 32030 3584 32036 3596
rect 31991 3556 32036 3584
rect 32030 3544 32036 3556
rect 32088 3544 32094 3596
rect 33410 3584 33416 3596
rect 33371 3556 33416 3584
rect 33410 3544 33416 3556
rect 33468 3544 33474 3596
rect 33888 3593 33916 3624
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 35206 3655 35264 3661
rect 35206 3652 35218 3655
rect 34664 3624 35218 3652
rect 34664 3612 34670 3624
rect 35206 3621 35218 3624
rect 35252 3621 35264 3655
rect 37090 3652 37096 3664
rect 37051 3624 37096 3652
rect 35206 3615 35264 3621
rect 37090 3612 37096 3624
rect 37148 3652 37154 3664
rect 37550 3652 37556 3664
rect 37148 3624 37556 3652
rect 37148 3612 37154 3624
rect 37550 3612 37556 3624
rect 37608 3612 37614 3664
rect 38120 3652 38148 3683
rect 38562 3680 38568 3732
rect 38620 3720 38626 3732
rect 39390 3720 39396 3732
rect 38620 3692 39205 3720
rect 39351 3692 39396 3720
rect 38620 3680 38626 3692
rect 38120 3624 38792 3652
rect 33873 3587 33931 3593
rect 33873 3553 33885 3587
rect 33919 3584 33931 3587
rect 35894 3584 35900 3596
rect 33919 3556 35900 3584
rect 33919 3553 33931 3556
rect 33873 3547 33931 3553
rect 35894 3544 35900 3556
rect 35952 3544 35958 3596
rect 36538 3544 36544 3596
rect 36596 3584 36602 3596
rect 36668 3587 36726 3593
rect 36668 3584 36680 3587
rect 36596 3556 36680 3584
rect 36596 3544 36602 3556
rect 36668 3553 36680 3556
rect 36714 3553 36726 3587
rect 38286 3584 38292 3596
rect 38247 3556 38292 3584
rect 36668 3547 36726 3553
rect 38286 3544 38292 3556
rect 38344 3544 38350 3596
rect 38764 3593 38792 3624
rect 38749 3587 38807 3593
rect 38749 3553 38761 3587
rect 38795 3553 38807 3587
rect 39177 3584 39205 3692
rect 39390 3680 39396 3692
rect 39448 3680 39454 3732
rect 40773 3723 40831 3729
rect 40773 3689 40785 3723
rect 40819 3720 40831 3723
rect 42794 3720 42800 3732
rect 40819 3692 42800 3720
rect 40819 3689 40831 3692
rect 40773 3683 40831 3689
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 43714 3680 43720 3732
rect 43772 3720 43778 3732
rect 44361 3723 44419 3729
rect 44361 3720 44373 3723
rect 43772 3692 44373 3720
rect 43772 3680 43778 3692
rect 44361 3689 44373 3692
rect 44407 3689 44419 3723
rect 44361 3683 44419 3689
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 39942 3652 39948 3664
rect 39632 3624 39948 3652
rect 39632 3612 39638 3624
rect 39942 3612 39948 3624
rect 40000 3652 40006 3664
rect 40174 3655 40232 3661
rect 40174 3652 40186 3655
rect 40000 3624 40186 3652
rect 40000 3612 40006 3624
rect 40174 3621 40186 3624
rect 40220 3621 40232 3655
rect 40174 3615 40232 3621
rect 41601 3655 41659 3661
rect 41601 3621 41613 3655
rect 41647 3652 41659 3655
rect 41782 3652 41788 3664
rect 41647 3624 41788 3652
rect 41647 3621 41659 3624
rect 41601 3615 41659 3621
rect 41782 3612 41788 3624
rect 41840 3612 41846 3664
rect 41877 3655 41935 3661
rect 41877 3621 41889 3655
rect 41923 3652 41935 3655
rect 41966 3652 41972 3664
rect 41923 3624 41972 3652
rect 41923 3621 41935 3624
rect 41877 3615 41935 3621
rect 41966 3612 41972 3624
rect 42024 3612 42030 3664
rect 42518 3612 42524 3664
rect 42576 3652 42582 3664
rect 43533 3655 43591 3661
rect 42576 3624 42794 3652
rect 42576 3612 42582 3624
rect 39853 3587 39911 3593
rect 39853 3584 39865 3587
rect 39177 3556 39865 3584
rect 38749 3547 38807 3553
rect 39853 3553 39865 3556
rect 39899 3584 39911 3587
rect 40034 3584 40040 3596
rect 39899 3556 40040 3584
rect 39899 3553 39911 3556
rect 39853 3547 39911 3553
rect 40034 3544 40040 3556
rect 40092 3544 40098 3596
rect 42429 3587 42487 3593
rect 42429 3553 42441 3587
rect 42475 3584 42487 3587
rect 42610 3584 42616 3596
rect 42475 3556 42616 3584
rect 42475 3553 42487 3556
rect 42429 3547 42487 3553
rect 42610 3544 42616 3556
rect 42668 3544 42674 3596
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3485 28227 3519
rect 30926 3516 30932 3528
rect 30887 3488 30932 3516
rect 28169 3479 28227 3485
rect 21361 3420 27476 3448
rect 21361 3417 21373 3420
rect 21315 3411 21373 3417
rect 28184 3392 28212 3479
rect 30926 3476 30932 3488
rect 30984 3476 30990 3528
rect 34057 3519 34115 3525
rect 34057 3485 34069 3519
rect 34103 3516 34115 3519
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34103 3488 34897 3516
rect 34103 3485 34115 3488
rect 34057 3479 34115 3485
rect 34885 3485 34897 3488
rect 34931 3516 34943 3519
rect 36078 3516 36084 3528
rect 34931 3488 36084 3516
rect 34931 3485 34943 3488
rect 34885 3479 34943 3485
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 39025 3519 39083 3525
rect 39025 3485 39037 3519
rect 39071 3516 39083 3519
rect 39758 3516 39764 3528
rect 39071 3488 39764 3516
rect 39071 3485 39083 3488
rect 39025 3479 39083 3485
rect 39758 3476 39764 3488
rect 39816 3476 39822 3528
rect 42766 3516 42794 3624
rect 43533 3621 43545 3655
rect 43579 3652 43591 3655
rect 43622 3652 43628 3664
rect 43579 3624 43628 3652
rect 43579 3621 43591 3624
rect 43533 3615 43591 3621
rect 43622 3612 43628 3624
rect 43680 3612 43686 3664
rect 43438 3516 43444 3528
rect 42766 3488 43444 3516
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 43990 3448 43996 3460
rect 43951 3420 43996 3448
rect 43990 3408 43996 3420
rect 44048 3408 44054 3460
rect 22002 3380 22008 3392
rect 21963 3352 22008 3380
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 24026 3380 24032 3392
rect 23987 3352 24032 3380
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 25961 3383 26019 3389
rect 25961 3380 25973 3383
rect 24452 3352 25973 3380
rect 24452 3340 24458 3352
rect 25961 3349 25973 3352
rect 26007 3380 26019 3383
rect 26050 3380 26056 3392
rect 26007 3352 26056 3380
rect 26007 3349 26019 3352
rect 25961 3343 26019 3349
rect 26050 3340 26056 3352
rect 26108 3340 26114 3392
rect 27614 3380 27620 3392
rect 27575 3352 27620 3380
rect 27614 3340 27620 3352
rect 27672 3340 27678 3392
rect 28077 3383 28135 3389
rect 28077 3349 28089 3383
rect 28123 3380 28135 3383
rect 28166 3380 28172 3392
rect 28123 3352 28172 3380
rect 28123 3349 28135 3352
rect 28077 3343 28135 3349
rect 28166 3340 28172 3352
rect 28224 3340 28230 3392
rect 29086 3380 29092 3392
rect 29047 3352 29092 3380
rect 29086 3340 29092 3352
rect 29144 3340 29150 3392
rect 34698 3380 34704 3392
rect 34659 3352 34704 3380
rect 34698 3340 34704 3352
rect 34756 3340 34762 3392
rect 35805 3383 35863 3389
rect 35805 3349 35817 3383
rect 35851 3380 35863 3383
rect 35986 3380 35992 3392
rect 35851 3352 35992 3380
rect 35851 3349 35863 3352
rect 35805 3343 35863 3349
rect 35986 3340 35992 3352
rect 36044 3340 36050 3392
rect 36170 3380 36176 3392
rect 36131 3352 36176 3380
rect 36170 3340 36176 3352
rect 36228 3340 36234 3392
rect 1104 3290 48852 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 48852 3290
rect 1104 3216 48852 3238
rect 20947 3179 21005 3185
rect 20947 3145 20959 3179
rect 20993 3176 21005 3179
rect 22554 3176 22560 3188
rect 20993 3148 22560 3176
rect 20993 3145 21005 3148
rect 20947 3139 21005 3145
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 24075 3179 24133 3185
rect 24075 3145 24087 3179
rect 24121 3176 24133 3179
rect 24394 3176 24400 3188
rect 24121 3148 24400 3176
rect 24121 3145 24133 3148
rect 24075 3139 24133 3145
rect 24394 3136 24400 3148
rect 24452 3136 24458 3188
rect 24489 3179 24547 3185
rect 24489 3145 24501 3179
rect 24535 3176 24547 3179
rect 24670 3176 24676 3188
rect 24535 3148 24676 3176
rect 24535 3145 24547 3148
rect 24489 3139 24547 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 26418 3136 26424 3188
rect 26476 3176 26482 3188
rect 26513 3179 26571 3185
rect 26513 3176 26525 3179
rect 26476 3148 26525 3176
rect 26476 3136 26482 3148
rect 26513 3145 26525 3148
rect 26559 3145 26571 3179
rect 26513 3139 26571 3145
rect 26602 3136 26608 3188
rect 26660 3176 26666 3188
rect 26881 3179 26939 3185
rect 26881 3176 26893 3179
rect 26660 3148 26893 3176
rect 26660 3136 26666 3148
rect 26881 3145 26893 3148
rect 26927 3145 26939 3179
rect 29086 3176 29092 3188
rect 29047 3148 29092 3176
rect 26881 3139 26939 3145
rect 29086 3136 29092 3148
rect 29144 3136 29150 3188
rect 29917 3179 29975 3185
rect 29917 3145 29929 3179
rect 29963 3176 29975 3179
rect 30190 3176 30196 3188
rect 29963 3148 30196 3176
rect 29963 3145 29975 3148
rect 29917 3139 29975 3145
rect 30190 3136 30196 3148
rect 30248 3176 30254 3188
rect 30834 3176 30840 3188
rect 30248 3148 30840 3176
rect 30248 3136 30254 3148
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 31665 3179 31723 3185
rect 31665 3145 31677 3179
rect 31711 3176 31723 3179
rect 32030 3176 32036 3188
rect 31711 3148 32036 3176
rect 31711 3145 31723 3148
rect 31665 3139 31723 3145
rect 32030 3136 32036 3148
rect 32088 3176 32094 3188
rect 32125 3179 32183 3185
rect 32125 3176 32137 3179
rect 32088 3148 32137 3176
rect 32088 3136 32094 3148
rect 32125 3145 32137 3148
rect 32171 3145 32183 3179
rect 32125 3139 32183 3145
rect 33686 3136 33692 3188
rect 33744 3176 33750 3188
rect 34241 3179 34299 3185
rect 34241 3176 34253 3179
rect 33744 3148 34253 3176
rect 33744 3136 33750 3148
rect 34241 3145 34253 3148
rect 34287 3176 34299 3179
rect 34606 3176 34612 3188
rect 34287 3148 34612 3176
rect 34287 3145 34299 3148
rect 34241 3139 34299 3145
rect 34606 3136 34612 3148
rect 34664 3136 34670 3188
rect 35805 3179 35863 3185
rect 35805 3145 35817 3179
rect 35851 3176 35863 3179
rect 36538 3176 36544 3188
rect 35851 3148 36544 3176
rect 35851 3145 35863 3148
rect 35805 3139 35863 3145
rect 36538 3136 36544 3148
rect 36596 3136 36602 3188
rect 39577 3179 39635 3185
rect 39577 3145 39589 3179
rect 39623 3176 39635 3179
rect 41230 3176 41236 3188
rect 39623 3148 41236 3176
rect 39623 3145 39635 3148
rect 39577 3139 39635 3145
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 41785 3179 41843 3185
rect 41785 3145 41797 3179
rect 41831 3176 41843 3179
rect 41966 3176 41972 3188
rect 41831 3148 41972 3176
rect 41831 3145 41843 3148
rect 41785 3139 41843 3145
rect 41966 3136 41972 3148
rect 42024 3136 42030 3188
rect 42058 3136 42064 3188
rect 42116 3176 42122 3188
rect 42426 3176 42432 3188
rect 42116 3148 42432 3176
rect 42116 3136 42122 3148
rect 42426 3136 42432 3148
rect 42484 3136 42490 3188
rect 43349 3179 43407 3185
rect 43349 3145 43361 3179
rect 43395 3176 43407 3179
rect 43622 3176 43628 3188
rect 43395 3148 43628 3176
rect 43395 3145 43407 3148
rect 43349 3139 43407 3145
rect 43622 3136 43628 3148
rect 43680 3136 43686 3188
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 22741 3111 22799 3117
rect 22741 3108 22753 3111
rect 20763 3080 22753 3108
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 20891 2981 20919 3080
rect 22741 3077 22753 3080
rect 22787 3077 22799 3111
rect 28353 3111 28411 3117
rect 28353 3108 28365 3111
rect 22741 3071 22799 3077
rect 23446 3080 28365 3108
rect 21358 3040 21364 3052
rect 21271 3012 21364 3040
rect 21358 3000 21364 3012
rect 21416 3040 21422 3052
rect 23446 3040 23474 3080
rect 28353 3077 28365 3080
rect 28399 3077 28411 3111
rect 28353 3071 28411 3077
rect 28442 3068 28448 3120
rect 28500 3108 28506 3120
rect 29411 3111 29469 3117
rect 29411 3108 29423 3111
rect 28500 3080 29423 3108
rect 28500 3068 28506 3080
rect 29411 3077 29423 3080
rect 29457 3077 29469 3111
rect 36078 3108 36084 3120
rect 29411 3071 29469 3077
rect 33106 3080 33732 3108
rect 36039 3080 36084 3108
rect 24946 3040 24952 3052
rect 21416 3012 23474 3040
rect 24907 3012 24952 3040
rect 21416 3000 21422 3012
rect 24946 3000 24952 3012
rect 25004 3000 25010 3052
rect 30745 3043 30803 3049
rect 30745 3009 30757 3043
rect 30791 3040 30803 3043
rect 30926 3040 30932 3052
rect 30791 3012 30932 3040
rect 30791 3009 30803 3012
rect 30745 3003 30803 3009
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 32769 3043 32827 3049
rect 32769 3009 32781 3043
rect 32815 3040 32827 3043
rect 33106 3040 33134 3080
rect 32815 3012 33134 3040
rect 32815 3009 32827 3012
rect 32769 3003 32827 3009
rect 20876 2975 20934 2981
rect 20876 2941 20888 2975
rect 20922 2941 20934 2975
rect 20876 2935 20934 2941
rect 21821 2975 21879 2981
rect 21821 2941 21833 2975
rect 21867 2972 21879 2975
rect 22554 2972 22560 2984
rect 21867 2944 22560 2972
rect 21867 2941 21879 2944
rect 21821 2935 21879 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24026 2981 24032 2984
rect 24004 2975 24032 2981
rect 24004 2972 24016 2975
rect 23939 2944 24016 2972
rect 24004 2941 24016 2944
rect 24084 2972 24090 2984
rect 25038 2972 25044 2984
rect 24084 2944 25044 2972
rect 24004 2935 24032 2941
rect 24026 2932 24032 2935
rect 24084 2932 24090 2944
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 27433 2975 27491 2981
rect 27433 2941 27445 2975
rect 27479 2972 27491 2975
rect 27614 2972 27620 2984
rect 27479 2944 27620 2972
rect 27479 2941 27491 2944
rect 27433 2935 27491 2941
rect 27614 2932 27620 2944
rect 27672 2972 27678 2984
rect 28258 2972 28264 2984
rect 27672 2944 28264 2972
rect 27672 2932 27678 2944
rect 28258 2932 28264 2944
rect 28316 2932 28322 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29308 2975 29366 2981
rect 29308 2972 29320 2975
rect 29144 2944 29320 2972
rect 29144 2932 29150 2944
rect 29308 2941 29320 2944
rect 29354 2941 29366 2975
rect 32784 2972 32812 3003
rect 29308 2935 29366 2941
rect 29426 2944 32812 2972
rect 33137 2975 33195 2981
rect 21729 2907 21787 2913
rect 21729 2873 21741 2907
rect 21775 2904 21787 2907
rect 22183 2907 22241 2913
rect 22183 2904 22195 2907
rect 21775 2876 22195 2904
rect 21775 2873 21787 2876
rect 21729 2867 21787 2873
rect 22183 2873 22195 2876
rect 22229 2904 22241 2907
rect 23106 2904 23112 2916
rect 22229 2876 23112 2904
rect 22229 2873 22241 2876
rect 22183 2867 22241 2873
rect 23106 2864 23112 2876
rect 23164 2904 23170 2916
rect 24762 2904 24768 2916
rect 23164 2876 24768 2904
rect 23164 2864 23170 2876
rect 24762 2864 24768 2876
rect 24820 2904 24826 2916
rect 24857 2907 24915 2913
rect 24857 2904 24869 2907
rect 24820 2876 24869 2904
rect 24820 2864 24826 2876
rect 24857 2873 24869 2876
rect 24903 2904 24915 2907
rect 25311 2907 25369 2913
rect 25311 2904 25323 2907
rect 24903 2876 25323 2904
rect 24903 2873 24915 2876
rect 24857 2867 24915 2873
rect 25311 2873 25323 2876
rect 25357 2904 25369 2907
rect 27341 2907 27399 2913
rect 27341 2904 27353 2907
rect 25357 2876 27353 2904
rect 25357 2873 25369 2876
rect 25311 2867 25369 2873
rect 27341 2873 27353 2876
rect 27387 2904 27399 2907
rect 27795 2907 27853 2913
rect 27795 2904 27807 2907
rect 27387 2876 27807 2904
rect 27387 2873 27399 2876
rect 27341 2867 27399 2873
rect 27795 2873 27807 2876
rect 27841 2873 27853 2907
rect 27795 2867 27853 2873
rect 23382 2836 23388 2848
rect 23343 2808 23388 2836
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 25866 2836 25872 2848
rect 25827 2808 25872 2836
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 27816 2836 27844 2867
rect 28350 2864 28356 2916
rect 28408 2904 28414 2916
rect 28718 2904 28724 2916
rect 28408 2876 28724 2904
rect 28408 2864 28414 2876
rect 28718 2864 28724 2876
rect 28776 2904 28782 2916
rect 29426 2904 29454 2944
rect 33137 2941 33149 2975
rect 33183 2972 33195 2975
rect 33410 2972 33416 2984
rect 33183 2944 33416 2972
rect 33183 2941 33195 2944
rect 33137 2935 33195 2941
rect 33410 2932 33416 2944
rect 33468 2932 33474 2984
rect 33704 2981 33732 3080
rect 36078 3068 36084 3080
rect 36136 3068 36142 3120
rect 39942 3108 39948 3120
rect 39903 3080 39948 3108
rect 39942 3068 39948 3080
rect 40000 3108 40006 3120
rect 40221 3111 40279 3117
rect 40221 3108 40233 3111
rect 40000 3080 40233 3108
rect 40000 3068 40006 3080
rect 40221 3077 40233 3080
rect 40267 3108 40279 3111
rect 44821 3111 44879 3117
rect 44821 3108 44833 3111
rect 40267 3080 40632 3108
rect 40267 3077 40279 3080
rect 40221 3071 40279 3077
rect 38105 3043 38163 3049
rect 38105 3040 38117 3043
rect 37108 3012 38117 3040
rect 33689 2975 33747 2981
rect 33689 2941 33701 2975
rect 33735 2941 33747 2975
rect 33689 2935 33747 2941
rect 34330 2932 34336 2984
rect 34388 2972 34394 2984
rect 34698 2972 34704 2984
rect 34388 2944 34704 2972
rect 34388 2932 34394 2944
rect 34698 2932 34704 2944
rect 34756 2972 34762 2984
rect 37108 2981 37136 3012
rect 38105 3009 38117 3012
rect 38151 3040 38163 3043
rect 38286 3040 38292 3052
rect 38151 3012 38292 3040
rect 38151 3009 38163 3012
rect 38105 3003 38163 3009
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 38657 3043 38715 3049
rect 38657 3009 38669 3043
rect 38703 3040 38715 3043
rect 39390 3040 39396 3052
rect 38703 3012 39396 3040
rect 38703 3009 38715 3012
rect 38657 3003 38715 3009
rect 39390 3000 39396 3012
rect 39448 3000 39454 3052
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 40494 3040 40500 3052
rect 39816 3012 40500 3040
rect 39816 3000 39822 3012
rect 40494 3000 40500 3012
rect 40552 3000 40558 3052
rect 34885 2975 34943 2981
rect 34885 2972 34897 2975
rect 34756 2944 34897 2972
rect 34756 2932 34762 2944
rect 34885 2941 34897 2944
rect 34931 2941 34943 2975
rect 34885 2935 34943 2941
rect 37001 2975 37059 2981
rect 37001 2941 37013 2975
rect 37047 2972 37059 2975
rect 37093 2975 37151 2981
rect 37093 2972 37105 2975
rect 37047 2944 37105 2972
rect 37047 2941 37059 2944
rect 37001 2935 37059 2941
rect 37093 2941 37105 2944
rect 37139 2941 37151 2975
rect 37550 2972 37556 2984
rect 37511 2944 37556 2972
rect 37093 2935 37151 2941
rect 37550 2932 37556 2944
rect 37608 2932 37614 2984
rect 30653 2907 30711 2913
rect 30653 2904 30665 2907
rect 28776 2876 29454 2904
rect 29564 2876 30665 2904
rect 28776 2864 28782 2876
rect 28626 2836 28632 2848
rect 27816 2808 28632 2836
rect 28626 2796 28632 2808
rect 28684 2836 28690 2848
rect 29564 2836 29592 2876
rect 30653 2873 30665 2876
rect 30699 2904 30711 2907
rect 31018 2904 31024 2916
rect 30699 2876 31024 2904
rect 30699 2873 30711 2876
rect 30653 2867 30711 2873
rect 31018 2864 31024 2876
rect 31076 2913 31082 2916
rect 31076 2907 31124 2913
rect 31076 2873 31078 2907
rect 31112 2873 31124 2907
rect 31076 2867 31124 2873
rect 33965 2907 34023 2913
rect 33965 2873 33977 2907
rect 34011 2904 34023 2907
rect 35066 2904 35072 2916
rect 34011 2876 35072 2904
rect 34011 2873 34023 2876
rect 33965 2867 34023 2873
rect 31076 2864 31082 2867
rect 35066 2864 35072 2876
rect 35124 2864 35130 2916
rect 37826 2904 37832 2916
rect 37787 2876 37832 2904
rect 37826 2864 37832 2876
rect 37884 2864 37890 2916
rect 39019 2907 39077 2913
rect 39019 2904 39031 2907
rect 38626 2876 39031 2904
rect 38626 2848 38654 2876
rect 39019 2873 39031 2876
rect 39065 2904 39077 2907
rect 39942 2904 39948 2916
rect 39065 2876 39948 2904
rect 39065 2873 39077 2876
rect 39019 2867 39077 2873
rect 39942 2864 39948 2876
rect 40000 2864 40006 2916
rect 40604 2904 40632 3080
rect 43916 3080 44833 3108
rect 43916 3052 43944 3080
rect 44821 3077 44833 3080
rect 44867 3077 44879 3111
rect 44821 3071 44879 3077
rect 41690 3000 41696 3052
rect 41748 3040 41754 3052
rect 42334 3040 42340 3052
rect 41748 3012 42340 3040
rect 41748 3000 41754 3012
rect 42334 3000 42340 3012
rect 42392 3000 42398 3052
rect 42610 3040 42616 3052
rect 42571 3012 42616 3040
rect 42610 3000 42616 3012
rect 42668 3000 42674 3052
rect 43898 3040 43904 3052
rect 43859 3012 43904 3040
rect 43898 3000 43904 3012
rect 43956 3000 43962 3052
rect 44082 3000 44088 3052
rect 44140 3040 44146 3052
rect 44177 3043 44235 3049
rect 44177 3040 44189 3043
rect 44140 3012 44189 3040
rect 44140 3000 44146 3012
rect 44177 3009 44189 3012
rect 44223 3009 44235 3043
rect 44177 3003 44235 3009
rect 41417 2975 41475 2981
rect 41417 2941 41429 2975
rect 41463 2972 41475 2975
rect 42058 2972 42064 2984
rect 41463 2944 42064 2972
rect 41463 2941 41475 2944
rect 41417 2935 41475 2941
rect 42058 2932 42064 2944
rect 42116 2932 42122 2984
rect 40818 2907 40876 2913
rect 40818 2904 40830 2907
rect 40604 2876 40830 2904
rect 40818 2873 40830 2876
rect 40864 2873 40876 2907
rect 40818 2867 40876 2873
rect 42426 2864 42432 2916
rect 42484 2904 42490 2916
rect 43993 2907 44051 2913
rect 42484 2876 42529 2904
rect 42484 2864 42490 2876
rect 43993 2873 44005 2907
rect 44039 2873 44051 2907
rect 43993 2867 44051 2873
rect 30282 2836 30288 2848
rect 28684 2808 29592 2836
rect 30243 2808 30288 2836
rect 28684 2796 28690 2808
rect 30282 2796 30288 2808
rect 30340 2796 30346 2848
rect 34606 2796 34612 2848
rect 34664 2836 34670 2848
rect 35253 2839 35311 2845
rect 35253 2836 35265 2839
rect 34664 2808 35265 2836
rect 34664 2796 34670 2808
rect 35253 2805 35265 2808
rect 35299 2836 35311 2839
rect 38473 2839 38531 2845
rect 38473 2836 38485 2839
rect 35299 2808 38485 2836
rect 35299 2805 35311 2808
rect 35253 2799 35311 2805
rect 38473 2805 38485 2808
rect 38519 2836 38531 2839
rect 38626 2836 38660 2848
rect 38519 2808 38660 2836
rect 38519 2805 38531 2808
rect 38473 2799 38531 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 43622 2796 43628 2848
rect 43680 2836 43686 2848
rect 44008 2836 44036 2867
rect 43680 2808 44036 2836
rect 43680 2796 43686 2808
rect 1104 2746 48852 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 48852 2746
rect 1104 2672 48852 2694
rect 21450 2592 21456 2644
rect 21508 2632 21514 2644
rect 21637 2635 21695 2641
rect 21637 2632 21649 2635
rect 21508 2604 21649 2632
rect 21508 2592 21514 2604
rect 21637 2601 21649 2604
rect 21683 2632 21695 2635
rect 22830 2632 22836 2644
rect 21683 2604 21864 2632
rect 22791 2604 22836 2632
rect 21683 2601 21695 2604
rect 21637 2595 21695 2601
rect 21836 2505 21864 2604
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 24489 2635 24547 2641
rect 24489 2601 24501 2635
rect 24535 2632 24547 2635
rect 24854 2632 24860 2644
rect 24535 2604 24860 2632
rect 24535 2601 24547 2604
rect 24489 2595 24547 2601
rect 24854 2592 24860 2604
rect 24912 2592 24918 2644
rect 25038 2592 25044 2644
rect 25096 2632 25102 2644
rect 25869 2635 25927 2641
rect 25869 2632 25881 2635
rect 25096 2604 25881 2632
rect 25096 2592 25102 2604
rect 25869 2601 25881 2604
rect 25915 2601 25927 2635
rect 25869 2595 25927 2601
rect 26602 2592 26608 2644
rect 26660 2632 26666 2644
rect 27019 2635 27077 2641
rect 27019 2632 27031 2635
rect 26660 2604 27031 2632
rect 26660 2592 26666 2604
rect 27019 2601 27031 2604
rect 27065 2601 27077 2635
rect 28166 2632 28172 2644
rect 28127 2604 28172 2632
rect 27019 2595 27077 2601
rect 28166 2592 28172 2604
rect 28224 2592 28230 2644
rect 28258 2592 28264 2644
rect 28316 2632 28322 2644
rect 29825 2635 29883 2641
rect 29825 2632 29837 2635
rect 28316 2604 29837 2632
rect 28316 2592 28322 2604
rect 29825 2601 29837 2604
rect 29871 2601 29883 2635
rect 29825 2595 29883 2601
rect 30837 2635 30895 2641
rect 30837 2601 30849 2635
rect 30883 2632 30895 2635
rect 30926 2632 30932 2644
rect 30883 2604 30932 2632
rect 30883 2601 30895 2604
rect 30837 2595 30895 2601
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 31202 2592 31208 2644
rect 31260 2632 31266 2644
rect 31435 2635 31493 2641
rect 31435 2632 31447 2635
rect 31260 2604 31447 2632
rect 31260 2592 31266 2604
rect 31435 2601 31447 2604
rect 31481 2601 31493 2635
rect 31435 2595 31493 2601
rect 32723 2635 32781 2641
rect 32723 2601 32735 2635
rect 32769 2632 32781 2635
rect 36170 2632 36176 2644
rect 32769 2604 36176 2632
rect 32769 2601 32781 2604
rect 32723 2595 32781 2601
rect 36170 2592 36176 2604
rect 36228 2592 36234 2644
rect 36998 2592 37004 2644
rect 37056 2632 37062 2644
rect 37323 2635 37381 2641
rect 37323 2632 37335 2635
rect 37056 2604 37335 2632
rect 37056 2592 37062 2604
rect 37323 2601 37335 2604
rect 37369 2601 37381 2635
rect 37323 2595 37381 2601
rect 37826 2592 37832 2644
rect 37884 2632 37890 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 37884 2604 38025 2632
rect 37884 2592 37890 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 22554 2564 22560 2576
rect 22467 2536 22560 2564
rect 22554 2524 22560 2536
rect 22612 2564 22618 2576
rect 23382 2564 23388 2576
rect 22612 2536 23388 2564
rect 22612 2524 22618 2536
rect 23382 2524 23388 2536
rect 23440 2524 23446 2576
rect 24762 2564 24768 2576
rect 24723 2536 24768 2564
rect 24762 2524 24768 2536
rect 24820 2564 24826 2576
rect 25270 2567 25328 2573
rect 25270 2564 25282 2567
rect 24820 2536 25282 2564
rect 24820 2524 24826 2536
rect 25270 2533 25282 2536
rect 25316 2533 25328 2567
rect 25270 2527 25328 2533
rect 27617 2567 27675 2573
rect 27617 2533 27629 2567
rect 27663 2564 27675 2567
rect 29181 2567 29239 2573
rect 29181 2564 29193 2567
rect 27663 2536 29193 2564
rect 27663 2533 27675 2536
rect 27617 2527 27675 2533
rect 21821 2499 21879 2505
rect 21821 2465 21833 2499
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 24949 2499 25007 2505
rect 24949 2465 24961 2499
rect 24995 2496 25007 2499
rect 25130 2496 25136 2508
rect 24995 2468 25136 2496
rect 24995 2465 25007 2468
rect 24949 2459 25007 2465
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 22002 2428 22008 2440
rect 21039 2400 22008 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 22002 2388 22008 2400
rect 22060 2428 22066 2440
rect 22296 2428 22324 2459
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 25866 2456 25872 2508
rect 25924 2496 25930 2508
rect 26605 2499 26663 2505
rect 26605 2496 26617 2499
rect 25924 2468 26617 2496
rect 25924 2456 25930 2468
rect 26605 2465 26617 2468
rect 26651 2496 26663 2499
rect 26916 2499 26974 2505
rect 26916 2496 26928 2499
rect 26651 2468 26928 2496
rect 26651 2465 26663 2468
rect 26605 2459 26663 2465
rect 26916 2465 26928 2468
rect 26962 2465 26974 2499
rect 26916 2459 26974 2465
rect 27985 2499 28043 2505
rect 27985 2465 27997 2499
rect 28031 2496 28043 2499
rect 28350 2496 28356 2508
rect 28031 2468 28356 2496
rect 28031 2465 28043 2468
rect 27985 2459 28043 2465
rect 28350 2456 28356 2468
rect 28408 2456 28414 2508
rect 28644 2505 28672 2536
rect 29181 2533 29193 2536
rect 29227 2564 29239 2567
rect 34330 2564 34336 2576
rect 29227 2536 30236 2564
rect 34291 2536 34336 2564
rect 29227 2533 29239 2536
rect 29181 2527 29239 2533
rect 30208 2508 30236 2536
rect 34330 2524 34336 2536
rect 34388 2524 34394 2576
rect 34606 2524 34612 2576
rect 34664 2564 34670 2576
rect 35161 2567 35219 2573
rect 35161 2564 35173 2567
rect 34664 2536 35173 2564
rect 34664 2524 34670 2536
rect 35161 2533 35173 2536
rect 35207 2564 35219 2567
rect 35758 2567 35816 2573
rect 35758 2564 35770 2567
rect 35207 2536 35770 2564
rect 35207 2533 35219 2536
rect 35161 2527 35219 2533
rect 35758 2533 35770 2536
rect 35804 2533 35816 2567
rect 35758 2527 35816 2533
rect 35986 2524 35992 2576
rect 36044 2564 36050 2576
rect 37645 2567 37703 2573
rect 37645 2564 37657 2567
rect 36044 2536 37657 2564
rect 36044 2524 36050 2536
rect 28629 2499 28687 2505
rect 28629 2465 28641 2499
rect 28675 2465 28687 2499
rect 28629 2459 28687 2465
rect 29549 2499 29607 2505
rect 29549 2465 29561 2499
rect 29595 2496 29607 2499
rect 30006 2496 30012 2508
rect 29595 2468 30012 2496
rect 29595 2465 29607 2468
rect 29549 2459 29607 2465
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 30190 2496 30196 2508
rect 30151 2468 30196 2496
rect 30190 2456 30196 2468
rect 30248 2456 30254 2508
rect 31205 2499 31263 2505
rect 31205 2465 31217 2499
rect 31251 2496 31263 2499
rect 31364 2499 31422 2505
rect 31364 2496 31376 2499
rect 31251 2468 31376 2496
rect 31251 2465 31263 2468
rect 31205 2459 31263 2465
rect 31364 2465 31376 2468
rect 31410 2496 31422 2499
rect 31938 2496 31944 2508
rect 31410 2468 31944 2496
rect 31410 2465 31422 2468
rect 31364 2459 31422 2465
rect 31938 2456 31944 2468
rect 31996 2456 32002 2508
rect 32033 2499 32091 2505
rect 32033 2465 32045 2499
rect 32079 2496 32091 2499
rect 32620 2499 32678 2505
rect 32620 2496 32632 2499
rect 32079 2468 32632 2496
rect 32079 2465 32091 2468
rect 32033 2459 32091 2465
rect 32620 2465 32632 2468
rect 32666 2496 32678 2499
rect 33321 2499 33379 2505
rect 32666 2468 33134 2496
rect 32666 2465 32678 2468
rect 32620 2459 32678 2465
rect 22060 2400 22324 2428
rect 25148 2428 25176 2456
rect 26145 2431 26203 2437
rect 26145 2428 26157 2431
rect 25148 2400 26157 2428
rect 22060 2388 22066 2400
rect 26145 2397 26157 2400
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 33106 2360 33134 2468
rect 33321 2465 33333 2499
rect 33367 2496 33379 2499
rect 33410 2496 33416 2508
rect 33367 2468 33416 2496
rect 33367 2465 33379 2468
rect 33321 2459 33379 2465
rect 33410 2456 33416 2468
rect 33468 2496 33474 2508
rect 33873 2499 33931 2505
rect 33873 2496 33885 2499
rect 33468 2468 33885 2496
rect 33468 2456 33474 2468
rect 33873 2465 33885 2468
rect 33919 2465 33931 2499
rect 33873 2459 33931 2465
rect 34149 2499 34207 2505
rect 34149 2465 34161 2499
rect 34195 2496 34207 2499
rect 34422 2496 34428 2508
rect 34195 2468 34428 2496
rect 34195 2465 34207 2468
rect 34149 2459 34207 2465
rect 33888 2428 33916 2459
rect 34422 2456 34428 2468
rect 34480 2456 34486 2508
rect 35066 2456 35072 2508
rect 35124 2496 35130 2508
rect 37235 2505 37263 2536
rect 37645 2533 37657 2536
rect 37691 2533 37703 2567
rect 37645 2527 37703 2533
rect 35437 2499 35495 2505
rect 35437 2496 35449 2499
rect 35124 2468 35449 2496
rect 35124 2456 35130 2468
rect 35437 2465 35449 2468
rect 35483 2496 35495 2499
rect 36633 2499 36691 2505
rect 36633 2496 36645 2499
rect 35483 2468 36645 2496
rect 35483 2465 35495 2468
rect 35437 2459 35495 2465
rect 36633 2465 36645 2468
rect 36679 2465 36691 2499
rect 37220 2499 37278 2505
rect 37220 2496 37232 2499
rect 37198 2468 37232 2496
rect 36633 2459 36691 2465
rect 37220 2465 37232 2468
rect 37266 2465 37278 2499
rect 38028 2496 38056 2595
rect 38654 2592 38660 2644
rect 38712 2632 38718 2644
rect 40034 2632 40040 2644
rect 38712 2604 38757 2632
rect 39995 2604 40040 2632
rect 38712 2592 38718 2604
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 40494 2632 40500 2644
rect 40455 2604 40500 2632
rect 40494 2592 40500 2604
rect 40552 2592 40558 2644
rect 40957 2635 41015 2641
rect 40957 2601 40969 2635
rect 41003 2632 41015 2635
rect 41046 2632 41052 2644
rect 41003 2604 41052 2632
rect 41003 2601 41015 2604
rect 40957 2595 41015 2601
rect 41046 2592 41052 2604
rect 41104 2592 41110 2644
rect 41601 2635 41659 2641
rect 41601 2601 41613 2635
rect 41647 2632 41659 2635
rect 41647 2604 41920 2632
rect 41647 2601 41659 2604
rect 41601 2595 41659 2601
rect 38672 2564 38700 2592
rect 39162 2567 39220 2573
rect 39162 2564 39174 2567
rect 38672 2536 39174 2564
rect 39162 2533 39174 2536
rect 39208 2533 39220 2567
rect 41064 2564 41092 2592
rect 41892 2573 41920 2604
rect 41785 2567 41843 2573
rect 41785 2564 41797 2567
rect 41064 2536 41797 2564
rect 39162 2527 39220 2533
rect 41785 2533 41797 2536
rect 41831 2533 41843 2567
rect 41785 2527 41843 2533
rect 41877 2567 41935 2573
rect 41877 2533 41889 2567
rect 41923 2564 41935 2567
rect 41966 2564 41972 2576
rect 41923 2536 41972 2564
rect 41923 2533 41935 2536
rect 41877 2527 41935 2533
rect 41966 2524 41972 2536
rect 42024 2524 42030 2576
rect 42429 2567 42487 2573
rect 42429 2533 42441 2567
rect 42475 2564 42487 2567
rect 43349 2567 43407 2573
rect 43349 2564 43361 2567
rect 42475 2536 43361 2564
rect 42475 2533 42487 2536
rect 42429 2527 42487 2533
rect 43349 2533 43361 2536
rect 43395 2564 43407 2567
rect 43438 2564 43444 2576
rect 43395 2536 43444 2564
rect 43395 2533 43407 2536
rect 43349 2527 43407 2533
rect 43438 2524 43444 2536
rect 43496 2524 43502 2576
rect 38841 2499 38899 2505
rect 38841 2496 38853 2499
rect 38028 2468 38853 2496
rect 37220 2459 37278 2465
rect 38841 2465 38853 2468
rect 38887 2465 38899 2499
rect 38841 2459 38899 2465
rect 39761 2499 39819 2505
rect 39761 2465 39773 2499
rect 39807 2496 39819 2499
rect 40770 2496 40776 2508
rect 39807 2468 40776 2496
rect 39807 2465 39819 2468
rect 39761 2459 39819 2465
rect 40770 2456 40776 2468
rect 40828 2456 40834 2508
rect 44028 2499 44086 2505
rect 44028 2496 44040 2499
rect 42766 2468 44040 2496
rect 34609 2431 34667 2437
rect 34609 2428 34621 2431
rect 33888 2400 34621 2428
rect 34609 2397 34621 2400
rect 34655 2397 34667 2431
rect 34609 2391 34667 2397
rect 42058 2388 42064 2440
rect 42116 2428 42122 2440
rect 42766 2428 42794 2468
rect 44028 2465 44040 2468
rect 44074 2496 44086 2499
rect 44453 2499 44511 2505
rect 44453 2496 44465 2499
rect 44074 2468 44465 2496
rect 44074 2465 44086 2468
rect 44028 2459 44086 2465
rect 44453 2465 44465 2468
rect 44499 2465 44511 2499
rect 44453 2459 44511 2465
rect 42116 2400 42794 2428
rect 42116 2388 42122 2400
rect 36357 2363 36415 2369
rect 36357 2360 36369 2363
rect 33106 2332 36369 2360
rect 36357 2329 36369 2332
rect 36403 2329 36415 2363
rect 36357 2323 36415 2329
rect 41874 2320 41880 2372
rect 41932 2360 41938 2372
rect 44131 2363 44189 2369
rect 44131 2360 44143 2363
rect 41932 2332 44143 2360
rect 41932 2320 41938 2332
rect 44131 2329 44143 2332
rect 44177 2329 44189 2363
rect 44131 2323 44189 2329
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 32401 2295 32459 2301
rect 32401 2292 32413 2295
rect 30340 2264 32413 2292
rect 30340 2252 30346 2264
rect 32401 2261 32413 2264
rect 32447 2292 32459 2295
rect 34422 2292 34428 2304
rect 32447 2264 34428 2292
rect 32447 2261 32459 2264
rect 32401 2255 32459 2261
rect 34422 2252 34428 2264
rect 34480 2252 34486 2304
rect 42334 2252 42340 2304
rect 42392 2292 42398 2304
rect 42705 2295 42763 2301
rect 42705 2292 42717 2295
rect 42392 2264 42717 2292
rect 42392 2252 42398 2264
rect 42705 2261 42717 2264
rect 42751 2261 42763 2295
rect 42705 2255 42763 2261
rect 1104 2202 48852 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 41052 47107 41104 47116
rect 41052 47073 41061 47107
rect 41061 47073 41095 47107
rect 41095 47073 41104 47107
rect 41052 47064 41104 47073
rect 41512 46860 41564 46912
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 36084 46588 36136 46640
rect 41052 46588 41104 46640
rect 41512 46563 41564 46572
rect 41512 46529 41521 46563
rect 41521 46529 41555 46563
rect 41555 46529 41564 46563
rect 41512 46520 41564 46529
rect 36268 46452 36320 46504
rect 41696 46384 41748 46436
rect 42340 46384 42392 46436
rect 28172 46316 28224 46368
rect 28448 46359 28500 46368
rect 28448 46325 28457 46359
rect 28457 46325 28491 46359
rect 28491 46325 28500 46359
rect 28448 46316 28500 46325
rect 34704 46316 34756 46368
rect 36360 46316 36412 46368
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 30196 46155 30248 46164
rect 30196 46121 30205 46155
rect 30205 46121 30239 46155
rect 30239 46121 30248 46155
rect 30196 46112 30248 46121
rect 36360 46112 36412 46164
rect 28724 46044 28776 46096
rect 34152 46044 34204 46096
rect 43720 46112 43772 46164
rect 41604 46044 41656 46096
rect 30380 46019 30432 46028
rect 30380 45985 30389 46019
rect 30389 45985 30423 46019
rect 30423 45985 30432 46019
rect 30380 45976 30432 45985
rect 31208 45976 31260 46028
rect 35624 45976 35676 46028
rect 36544 45976 36596 46028
rect 39856 46019 39908 46028
rect 39856 45985 39865 46019
rect 39865 45985 39899 46019
rect 39899 45985 39908 46019
rect 39856 45976 39908 45985
rect 28632 45908 28684 45960
rect 29000 45951 29052 45960
rect 29000 45917 29009 45951
rect 29009 45917 29043 45951
rect 29043 45917 29052 45951
rect 29000 45908 29052 45917
rect 25320 45815 25372 45824
rect 25320 45781 25329 45815
rect 25329 45781 25363 45815
rect 25363 45781 25372 45815
rect 25320 45772 25372 45781
rect 32864 45815 32916 45824
rect 32864 45781 32873 45815
rect 32873 45781 32907 45815
rect 32907 45781 32916 45815
rect 32864 45772 32916 45781
rect 33324 45772 33376 45824
rect 36084 45908 36136 45960
rect 41788 45951 41840 45960
rect 41788 45917 41797 45951
rect 41797 45917 41831 45951
rect 41831 45917 41840 45951
rect 41788 45908 41840 45917
rect 38108 45840 38160 45892
rect 42340 45883 42392 45892
rect 42340 45849 42349 45883
rect 42349 45849 42383 45883
rect 42383 45849 42392 45883
rect 42340 45840 42392 45849
rect 36452 45772 36504 45824
rect 40592 45772 40644 45824
rect 40684 45772 40736 45824
rect 41696 45772 41748 45824
rect 42156 45772 42208 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 18880 45568 18932 45620
rect 21548 45568 21600 45620
rect 28632 45611 28684 45620
rect 28632 45577 28641 45611
rect 28641 45577 28675 45611
rect 28675 45577 28684 45611
rect 28632 45568 28684 45577
rect 28724 45568 28776 45620
rect 28724 45432 28776 45484
rect 25320 45339 25372 45348
rect 25320 45305 25329 45339
rect 25329 45305 25363 45339
rect 25363 45305 25372 45339
rect 25320 45296 25372 45305
rect 25412 45339 25464 45348
rect 25412 45305 25421 45339
rect 25421 45305 25455 45339
rect 25455 45305 25464 45339
rect 25412 45296 25464 45305
rect 27712 45339 27764 45348
rect 27712 45305 27721 45339
rect 27721 45305 27755 45339
rect 27755 45305 27764 45339
rect 27712 45296 27764 45305
rect 30380 45568 30432 45620
rect 34704 45611 34756 45620
rect 34704 45577 34713 45611
rect 34713 45577 34747 45611
rect 34747 45577 34756 45611
rect 34704 45568 34756 45577
rect 29368 45432 29420 45484
rect 30196 45432 30248 45484
rect 36268 45568 36320 45620
rect 39856 45611 39908 45620
rect 39856 45577 39865 45611
rect 39865 45577 39899 45611
rect 39899 45577 39908 45611
rect 39856 45568 39908 45577
rect 42156 45611 42208 45620
rect 42156 45577 42165 45611
rect 42165 45577 42199 45611
rect 42199 45577 42208 45611
rect 42156 45568 42208 45577
rect 42524 45568 42576 45620
rect 36360 45432 36412 45484
rect 41788 45500 41840 45552
rect 36820 45475 36872 45484
rect 36820 45441 36829 45475
rect 36829 45441 36863 45475
rect 36863 45441 36872 45475
rect 36820 45432 36872 45441
rect 38108 45475 38160 45484
rect 38108 45441 38117 45475
rect 38117 45441 38151 45475
rect 38151 45441 38160 45475
rect 38108 45432 38160 45441
rect 38384 45475 38436 45484
rect 38384 45441 38393 45475
rect 38393 45441 38427 45475
rect 38427 45441 38436 45475
rect 38384 45432 38436 45441
rect 40592 45475 40644 45484
rect 40592 45441 40601 45475
rect 40601 45441 40635 45475
rect 40635 45441 40644 45475
rect 40592 45432 40644 45441
rect 42432 45475 42484 45484
rect 42432 45441 42441 45475
rect 42441 45441 42475 45475
rect 42475 45441 42484 45475
rect 42432 45432 42484 45441
rect 32864 45364 32916 45416
rect 25136 45271 25188 45280
rect 25136 45237 25145 45271
rect 25145 45237 25179 45271
rect 25179 45237 25188 45271
rect 25136 45228 25188 45237
rect 27620 45228 27672 45280
rect 30196 45296 30248 45348
rect 34152 45339 34204 45348
rect 31208 45228 31260 45280
rect 31300 45228 31352 45280
rect 32220 45228 32272 45280
rect 34152 45305 34161 45339
rect 34161 45305 34195 45339
rect 34195 45305 34204 45339
rect 34152 45296 34204 45305
rect 35256 45296 35308 45348
rect 40684 45339 40736 45348
rect 33416 45228 33468 45280
rect 36084 45271 36136 45280
rect 36084 45237 36093 45271
rect 36093 45237 36127 45271
rect 36127 45237 36136 45271
rect 36084 45228 36136 45237
rect 36452 45228 36504 45280
rect 40684 45305 40693 45339
rect 40693 45305 40727 45339
rect 40727 45305 40736 45339
rect 40684 45296 40736 45305
rect 41512 45296 41564 45348
rect 42524 45339 42576 45348
rect 39580 45228 39632 45280
rect 41604 45228 41656 45280
rect 42524 45305 42533 45339
rect 42533 45305 42567 45339
rect 42567 45305 42576 45339
rect 42524 45296 42576 45305
rect 43720 45296 43772 45348
rect 43812 45228 43864 45280
rect 44824 45228 44876 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 27620 45067 27672 45076
rect 27620 45033 27629 45067
rect 27629 45033 27663 45067
rect 27663 45033 27672 45067
rect 27620 45024 27672 45033
rect 29368 45067 29420 45076
rect 29368 45033 29377 45067
rect 29377 45033 29411 45067
rect 29411 45033 29420 45067
rect 29368 45024 29420 45033
rect 30380 45024 30432 45076
rect 25136 44956 25188 45008
rect 25412 44956 25464 45008
rect 28172 44956 28224 45008
rect 28448 44999 28500 45008
rect 28448 44965 28457 44999
rect 28457 44965 28491 44999
rect 28491 44965 28500 44999
rect 29000 44999 29052 45008
rect 28448 44956 28500 44965
rect 29000 44965 29009 44999
rect 29009 44965 29043 44999
rect 29043 44965 29052 44999
rect 29000 44956 29052 44965
rect 32220 45024 32272 45076
rect 36084 45024 36136 45076
rect 32864 44999 32916 45008
rect 32864 44965 32873 44999
rect 32873 44965 32907 44999
rect 32907 44965 32916 44999
rect 32864 44956 32916 44965
rect 34152 44999 34204 45008
rect 34152 44965 34161 44999
rect 34161 44965 34195 44999
rect 34195 44965 34204 44999
rect 34152 44956 34204 44965
rect 34796 44956 34848 45008
rect 38384 45024 38436 45076
rect 40592 45067 40644 45076
rect 40592 45033 40601 45067
rect 40601 45033 40635 45067
rect 40635 45033 40644 45067
rect 40592 45024 40644 45033
rect 42432 45067 42484 45076
rect 42432 45033 42441 45067
rect 42441 45033 42475 45067
rect 42475 45033 42484 45067
rect 42432 45024 42484 45033
rect 36452 44956 36504 45008
rect 36544 44956 36596 45008
rect 39948 44956 40000 45008
rect 40224 44956 40276 45008
rect 41604 44956 41656 45008
rect 43812 44956 43864 45008
rect 23848 44931 23900 44940
rect 23848 44897 23857 44931
rect 23857 44897 23891 44931
rect 23891 44897 23900 44931
rect 23848 44888 23900 44897
rect 27068 44888 27120 44940
rect 30380 44931 30432 44940
rect 30380 44897 30389 44931
rect 30389 44897 30423 44931
rect 30423 44897 30432 44931
rect 30380 44888 30432 44897
rect 31208 44888 31260 44940
rect 32128 44931 32180 44940
rect 32128 44897 32137 44931
rect 32137 44897 32171 44931
rect 32171 44897 32180 44931
rect 32128 44888 32180 44897
rect 32220 44888 32272 44940
rect 37740 44888 37792 44940
rect 24952 44863 25004 44872
rect 24952 44829 24961 44863
rect 24961 44829 24995 44863
rect 24995 44829 25004 44863
rect 24952 44820 25004 44829
rect 25872 44820 25924 44872
rect 27804 44820 27856 44872
rect 30748 44820 30800 44872
rect 34060 44863 34112 44872
rect 34060 44829 34069 44863
rect 34069 44829 34103 44863
rect 34103 44829 34112 44863
rect 34060 44820 34112 44829
rect 36176 44863 36228 44872
rect 36176 44829 36185 44863
rect 36185 44829 36219 44863
rect 36219 44829 36228 44863
rect 36176 44820 36228 44829
rect 39304 44863 39356 44872
rect 39304 44829 39313 44863
rect 39313 44829 39347 44863
rect 39347 44829 39356 44863
rect 39304 44820 39356 44829
rect 41512 44863 41564 44872
rect 35256 44752 35308 44804
rect 41512 44829 41521 44863
rect 41521 44829 41555 44863
rect 41555 44829 41564 44863
rect 41512 44820 41564 44829
rect 43444 44863 43496 44872
rect 43444 44829 43453 44863
rect 43453 44829 43487 44863
rect 43487 44829 43496 44863
rect 43444 44820 43496 44829
rect 43720 44863 43772 44872
rect 43720 44829 43729 44863
rect 43729 44829 43763 44863
rect 43763 44829 43772 44863
rect 43720 44820 43772 44829
rect 41328 44752 41380 44804
rect 27436 44684 27488 44736
rect 31392 44727 31444 44736
rect 31392 44693 31401 44727
rect 31401 44693 31435 44727
rect 31435 44693 31444 44727
rect 31392 44684 31444 44693
rect 35348 44727 35400 44736
rect 35348 44693 35357 44727
rect 35357 44693 35391 44727
rect 35391 44693 35400 44727
rect 35348 44684 35400 44693
rect 38568 44684 38620 44736
rect 40224 44727 40276 44736
rect 40224 44693 40233 44727
rect 40233 44693 40267 44727
rect 40267 44693 40276 44727
rect 40224 44684 40276 44693
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 22284 44523 22336 44532
rect 22284 44489 22293 44523
rect 22293 44489 22327 44523
rect 22327 44489 22336 44523
rect 22284 44480 22336 44489
rect 24952 44480 25004 44532
rect 28172 44480 28224 44532
rect 30380 44480 30432 44532
rect 32220 44523 32272 44532
rect 32220 44489 32229 44523
rect 32229 44489 32263 44523
rect 32263 44489 32272 44523
rect 32220 44480 32272 44489
rect 33324 44480 33376 44532
rect 34060 44480 34112 44532
rect 39580 44523 39632 44532
rect 39580 44489 39589 44523
rect 39589 44489 39623 44523
rect 39623 44489 39632 44523
rect 39580 44480 39632 44489
rect 40224 44523 40276 44532
rect 40224 44489 40233 44523
rect 40233 44489 40267 44523
rect 40267 44489 40276 44523
rect 40224 44480 40276 44489
rect 41788 44480 41840 44532
rect 42156 44480 42208 44532
rect 27712 44412 27764 44464
rect 21548 44344 21600 44396
rect 25688 44387 25740 44396
rect 19156 44276 19208 44328
rect 22284 44276 22336 44328
rect 25688 44353 25697 44387
rect 25697 44353 25731 44387
rect 25731 44353 25740 44387
rect 25688 44344 25740 44353
rect 27436 44387 27488 44396
rect 27436 44353 27445 44387
rect 27445 44353 27479 44387
rect 27479 44353 27488 44387
rect 27436 44344 27488 44353
rect 27804 44387 27856 44396
rect 27804 44353 27813 44387
rect 27813 44353 27847 44387
rect 27847 44353 27856 44387
rect 27804 44344 27856 44353
rect 30840 44344 30892 44396
rect 31392 44344 31444 44396
rect 32956 44319 33008 44328
rect 32956 44285 32965 44319
rect 32965 44285 32999 44319
rect 32999 44285 33008 44319
rect 32956 44276 33008 44285
rect 35348 44344 35400 44396
rect 35992 44344 36044 44396
rect 21364 44208 21416 44260
rect 23848 44251 23900 44260
rect 23848 44217 23857 44251
rect 23857 44217 23891 44251
rect 23891 44217 23900 44251
rect 23848 44208 23900 44217
rect 25228 44251 25280 44260
rect 25228 44217 25237 44251
rect 25237 44217 25271 44251
rect 25271 44217 25280 44251
rect 25228 44208 25280 44217
rect 19248 44183 19300 44192
rect 19248 44149 19257 44183
rect 19257 44149 19291 44183
rect 19291 44149 19300 44183
rect 19248 44140 19300 44149
rect 22008 44140 22060 44192
rect 25412 44208 25464 44260
rect 27620 44208 27672 44260
rect 30196 44208 30248 44260
rect 35256 44208 35308 44260
rect 36544 44251 36596 44260
rect 36544 44217 36553 44251
rect 36553 44217 36587 44251
rect 36587 44217 36596 44251
rect 36544 44208 36596 44217
rect 39948 44455 40000 44464
rect 37832 44387 37884 44396
rect 37832 44353 37841 44387
rect 37841 44353 37875 44387
rect 37875 44353 37884 44387
rect 37832 44344 37884 44353
rect 38568 44276 38620 44328
rect 39948 44421 39957 44455
rect 39957 44421 39991 44455
rect 39991 44421 40000 44455
rect 39948 44412 40000 44421
rect 49516 44412 49568 44464
rect 42708 44344 42760 44396
rect 43812 44344 43864 44396
rect 27068 44183 27120 44192
rect 27068 44149 27077 44183
rect 27077 44149 27111 44183
rect 27111 44149 27120 44183
rect 27068 44140 27120 44149
rect 27160 44140 27212 44192
rect 28448 44183 28500 44192
rect 28448 44149 28457 44183
rect 28457 44149 28491 44183
rect 28491 44149 28500 44183
rect 28448 44140 28500 44149
rect 36452 44140 36504 44192
rect 37832 44140 37884 44192
rect 41328 44183 41380 44192
rect 41328 44149 41337 44183
rect 41337 44149 41371 44183
rect 41371 44149 41380 44183
rect 41328 44140 41380 44149
rect 43720 44276 43772 44328
rect 44272 44276 44324 44328
rect 43444 44208 43496 44260
rect 42156 44140 42208 44192
rect 43628 44140 43680 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 25320 43936 25372 43988
rect 25412 43979 25464 43988
rect 25412 43945 25421 43979
rect 25421 43945 25455 43979
rect 25455 43945 25464 43979
rect 25412 43936 25464 43945
rect 27160 43936 27212 43988
rect 27436 43936 27488 43988
rect 19340 43868 19392 43920
rect 22100 43868 22152 43920
rect 25228 43868 25280 43920
rect 31300 43936 31352 43988
rect 32128 43936 32180 43988
rect 33416 43979 33468 43988
rect 28448 43911 28500 43920
rect 24768 43800 24820 43852
rect 25320 43800 25372 43852
rect 28448 43877 28457 43911
rect 28457 43877 28491 43911
rect 28491 43877 28500 43911
rect 28448 43868 28500 43877
rect 29000 43911 29052 43920
rect 29000 43877 29009 43911
rect 29009 43877 29043 43911
rect 29043 43877 29052 43911
rect 29000 43868 29052 43877
rect 30196 43868 30248 43920
rect 26792 43800 26844 43852
rect 27436 43843 27488 43852
rect 27436 43809 27445 43843
rect 27445 43809 27479 43843
rect 27479 43809 27488 43843
rect 27436 43800 27488 43809
rect 27620 43800 27672 43852
rect 30748 43800 30800 43852
rect 19156 43775 19208 43784
rect 19156 43741 19165 43775
rect 19165 43741 19199 43775
rect 19199 43741 19208 43775
rect 19156 43732 19208 43741
rect 21916 43775 21968 43784
rect 21916 43741 21925 43775
rect 21925 43741 21959 43775
rect 21959 43741 21968 43775
rect 21916 43732 21968 43741
rect 18052 43664 18104 43716
rect 23388 43732 23440 43784
rect 28356 43775 28408 43784
rect 28356 43741 28365 43775
rect 28365 43741 28399 43775
rect 28399 43741 28408 43775
rect 28356 43732 28408 43741
rect 33416 43945 33425 43979
rect 33425 43945 33459 43979
rect 33459 43945 33468 43979
rect 33416 43936 33468 43945
rect 35348 43936 35400 43988
rect 36176 43936 36228 43988
rect 41328 43936 41380 43988
rect 42708 43979 42760 43988
rect 42708 43945 42717 43979
rect 42717 43945 42751 43979
rect 42751 43945 42760 43979
rect 42708 43936 42760 43945
rect 35256 43911 35308 43920
rect 35256 43877 35265 43911
rect 35265 43877 35299 43911
rect 35299 43877 35308 43911
rect 35256 43868 35308 43877
rect 39304 43868 39356 43920
rect 43444 43868 43496 43920
rect 43812 43868 43864 43920
rect 44088 43868 44140 43920
rect 34704 43800 34756 43852
rect 36176 43843 36228 43852
rect 36176 43809 36185 43843
rect 36185 43809 36219 43843
rect 36219 43809 36228 43843
rect 36176 43800 36228 43809
rect 36544 43800 36596 43852
rect 38936 43843 38988 43852
rect 33048 43775 33100 43784
rect 33048 43741 33057 43775
rect 33057 43741 33091 43775
rect 33091 43741 33100 43775
rect 33048 43732 33100 43741
rect 38384 43664 38436 43716
rect 38936 43809 38945 43843
rect 38945 43809 38979 43843
rect 38979 43809 38988 43843
rect 38936 43800 38988 43809
rect 41052 43843 41104 43852
rect 41052 43809 41061 43843
rect 41061 43809 41095 43843
rect 41095 43809 41104 43843
rect 41052 43800 41104 43809
rect 42524 43800 42576 43852
rect 41880 43732 41932 43784
rect 43628 43732 43680 43784
rect 43720 43775 43772 43784
rect 43720 43741 43729 43775
rect 43729 43741 43763 43775
rect 43763 43741 43772 43775
rect 43720 43732 43772 43741
rect 42156 43664 42208 43716
rect 42708 43664 42760 43716
rect 16488 43639 16540 43648
rect 16488 43605 16497 43639
rect 16497 43605 16531 43639
rect 16531 43605 16540 43639
rect 16488 43596 16540 43605
rect 26608 43596 26660 43648
rect 30932 43639 30984 43648
rect 30932 43605 30941 43639
rect 30941 43605 30975 43639
rect 30975 43605 30984 43639
rect 30932 43596 30984 43605
rect 31208 43639 31260 43648
rect 31208 43605 31217 43639
rect 31217 43605 31251 43639
rect 31251 43605 31260 43639
rect 31208 43596 31260 43605
rect 34244 43596 34296 43648
rect 36636 43639 36688 43648
rect 36636 43605 36645 43639
rect 36645 43605 36679 43639
rect 36679 43605 36688 43639
rect 36636 43596 36688 43605
rect 41788 43596 41840 43648
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 19156 43392 19208 43444
rect 24768 43435 24820 43444
rect 18052 43324 18104 43376
rect 16488 43299 16540 43308
rect 16488 43265 16497 43299
rect 16497 43265 16531 43299
rect 16531 43265 16540 43299
rect 16488 43256 16540 43265
rect 17224 43256 17276 43308
rect 16580 43163 16632 43172
rect 16580 43129 16589 43163
rect 16589 43129 16623 43163
rect 16623 43129 16632 43163
rect 16580 43120 16632 43129
rect 18972 43120 19024 43172
rect 24768 43401 24777 43435
rect 24777 43401 24811 43435
rect 24811 43401 24820 43435
rect 24768 43392 24820 43401
rect 26608 43435 26660 43444
rect 26608 43401 26617 43435
rect 26617 43401 26651 43435
rect 26651 43401 26660 43435
rect 26608 43392 26660 43401
rect 28356 43392 28408 43444
rect 28632 43435 28684 43444
rect 28632 43401 28641 43435
rect 28641 43401 28675 43435
rect 28675 43401 28684 43435
rect 28632 43392 28684 43401
rect 30748 43435 30800 43444
rect 30748 43401 30757 43435
rect 30757 43401 30791 43435
rect 30791 43401 30800 43435
rect 30748 43392 30800 43401
rect 34244 43435 34296 43444
rect 34244 43401 34253 43435
rect 34253 43401 34287 43435
rect 34287 43401 34296 43435
rect 34244 43392 34296 43401
rect 34704 43435 34756 43444
rect 34704 43401 34713 43435
rect 34713 43401 34747 43435
rect 34747 43401 34756 43435
rect 34704 43392 34756 43401
rect 36176 43392 36228 43444
rect 42156 43392 42208 43444
rect 43628 43392 43680 43444
rect 44088 43435 44140 43444
rect 44088 43401 44097 43435
rect 44097 43401 44131 43435
rect 44131 43401 44140 43435
rect 44088 43392 44140 43401
rect 21916 43324 21968 43376
rect 22376 43256 22428 43308
rect 30380 43324 30432 43376
rect 27620 43299 27672 43308
rect 27620 43265 27629 43299
rect 27629 43265 27663 43299
rect 27663 43265 27672 43299
rect 27620 43256 27672 43265
rect 28448 43256 28500 43308
rect 29000 43256 29052 43308
rect 29644 43299 29696 43308
rect 29644 43265 29653 43299
rect 29653 43265 29687 43299
rect 29687 43265 29696 43299
rect 29644 43256 29696 43265
rect 18420 43052 18472 43104
rect 18604 43095 18656 43104
rect 18604 43061 18613 43095
rect 18613 43061 18647 43095
rect 18647 43061 18656 43095
rect 18604 43052 18656 43061
rect 18880 43095 18932 43104
rect 18880 43061 18889 43095
rect 18889 43061 18923 43095
rect 18923 43061 18932 43095
rect 21732 43120 21784 43172
rect 18880 43052 18932 43061
rect 21180 43052 21232 43104
rect 22100 43120 22152 43172
rect 22928 43095 22980 43104
rect 22928 43061 22937 43095
rect 22937 43061 22971 43095
rect 22971 43061 22980 43095
rect 22928 43052 22980 43061
rect 24216 43052 24268 43104
rect 32036 43188 32088 43240
rect 37464 43324 37516 43376
rect 32220 43256 32272 43308
rect 33048 43299 33100 43308
rect 33048 43265 33057 43299
rect 33057 43265 33091 43299
rect 33091 43265 33100 43299
rect 33048 43256 33100 43265
rect 35348 43299 35400 43308
rect 35348 43265 35357 43299
rect 35357 43265 35391 43299
rect 35391 43265 35400 43299
rect 35348 43256 35400 43265
rect 36820 43299 36872 43308
rect 36820 43265 36829 43299
rect 36829 43265 36863 43299
rect 36863 43265 36872 43299
rect 36820 43256 36872 43265
rect 39764 43256 39816 43308
rect 41052 43299 41104 43308
rect 41052 43265 41061 43299
rect 41061 43265 41095 43299
rect 41095 43265 41104 43299
rect 41052 43256 41104 43265
rect 41788 43299 41840 43308
rect 41788 43265 41797 43299
rect 41797 43265 41831 43299
rect 41831 43265 41840 43299
rect 41788 43256 41840 43265
rect 38936 43231 38988 43240
rect 38936 43197 38945 43231
rect 38945 43197 38979 43231
rect 38979 43197 38988 43231
rect 38936 43188 38988 43197
rect 24768 43120 24820 43172
rect 25596 43163 25648 43172
rect 24492 43052 24544 43104
rect 25596 43129 25605 43163
rect 25605 43129 25639 43163
rect 25639 43129 25648 43163
rect 25596 43120 25648 43129
rect 27436 43163 27488 43172
rect 27436 43129 27445 43163
rect 27445 43129 27479 43163
rect 27479 43129 27488 43163
rect 27436 43120 27488 43129
rect 25964 43095 26016 43104
rect 25964 43061 25973 43095
rect 25973 43061 26007 43095
rect 26007 43061 26016 43095
rect 25964 43052 26016 43061
rect 26792 43052 26844 43104
rect 30932 43120 30984 43172
rect 34980 43163 35032 43172
rect 34980 43129 34989 43163
rect 34989 43129 35023 43163
rect 35023 43129 35032 43163
rect 34980 43120 35032 43129
rect 36544 43163 36596 43172
rect 30196 43052 30248 43104
rect 33048 43052 33100 43104
rect 33416 43052 33468 43104
rect 34244 43052 34296 43104
rect 36544 43129 36553 43163
rect 36553 43129 36587 43163
rect 36587 43129 36596 43163
rect 36544 43120 36596 43129
rect 36636 43163 36688 43172
rect 36636 43129 36645 43163
rect 36645 43129 36679 43163
rect 36679 43129 36688 43163
rect 36636 43120 36688 43129
rect 38108 43052 38160 43104
rect 38476 43095 38528 43104
rect 38476 43061 38485 43095
rect 38485 43061 38519 43095
rect 38519 43061 38528 43095
rect 38476 43052 38528 43061
rect 39488 43052 39540 43104
rect 42616 43188 42668 43240
rect 42064 43120 42116 43172
rect 40868 43052 40920 43104
rect 41788 43052 41840 43104
rect 42340 43052 42392 43104
rect 42524 43120 42576 43172
rect 43996 43120 44048 43172
rect 43536 43052 43588 43104
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 16488 42848 16540 42900
rect 18420 42848 18472 42900
rect 18972 42891 19024 42900
rect 18972 42857 18981 42891
rect 18981 42857 19015 42891
rect 19015 42857 19024 42891
rect 18972 42848 19024 42857
rect 21916 42848 21968 42900
rect 24768 42891 24820 42900
rect 24768 42857 24777 42891
rect 24777 42857 24811 42891
rect 24811 42857 24820 42891
rect 24768 42848 24820 42857
rect 26884 42891 26936 42900
rect 26884 42857 26893 42891
rect 26893 42857 26927 42891
rect 26927 42857 26936 42891
rect 26884 42848 26936 42857
rect 32220 42848 32272 42900
rect 33048 42891 33100 42900
rect 33048 42857 33057 42891
rect 33057 42857 33091 42891
rect 33091 42857 33100 42891
rect 33048 42848 33100 42857
rect 36544 42848 36596 42900
rect 38200 42848 38252 42900
rect 40776 42891 40828 42900
rect 16304 42780 16356 42832
rect 16580 42823 16632 42832
rect 16580 42789 16589 42823
rect 16589 42789 16623 42823
rect 16623 42789 16632 42823
rect 16580 42780 16632 42789
rect 18880 42780 18932 42832
rect 19248 42823 19300 42832
rect 19248 42789 19257 42823
rect 19257 42789 19291 42823
rect 19291 42789 19300 42823
rect 19248 42780 19300 42789
rect 19432 42780 19484 42832
rect 15936 42712 15988 42764
rect 18972 42712 19024 42764
rect 21180 42780 21232 42832
rect 21824 42780 21876 42832
rect 22100 42823 22152 42832
rect 22100 42789 22109 42823
rect 22109 42789 22143 42823
rect 22143 42789 22152 42823
rect 22100 42780 22152 42789
rect 22928 42780 22980 42832
rect 24952 42780 25004 42832
rect 25964 42780 26016 42832
rect 28448 42780 28500 42832
rect 28816 42823 28868 42832
rect 28816 42789 28825 42823
rect 28825 42789 28859 42823
rect 28859 42789 28868 42823
rect 28816 42780 28868 42789
rect 29644 42780 29696 42832
rect 30196 42780 30248 42832
rect 34796 42823 34848 42832
rect 34796 42789 34805 42823
rect 34805 42789 34839 42823
rect 34839 42789 34848 42823
rect 34796 42780 34848 42789
rect 34980 42780 35032 42832
rect 36728 42780 36780 42832
rect 40776 42857 40785 42891
rect 40785 42857 40819 42891
rect 40819 42857 40828 42891
rect 40776 42848 40828 42857
rect 41512 42848 41564 42900
rect 40868 42780 40920 42832
rect 41144 42823 41196 42832
rect 41144 42789 41153 42823
rect 41153 42789 41187 42823
rect 41187 42789 41196 42823
rect 41144 42780 41196 42789
rect 43536 42823 43588 42832
rect 43536 42789 43545 42823
rect 43545 42789 43579 42823
rect 43579 42789 43588 42823
rect 43536 42780 43588 42789
rect 21364 42712 21416 42764
rect 23848 42755 23900 42764
rect 23848 42721 23857 42755
rect 23857 42721 23891 42755
rect 23891 42721 23900 42755
rect 23848 42712 23900 42721
rect 25596 42755 25648 42764
rect 25596 42721 25605 42755
rect 25605 42721 25639 42755
rect 25639 42721 25648 42755
rect 25596 42712 25648 42721
rect 27160 42712 27212 42764
rect 27344 42755 27396 42764
rect 27344 42721 27353 42755
rect 27353 42721 27387 42755
rect 27387 42721 27396 42755
rect 27344 42712 27396 42721
rect 28356 42712 28408 42764
rect 35348 42755 35400 42764
rect 35348 42721 35357 42755
rect 35357 42721 35391 42755
rect 35391 42721 35400 42755
rect 35348 42712 35400 42721
rect 36084 42712 36136 42764
rect 36176 42755 36228 42764
rect 36176 42721 36185 42755
rect 36185 42721 36219 42755
rect 36219 42721 36228 42755
rect 36176 42712 36228 42721
rect 38016 42712 38068 42764
rect 38108 42712 38160 42764
rect 38844 42712 38896 42764
rect 16212 42644 16264 42696
rect 19156 42687 19208 42696
rect 19156 42653 19165 42687
rect 19165 42653 19199 42687
rect 19199 42653 19208 42687
rect 19156 42644 19208 42653
rect 24216 42644 24268 42696
rect 24676 42644 24728 42696
rect 28724 42687 28776 42696
rect 28724 42653 28733 42687
rect 28733 42653 28767 42687
rect 28767 42653 28776 42687
rect 28724 42644 28776 42653
rect 30748 42644 30800 42696
rect 32680 42687 32732 42696
rect 32680 42653 32689 42687
rect 32689 42653 32723 42687
rect 32723 42653 32732 42687
rect 32680 42644 32732 42653
rect 34704 42687 34756 42696
rect 34704 42653 34713 42687
rect 34713 42653 34747 42687
rect 34747 42653 34756 42687
rect 34704 42644 34756 42653
rect 36820 42644 36872 42696
rect 38476 42644 38528 42696
rect 39212 42687 39264 42696
rect 39212 42653 39221 42687
rect 39221 42653 39255 42687
rect 39255 42653 39264 42687
rect 39212 42644 39264 42653
rect 17132 42576 17184 42628
rect 22560 42619 22612 42628
rect 22560 42585 22569 42619
rect 22569 42585 22603 42619
rect 22603 42585 22612 42619
rect 22560 42576 22612 42585
rect 27068 42576 27120 42628
rect 28080 42576 28132 42628
rect 32956 42576 33008 42628
rect 36176 42576 36228 42628
rect 40316 42576 40368 42628
rect 42616 42644 42668 42696
rect 43444 42687 43496 42696
rect 43444 42653 43453 42687
rect 43453 42653 43487 42687
rect 43487 42653 43496 42687
rect 43444 42644 43496 42653
rect 41788 42576 41840 42628
rect 15936 42551 15988 42560
rect 15936 42517 15945 42551
rect 15945 42517 15979 42551
rect 15979 42517 15988 42551
rect 15936 42508 15988 42517
rect 21732 42551 21784 42560
rect 21732 42517 21741 42551
rect 21741 42517 21775 42551
rect 21775 42517 21784 42551
rect 21732 42508 21784 42517
rect 28816 42508 28868 42560
rect 29092 42508 29144 42560
rect 36544 42508 36596 42560
rect 38476 42551 38528 42560
rect 38476 42517 38485 42551
rect 38485 42517 38519 42551
rect 38519 42517 38528 42551
rect 38476 42508 38528 42517
rect 40132 42551 40184 42560
rect 40132 42517 40141 42551
rect 40141 42517 40175 42551
rect 40175 42517 40184 42551
rect 40132 42508 40184 42517
rect 42340 42551 42392 42560
rect 42340 42517 42349 42551
rect 42349 42517 42383 42551
rect 42383 42517 42392 42551
rect 42340 42508 42392 42517
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 16212 42304 16264 42356
rect 16304 42304 16356 42356
rect 16672 42304 16724 42356
rect 19156 42304 19208 42356
rect 21364 42347 21416 42356
rect 21364 42313 21373 42347
rect 21373 42313 21407 42347
rect 21407 42313 21416 42347
rect 21364 42304 21416 42313
rect 22928 42347 22980 42356
rect 22928 42313 22937 42347
rect 22937 42313 22971 42347
rect 22971 42313 22980 42347
rect 22928 42304 22980 42313
rect 27344 42304 27396 42356
rect 28632 42304 28684 42356
rect 29092 42347 29144 42356
rect 29092 42313 29101 42347
rect 29101 42313 29135 42347
rect 29135 42313 29144 42347
rect 29092 42304 29144 42313
rect 32220 42304 32272 42356
rect 36176 42304 36228 42356
rect 40132 42304 40184 42356
rect 21732 42236 21784 42288
rect 21824 42236 21876 42288
rect 24952 42236 25004 42288
rect 27160 42236 27212 42288
rect 22008 42211 22060 42220
rect 22008 42177 22017 42211
rect 22017 42177 22051 42211
rect 22051 42177 22060 42211
rect 22008 42168 22060 42177
rect 28356 42168 28408 42220
rect 15568 42143 15620 42152
rect 15568 42109 15577 42143
rect 15577 42109 15611 42143
rect 15611 42109 15620 42143
rect 15568 42100 15620 42109
rect 20168 42100 20220 42152
rect 21548 42100 21600 42152
rect 16212 42032 16264 42084
rect 14924 41964 14976 42016
rect 18972 41964 19024 42016
rect 19340 41964 19392 42016
rect 19892 42032 19944 42084
rect 22100 42075 22152 42084
rect 22100 42041 22109 42075
rect 22109 42041 22143 42075
rect 22143 42041 22152 42075
rect 22652 42075 22704 42084
rect 22100 42032 22152 42041
rect 22652 42041 22661 42075
rect 22661 42041 22695 42075
rect 22695 42041 22704 42075
rect 22652 42032 22704 42041
rect 25780 42143 25832 42152
rect 25780 42109 25789 42143
rect 25789 42109 25823 42143
rect 25823 42109 25832 42143
rect 25780 42100 25832 42109
rect 26516 42100 26568 42152
rect 27620 42100 27672 42152
rect 25136 42075 25188 42084
rect 25136 42041 25145 42075
rect 25145 42041 25179 42075
rect 25179 42041 25188 42075
rect 25136 42032 25188 42041
rect 23848 42007 23900 42016
rect 23848 41973 23857 42007
rect 23857 41973 23891 42007
rect 23891 41973 23900 42007
rect 23848 41964 23900 41973
rect 24584 42007 24636 42016
rect 24584 41973 24593 42007
rect 24593 41973 24627 42007
rect 24627 41973 24636 42007
rect 24584 41964 24636 41973
rect 25044 41964 25096 42016
rect 26976 42032 27028 42084
rect 25964 41964 26016 42016
rect 26516 41964 26568 42016
rect 27896 42032 27948 42084
rect 31208 42100 31260 42152
rect 33508 42236 33560 42288
rect 37924 42236 37976 42288
rect 43536 42304 43588 42356
rect 43076 42236 43128 42288
rect 43720 42236 43772 42288
rect 43812 42236 43864 42288
rect 44180 42236 44232 42288
rect 32680 42211 32732 42220
rect 32680 42177 32689 42211
rect 32689 42177 32723 42211
rect 32723 42177 32732 42211
rect 32680 42168 32732 42177
rect 35624 42211 35676 42220
rect 35624 42177 35633 42211
rect 35633 42177 35667 42211
rect 35667 42177 35676 42211
rect 35624 42168 35676 42177
rect 36544 42211 36596 42220
rect 36544 42177 36553 42211
rect 36553 42177 36587 42211
rect 36587 42177 36596 42211
rect 36544 42168 36596 42177
rect 36820 42211 36872 42220
rect 36820 42177 36829 42211
rect 36829 42177 36863 42211
rect 36863 42177 36872 42211
rect 36820 42168 36872 42177
rect 38016 42168 38068 42220
rect 39488 42168 39540 42220
rect 40776 42211 40828 42220
rect 40776 42177 40785 42211
rect 40785 42177 40819 42211
rect 40819 42177 40828 42211
rect 40776 42168 40828 42177
rect 43444 42168 43496 42220
rect 32220 42100 32272 42152
rect 34060 42100 34112 42152
rect 38200 42143 38252 42152
rect 28816 41964 28868 42016
rect 30196 42007 30248 42016
rect 30196 41973 30205 42007
rect 30205 41973 30239 42007
rect 30239 41973 30248 42007
rect 30196 41964 30248 41973
rect 30748 41964 30800 42016
rect 33048 42007 33100 42016
rect 33048 41973 33057 42007
rect 33057 41973 33091 42007
rect 33091 41973 33100 42007
rect 33048 41964 33100 41973
rect 33968 41964 34020 42016
rect 34152 42007 34204 42016
rect 34152 41973 34161 42007
rect 34161 41973 34195 42007
rect 34195 41973 34204 42007
rect 34152 41964 34204 41973
rect 38200 42109 38209 42143
rect 38209 42109 38243 42143
rect 38243 42109 38252 42143
rect 38200 42100 38252 42109
rect 34980 42075 35032 42084
rect 34980 42041 34989 42075
rect 34989 42041 35023 42075
rect 35023 42041 35032 42075
rect 34980 42032 35032 42041
rect 36636 42075 36688 42084
rect 36636 42041 36645 42075
rect 36645 42041 36679 42075
rect 36679 42041 36688 42075
rect 36636 42032 36688 42041
rect 38292 42032 38344 42084
rect 40132 42032 40184 42084
rect 41972 42032 42024 42084
rect 42340 42075 42392 42084
rect 42340 42041 42349 42075
rect 42349 42041 42383 42075
rect 42383 42041 42392 42075
rect 42340 42032 42392 42041
rect 43904 42075 43956 42084
rect 39580 42007 39632 42016
rect 39580 41973 39589 42007
rect 39589 41973 39623 42007
rect 39623 41973 39632 42007
rect 39580 41964 39632 41973
rect 39948 42007 40000 42016
rect 39948 41973 39957 42007
rect 39957 41973 39991 42007
rect 39991 41973 40000 42007
rect 39948 41964 40000 41973
rect 41328 41964 41380 42016
rect 42064 42007 42116 42016
rect 42064 41973 42073 42007
rect 42073 41973 42107 42007
rect 42107 41973 42116 42007
rect 43904 42041 43913 42075
rect 43913 42041 43947 42075
rect 43947 42041 43956 42075
rect 43904 42032 43956 42041
rect 43996 42075 44048 42084
rect 43996 42041 44005 42075
rect 44005 42041 44039 42075
rect 44039 42041 44048 42075
rect 43996 42032 44048 42041
rect 42064 41964 42116 41973
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 19340 41760 19392 41812
rect 21272 41803 21324 41812
rect 21272 41769 21281 41803
rect 21281 41769 21315 41803
rect 21315 41769 21324 41803
rect 21272 41760 21324 41769
rect 22100 41803 22152 41812
rect 22100 41769 22109 41803
rect 22109 41769 22143 41803
rect 22143 41769 22152 41803
rect 22100 41760 22152 41769
rect 24676 41803 24728 41812
rect 24676 41769 24685 41803
rect 24685 41769 24719 41803
rect 24719 41769 24728 41803
rect 24676 41760 24728 41769
rect 26976 41803 27028 41812
rect 26976 41769 26985 41803
rect 26985 41769 27019 41803
rect 27019 41769 27028 41803
rect 26976 41760 27028 41769
rect 28724 41760 28776 41812
rect 30748 41803 30800 41812
rect 30748 41769 30757 41803
rect 30757 41769 30791 41803
rect 30791 41769 30800 41803
rect 30748 41760 30800 41769
rect 16672 41735 16724 41744
rect 16672 41701 16681 41735
rect 16681 41701 16715 41735
rect 16715 41701 16724 41735
rect 16672 41692 16724 41701
rect 17224 41735 17276 41744
rect 17224 41701 17233 41735
rect 17233 41701 17267 41735
rect 17267 41701 17276 41735
rect 17224 41692 17276 41701
rect 18696 41692 18748 41744
rect 22008 41692 22060 41744
rect 22836 41735 22888 41744
rect 22836 41701 22845 41735
rect 22845 41701 22879 41735
rect 22879 41701 22888 41735
rect 22836 41692 22888 41701
rect 23388 41735 23440 41744
rect 23388 41701 23397 41735
rect 23397 41701 23431 41735
rect 23431 41701 23440 41735
rect 23388 41692 23440 41701
rect 24952 41692 25004 41744
rect 25872 41692 25924 41744
rect 27988 41735 28040 41744
rect 27988 41701 27997 41735
rect 27997 41701 28031 41735
rect 28031 41701 28040 41735
rect 27988 41692 28040 41701
rect 29552 41735 29604 41744
rect 29552 41701 29561 41735
rect 29561 41701 29595 41735
rect 29595 41701 29604 41735
rect 29552 41692 29604 41701
rect 31208 41760 31260 41812
rect 34796 41760 34848 41812
rect 36636 41760 36688 41812
rect 38200 41803 38252 41812
rect 38200 41769 38209 41803
rect 38209 41769 38243 41803
rect 38243 41769 38252 41803
rect 38200 41760 38252 41769
rect 39212 41803 39264 41812
rect 39212 41769 39221 41803
rect 39221 41769 39255 41803
rect 39255 41769 39264 41803
rect 39212 41760 39264 41769
rect 40868 41760 40920 41812
rect 43904 41760 43956 41812
rect 33968 41735 34020 41744
rect 33968 41701 33977 41735
rect 33977 41701 34011 41735
rect 34011 41701 34020 41735
rect 33968 41692 34020 41701
rect 34060 41735 34112 41744
rect 34060 41701 34069 41735
rect 34069 41701 34103 41735
rect 34103 41701 34112 41735
rect 34060 41692 34112 41701
rect 34704 41692 34756 41744
rect 35624 41735 35676 41744
rect 35624 41701 35633 41735
rect 35633 41701 35667 41735
rect 35667 41701 35676 41735
rect 35624 41692 35676 41701
rect 39948 41692 40000 41744
rect 40776 41692 40828 41744
rect 41972 41692 42024 41744
rect 42616 41692 42668 41744
rect 26516 41624 26568 41676
rect 31392 41624 31444 41676
rect 32312 41624 32364 41676
rect 37924 41667 37976 41676
rect 37924 41633 37933 41667
rect 37933 41633 37967 41667
rect 37967 41633 37976 41667
rect 37924 41624 37976 41633
rect 38108 41624 38160 41676
rect 43352 41624 43404 41676
rect 17408 41556 17460 41608
rect 18880 41556 18932 41608
rect 21180 41556 21232 41608
rect 23388 41556 23440 41608
rect 24400 41556 24452 41608
rect 27896 41599 27948 41608
rect 27896 41565 27905 41599
rect 27905 41565 27939 41599
rect 27939 41565 27948 41599
rect 27896 41556 27948 41565
rect 29460 41599 29512 41608
rect 29460 41565 29469 41599
rect 29469 41565 29503 41599
rect 29503 41565 29512 41599
rect 29460 41556 29512 41565
rect 29644 41556 29696 41608
rect 15384 41531 15436 41540
rect 15384 41497 15393 41531
rect 15393 41497 15427 41531
rect 15427 41497 15436 41531
rect 15384 41488 15436 41497
rect 26792 41488 26844 41540
rect 35992 41599 36044 41608
rect 35992 41565 36001 41599
rect 36001 41565 36035 41599
rect 36035 41565 36044 41599
rect 35992 41556 36044 41565
rect 39856 41599 39908 41608
rect 39856 41565 39865 41599
rect 39865 41565 39899 41599
rect 39899 41565 39908 41599
rect 39856 41556 39908 41565
rect 41604 41556 41656 41608
rect 41788 41599 41840 41608
rect 41788 41565 41797 41599
rect 41797 41565 41831 41599
rect 41831 41565 41840 41599
rect 41788 41556 41840 41565
rect 43996 41556 44048 41608
rect 34980 41488 35032 41540
rect 42064 41488 42116 41540
rect 13912 41420 13964 41472
rect 15568 41420 15620 41472
rect 25136 41420 25188 41472
rect 27620 41420 27672 41472
rect 32680 41463 32732 41472
rect 32680 41429 32689 41463
rect 32689 41429 32723 41463
rect 32723 41429 32732 41463
rect 32680 41420 32732 41429
rect 34612 41420 34664 41472
rect 34796 41420 34848 41472
rect 37372 41463 37424 41472
rect 37372 41429 37381 41463
rect 37381 41429 37415 41463
rect 37415 41429 37424 41463
rect 37372 41420 37424 41429
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 16672 41216 16724 41268
rect 17408 41259 17460 41268
rect 17408 41225 17417 41259
rect 17417 41225 17451 41259
rect 17451 41225 17460 41259
rect 17408 41216 17460 41225
rect 18696 41259 18748 41268
rect 18696 41225 18705 41259
rect 18705 41225 18739 41259
rect 18739 41225 18748 41259
rect 18696 41216 18748 41225
rect 22192 41216 22244 41268
rect 22836 41216 22888 41268
rect 25136 41216 25188 41268
rect 25872 41216 25924 41268
rect 21272 41148 21324 41200
rect 24952 41148 25004 41200
rect 17132 41080 17184 41132
rect 19892 41123 19944 41132
rect 19892 41089 19901 41123
rect 19901 41089 19935 41123
rect 19935 41089 19944 41123
rect 19892 41080 19944 41089
rect 22560 41123 22612 41132
rect 22560 41089 22569 41123
rect 22569 41089 22603 41123
rect 22603 41089 22612 41123
rect 22560 41080 22612 41089
rect 23020 41080 23072 41132
rect 14004 40876 14056 40928
rect 15384 40876 15436 40928
rect 16396 40876 16448 40928
rect 17960 40944 18012 40996
rect 19432 40944 19484 40996
rect 20536 40987 20588 40996
rect 20536 40953 20545 40987
rect 20545 40953 20579 40987
rect 20579 40953 20588 40987
rect 20536 40944 20588 40953
rect 21732 40944 21784 40996
rect 22192 40987 22244 40996
rect 22192 40953 22201 40987
rect 22201 40953 22235 40987
rect 22235 40953 22244 40987
rect 22192 40944 22244 40953
rect 22468 40944 22520 40996
rect 24768 41080 24820 41132
rect 26884 41080 26936 41132
rect 27988 41216 28040 41268
rect 29552 41259 29604 41268
rect 29552 41225 29561 41259
rect 29561 41225 29595 41259
rect 29595 41225 29604 41259
rect 29552 41216 29604 41225
rect 28448 41148 28500 41200
rect 33968 41216 34020 41268
rect 34612 41259 34664 41268
rect 34612 41225 34621 41259
rect 34621 41225 34655 41259
rect 34655 41225 34664 41259
rect 34612 41216 34664 41225
rect 38108 41216 38160 41268
rect 39580 41216 39632 41268
rect 40776 41259 40828 41268
rect 40776 41225 40785 41259
rect 40785 41225 40819 41259
rect 40819 41225 40828 41259
rect 40776 41216 40828 41225
rect 42340 41216 42392 41268
rect 43076 41259 43128 41268
rect 34060 41148 34112 41200
rect 35624 41148 35676 41200
rect 29460 41080 29512 41132
rect 32312 41080 32364 41132
rect 32680 41123 32732 41132
rect 32680 41089 32689 41123
rect 32689 41089 32723 41123
rect 32723 41089 32732 41123
rect 32680 41080 32732 41089
rect 35992 41080 36044 41132
rect 36084 41123 36136 41132
rect 36084 41089 36093 41123
rect 36093 41089 36127 41123
rect 36127 41089 36136 41123
rect 37372 41123 37424 41132
rect 36084 41080 36136 41089
rect 37372 41089 37381 41123
rect 37381 41089 37415 41123
rect 37415 41089 37424 41123
rect 37372 41080 37424 41089
rect 37924 41148 37976 41200
rect 42616 41191 42668 41200
rect 42616 41157 42625 41191
rect 42625 41157 42659 41191
rect 42659 41157 42668 41191
rect 42616 41148 42668 41157
rect 38108 41080 38160 41132
rect 38936 41080 38988 41132
rect 27620 41012 27672 41064
rect 30564 41012 30616 41064
rect 39856 41080 39908 41132
rect 43076 41225 43085 41259
rect 43085 41225 43119 41259
rect 43119 41225 43128 41259
rect 43076 41216 43128 41225
rect 43352 41123 43404 41132
rect 43352 41089 43361 41123
rect 43361 41089 43395 41123
rect 43395 41089 43404 41123
rect 43352 41080 43404 41089
rect 25136 40944 25188 40996
rect 28540 40944 28592 40996
rect 30196 40944 30248 40996
rect 33048 40987 33100 40996
rect 33048 40953 33051 40987
rect 33051 40953 33085 40987
rect 33085 40953 33100 40987
rect 33048 40944 33100 40953
rect 33324 40944 33376 40996
rect 35900 40987 35952 40996
rect 35900 40953 35909 40987
rect 35909 40953 35943 40987
rect 35943 40953 35952 40987
rect 35900 40944 35952 40953
rect 36636 40944 36688 40996
rect 37188 40944 37240 40996
rect 18880 40876 18932 40928
rect 21180 40876 21232 40928
rect 23388 40919 23440 40928
rect 23388 40885 23397 40919
rect 23397 40885 23431 40919
rect 23431 40885 23440 40919
rect 23388 40876 23440 40885
rect 26516 40919 26568 40928
rect 26516 40885 26525 40919
rect 26525 40885 26559 40919
rect 26559 40885 26568 40919
rect 26516 40876 26568 40885
rect 31392 40876 31444 40928
rect 35164 40919 35216 40928
rect 35164 40885 35173 40919
rect 35173 40885 35207 40919
rect 35207 40885 35216 40919
rect 35164 40876 35216 40885
rect 38384 40876 38436 40928
rect 39672 41012 39724 41064
rect 41420 41055 41472 41064
rect 41420 41021 41429 41055
rect 41429 41021 41463 41055
rect 41463 41021 41472 41055
rect 41420 41012 41472 41021
rect 39120 40876 39172 40928
rect 39948 40876 40000 40928
rect 41696 40876 41748 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 16396 40715 16448 40724
rect 16396 40681 16405 40715
rect 16405 40681 16439 40715
rect 16439 40681 16448 40715
rect 16396 40672 16448 40681
rect 17132 40715 17184 40724
rect 17132 40681 17141 40715
rect 17141 40681 17175 40715
rect 17175 40681 17184 40715
rect 17132 40672 17184 40681
rect 18144 40672 18196 40724
rect 19064 40672 19116 40724
rect 21732 40715 21784 40724
rect 21732 40681 21741 40715
rect 21741 40681 21775 40715
rect 21775 40681 21784 40715
rect 21732 40672 21784 40681
rect 22192 40672 22244 40724
rect 24400 40715 24452 40724
rect 16212 40604 16264 40656
rect 17408 40647 17460 40656
rect 17408 40613 17417 40647
rect 17417 40613 17451 40647
rect 17451 40613 17460 40647
rect 17408 40604 17460 40613
rect 19892 40647 19944 40656
rect 19892 40613 19901 40647
rect 19901 40613 19935 40647
rect 19935 40613 19944 40647
rect 19892 40604 19944 40613
rect 24400 40681 24409 40715
rect 24409 40681 24443 40715
rect 24443 40681 24452 40715
rect 24400 40672 24452 40681
rect 24768 40715 24820 40724
rect 24768 40681 24777 40715
rect 24777 40681 24811 40715
rect 24811 40681 24820 40715
rect 24768 40672 24820 40681
rect 27896 40715 27948 40724
rect 27896 40681 27905 40715
rect 27905 40681 27939 40715
rect 27939 40681 27948 40715
rect 27896 40672 27948 40681
rect 28540 40672 28592 40724
rect 29552 40672 29604 40724
rect 30564 40715 30616 40724
rect 30564 40681 30573 40715
rect 30573 40681 30607 40715
rect 30607 40681 30616 40715
rect 30564 40672 30616 40681
rect 34796 40672 34848 40724
rect 35164 40672 35216 40724
rect 35900 40672 35952 40724
rect 35992 40715 36044 40724
rect 35992 40681 36001 40715
rect 36001 40681 36035 40715
rect 36035 40681 36044 40715
rect 35992 40672 36044 40681
rect 37372 40672 37424 40724
rect 38936 40715 38988 40724
rect 38936 40681 38945 40715
rect 38945 40681 38979 40715
rect 38979 40681 38988 40715
rect 38936 40672 38988 40681
rect 41604 40715 41656 40724
rect 41604 40681 41613 40715
rect 41613 40681 41647 40715
rect 41647 40681 41656 40715
rect 41604 40672 41656 40681
rect 22652 40604 22704 40656
rect 25044 40647 25096 40656
rect 25044 40613 25053 40647
rect 25053 40613 25087 40647
rect 25087 40613 25096 40647
rect 25044 40604 25096 40613
rect 25872 40604 25924 40656
rect 33324 40604 33376 40656
rect 35256 40604 35308 40656
rect 37188 40604 37240 40656
rect 41880 40647 41932 40656
rect 41880 40613 41889 40647
rect 41889 40613 41923 40647
rect 41923 40613 41932 40647
rect 41880 40604 41932 40613
rect 42432 40647 42484 40656
rect 42432 40613 42441 40647
rect 42441 40613 42475 40647
rect 42475 40613 42484 40647
rect 42432 40604 42484 40613
rect 42616 40604 42668 40656
rect 18604 40536 18656 40588
rect 21548 40536 21600 40588
rect 24308 40536 24360 40588
rect 26976 40579 27028 40588
rect 26976 40545 26985 40579
rect 26985 40545 27019 40579
rect 27019 40545 27028 40579
rect 26976 40536 27028 40545
rect 27344 40536 27396 40588
rect 30564 40579 30616 40588
rect 30564 40545 30573 40579
rect 30573 40545 30607 40579
rect 30607 40545 30616 40579
rect 30564 40536 30616 40545
rect 31392 40536 31444 40588
rect 15292 40468 15344 40520
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 17960 40511 18012 40520
rect 17960 40477 17969 40511
rect 17969 40477 18003 40511
rect 18003 40477 18012 40511
rect 17960 40468 18012 40477
rect 18696 40468 18748 40520
rect 22744 40468 22796 40520
rect 24952 40511 25004 40520
rect 24952 40477 24961 40511
rect 24961 40477 24995 40511
rect 24995 40477 25004 40511
rect 24952 40468 25004 40477
rect 28908 40468 28960 40520
rect 32220 40536 32272 40588
rect 34244 40536 34296 40588
rect 27160 40400 27212 40452
rect 32496 40468 32548 40520
rect 32680 40511 32732 40520
rect 32680 40477 32689 40511
rect 32689 40477 32723 40511
rect 32723 40477 32732 40511
rect 32680 40468 32732 40477
rect 34704 40511 34756 40520
rect 34704 40477 34713 40511
rect 34713 40477 34747 40511
rect 34747 40477 34756 40511
rect 34704 40468 34756 40477
rect 36544 40536 36596 40588
rect 38936 40536 38988 40588
rect 39580 40579 39632 40588
rect 39580 40545 39589 40579
rect 39589 40545 39623 40579
rect 39623 40545 39632 40579
rect 39580 40536 39632 40545
rect 43812 40536 43864 40588
rect 39672 40468 39724 40520
rect 39856 40511 39908 40520
rect 39856 40477 39865 40511
rect 39865 40477 39899 40511
rect 39899 40477 39908 40511
rect 39856 40468 39908 40477
rect 41788 40511 41840 40520
rect 41788 40477 41797 40511
rect 41797 40477 41831 40511
rect 41831 40477 41840 40511
rect 41788 40468 41840 40477
rect 38384 40400 38436 40452
rect 16120 40332 16172 40384
rect 19156 40375 19208 40384
rect 19156 40341 19165 40375
rect 19165 40341 19199 40375
rect 19199 40341 19208 40375
rect 19156 40332 19208 40341
rect 38016 40375 38068 40384
rect 38016 40341 38025 40375
rect 38025 40341 38059 40375
rect 38059 40341 38068 40375
rect 38016 40332 38068 40341
rect 40500 40375 40552 40384
rect 40500 40341 40509 40375
rect 40509 40341 40543 40375
rect 40543 40341 40552 40375
rect 40500 40332 40552 40341
rect 42800 40332 42852 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 17408 40171 17460 40180
rect 17408 40137 17417 40171
rect 17417 40137 17451 40171
rect 17451 40137 17460 40171
rect 17408 40128 17460 40137
rect 18604 40171 18656 40180
rect 18604 40137 18613 40171
rect 18613 40137 18647 40171
rect 18647 40137 18656 40171
rect 18604 40128 18656 40137
rect 19432 40128 19484 40180
rect 17316 40060 17368 40112
rect 22468 40128 22520 40180
rect 22836 40128 22888 40180
rect 25044 40128 25096 40180
rect 27344 40128 27396 40180
rect 28540 40171 28592 40180
rect 28540 40137 28549 40171
rect 28549 40137 28583 40171
rect 28583 40137 28592 40171
rect 28540 40128 28592 40137
rect 28908 40171 28960 40180
rect 28908 40137 28917 40171
rect 28917 40137 28951 40171
rect 28951 40137 28960 40171
rect 28908 40128 28960 40137
rect 32220 40171 32272 40180
rect 32220 40137 32229 40171
rect 32229 40137 32263 40171
rect 32263 40137 32272 40171
rect 32220 40128 32272 40137
rect 32864 40128 32916 40180
rect 34244 40171 34296 40180
rect 16120 39967 16172 39976
rect 16120 39933 16129 39967
rect 16129 39933 16163 39967
rect 16163 39933 16172 39967
rect 16120 39924 16172 39933
rect 19064 39967 19116 39976
rect 19064 39933 19073 39967
rect 19073 39933 19107 39967
rect 19107 39933 19116 39967
rect 19064 39924 19116 39933
rect 20260 39924 20312 39976
rect 22376 40060 22428 40112
rect 23112 40060 23164 40112
rect 26976 40103 27028 40112
rect 26976 40069 26985 40103
rect 26985 40069 27019 40103
rect 27019 40069 27028 40103
rect 26976 40060 27028 40069
rect 32496 40103 32548 40112
rect 32496 40069 32505 40103
rect 32505 40069 32539 40103
rect 32539 40069 32548 40103
rect 32496 40060 32548 40069
rect 27712 39992 27764 40044
rect 23756 39924 23808 39976
rect 16212 39856 16264 39908
rect 20628 39856 20680 39908
rect 22192 39899 22244 39908
rect 22192 39865 22201 39899
rect 22201 39865 22235 39899
rect 22235 39865 22244 39899
rect 22192 39856 22244 39865
rect 24952 39856 25004 39908
rect 15292 39788 15344 39840
rect 21548 39788 21600 39840
rect 22652 39788 22704 39840
rect 23848 39788 23900 39840
rect 24308 39788 24360 39840
rect 26792 39924 26844 39976
rect 26056 39856 26108 39908
rect 30932 39967 30984 39976
rect 30932 39933 30941 39967
rect 30941 39933 30975 39967
rect 30975 39933 30984 39967
rect 30932 39924 30984 39933
rect 31392 39967 31444 39976
rect 31392 39933 31401 39967
rect 31401 39933 31435 39967
rect 31435 39933 31444 39967
rect 31392 39924 31444 39933
rect 33232 39967 33284 39976
rect 33232 39933 33241 39967
rect 33241 39933 33275 39967
rect 33275 39933 33284 39967
rect 33232 39924 33284 39933
rect 34244 40137 34253 40171
rect 34253 40137 34287 40171
rect 34287 40137 34296 40171
rect 34244 40128 34296 40137
rect 35256 40128 35308 40180
rect 35348 40128 35400 40180
rect 37924 40128 37976 40180
rect 39580 40171 39632 40180
rect 39580 40137 39589 40171
rect 39589 40137 39623 40171
rect 39623 40137 39632 40171
rect 39580 40128 39632 40137
rect 41696 40128 41748 40180
rect 41788 40128 41840 40180
rect 44180 40128 44232 40180
rect 36544 40060 36596 40112
rect 42248 40060 42300 40112
rect 34704 39992 34756 40044
rect 35532 39992 35584 40044
rect 36912 39992 36964 40044
rect 38568 40035 38620 40044
rect 38568 40001 38577 40035
rect 38577 40001 38611 40035
rect 38611 40001 38620 40035
rect 38568 39992 38620 40001
rect 39120 39992 39172 40044
rect 35808 39967 35860 39976
rect 35808 39933 35817 39967
rect 35817 39933 35851 39967
rect 35851 39933 35860 39967
rect 35808 39924 35860 39933
rect 37924 39967 37976 39976
rect 37924 39933 37933 39967
rect 37933 39933 37967 39967
rect 37967 39933 37976 39967
rect 37924 39924 37976 39933
rect 38016 39924 38068 39976
rect 39580 39924 39632 39976
rect 40500 39967 40552 39976
rect 40500 39933 40509 39967
rect 40509 39933 40543 39967
rect 40543 39933 40552 39967
rect 40500 39924 40552 39933
rect 41880 39992 41932 40044
rect 42800 40035 42852 40044
rect 42800 40001 42809 40035
rect 42809 40001 42843 40035
rect 42843 40001 42852 40035
rect 43076 40035 43128 40044
rect 42800 39992 42852 40001
rect 43076 40001 43085 40035
rect 43085 40001 43119 40035
rect 43119 40001 43128 40035
rect 43076 39992 43128 40001
rect 25504 39788 25556 39840
rect 27436 39831 27488 39840
rect 27436 39797 27445 39831
rect 27445 39797 27479 39831
rect 27479 39797 27488 39831
rect 27436 39788 27488 39797
rect 27620 39831 27672 39840
rect 27620 39797 27629 39831
rect 27629 39797 27663 39831
rect 27663 39797 27672 39831
rect 27620 39788 27672 39797
rect 30196 39831 30248 39840
rect 30196 39797 30205 39831
rect 30205 39797 30239 39831
rect 30239 39797 30248 39831
rect 30196 39788 30248 39797
rect 30564 39831 30616 39840
rect 30564 39797 30573 39831
rect 30573 39797 30607 39831
rect 30607 39797 30616 39831
rect 30564 39788 30616 39797
rect 30840 39788 30892 39840
rect 36636 39856 36688 39908
rect 40776 39899 40828 39908
rect 40776 39865 40794 39899
rect 40794 39865 40828 39899
rect 40776 39856 40828 39865
rect 36820 39788 36872 39840
rect 38936 39788 38988 39840
rect 41328 39788 41380 39840
rect 43352 39788 43404 39840
rect 43812 39831 43864 39840
rect 43812 39797 43821 39831
rect 43821 39797 43855 39831
rect 43855 39797 43864 39831
rect 43812 39788 43864 39797
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 17960 39584 18012 39636
rect 16212 39516 16264 39568
rect 18052 39559 18104 39568
rect 18052 39525 18061 39559
rect 18061 39525 18095 39559
rect 18095 39525 18104 39559
rect 18052 39516 18104 39525
rect 22192 39584 22244 39636
rect 22744 39627 22796 39636
rect 22744 39593 22753 39627
rect 22753 39593 22787 39627
rect 22787 39593 22796 39627
rect 22744 39584 22796 39593
rect 24952 39627 25004 39636
rect 24952 39593 24961 39627
rect 24961 39593 24995 39627
rect 24995 39593 25004 39627
rect 24952 39584 25004 39593
rect 25964 39584 26016 39636
rect 27712 39627 27764 39636
rect 27712 39593 27721 39627
rect 27721 39593 27755 39627
rect 27755 39593 27764 39627
rect 27712 39584 27764 39593
rect 28540 39584 28592 39636
rect 30932 39627 30984 39636
rect 30932 39593 30941 39627
rect 30941 39593 30975 39627
rect 30975 39593 30984 39627
rect 30932 39584 30984 39593
rect 32220 39627 32272 39636
rect 32220 39593 32229 39627
rect 32229 39593 32263 39627
rect 32263 39593 32272 39627
rect 32220 39584 32272 39593
rect 33232 39627 33284 39636
rect 33232 39593 33241 39627
rect 33241 39593 33275 39627
rect 33275 39593 33284 39627
rect 33232 39584 33284 39593
rect 33416 39584 33468 39636
rect 18696 39559 18748 39568
rect 18696 39525 18705 39559
rect 18705 39525 18739 39559
rect 18739 39525 18748 39559
rect 18696 39516 18748 39525
rect 20628 39516 20680 39568
rect 22008 39516 22060 39568
rect 19616 39448 19668 39500
rect 20536 39448 20588 39500
rect 23296 39448 23348 39500
rect 24124 39448 24176 39500
rect 24584 39448 24636 39500
rect 27160 39516 27212 39568
rect 30196 39516 30248 39568
rect 31392 39516 31444 39568
rect 33324 39516 33376 39568
rect 36636 39584 36688 39636
rect 36820 39627 36872 39636
rect 36820 39593 36829 39627
rect 36829 39593 36863 39627
rect 36863 39593 36872 39627
rect 36820 39584 36872 39593
rect 38108 39584 38160 39636
rect 39120 39627 39172 39636
rect 39120 39593 39129 39627
rect 39129 39593 39163 39627
rect 39163 39593 39172 39627
rect 39120 39584 39172 39593
rect 41328 39584 41380 39636
rect 41880 39584 41932 39636
rect 42800 39627 42852 39636
rect 42800 39593 42809 39627
rect 42809 39593 42843 39627
rect 42843 39593 42852 39627
rect 42800 39584 42852 39593
rect 38660 39516 38712 39568
rect 38936 39516 38988 39568
rect 40776 39559 40828 39568
rect 40776 39525 40785 39559
rect 40785 39525 40819 39559
rect 40819 39525 40828 39559
rect 40776 39516 40828 39525
rect 41788 39559 41840 39568
rect 41788 39525 41797 39559
rect 41797 39525 41831 39559
rect 41831 39525 41840 39559
rect 41788 39516 41840 39525
rect 42432 39516 42484 39568
rect 43444 39516 43496 39568
rect 44180 39516 44232 39568
rect 16764 39380 16816 39432
rect 21456 39423 21508 39432
rect 21456 39389 21465 39423
rect 21465 39389 21499 39423
rect 21499 39389 21508 39423
rect 21456 39380 21508 39389
rect 21364 39312 21416 39364
rect 27252 39448 27304 39500
rect 31024 39491 31076 39500
rect 31024 39457 31033 39491
rect 31033 39457 31067 39491
rect 31067 39457 31076 39491
rect 31024 39448 31076 39457
rect 32036 39448 32088 39500
rect 34612 39491 34664 39500
rect 28264 39423 28316 39432
rect 28264 39389 28273 39423
rect 28273 39389 28307 39423
rect 28307 39389 28316 39423
rect 28264 39380 28316 39389
rect 32312 39380 32364 39432
rect 31852 39312 31904 39364
rect 34612 39457 34621 39491
rect 34621 39457 34655 39491
rect 34655 39457 34664 39491
rect 34612 39448 34664 39457
rect 38016 39448 38068 39500
rect 39856 39448 39908 39500
rect 40224 39448 40276 39500
rect 42248 39491 42300 39500
rect 42248 39457 42257 39491
rect 42257 39457 42291 39491
rect 42291 39457 42300 39491
rect 42248 39448 42300 39457
rect 33692 39423 33744 39432
rect 33692 39389 33701 39423
rect 33701 39389 33735 39423
rect 33735 39389 33744 39423
rect 33692 39380 33744 39389
rect 35532 39423 35584 39432
rect 35532 39389 35541 39423
rect 35541 39389 35575 39423
rect 35575 39389 35584 39423
rect 35532 39380 35584 39389
rect 38752 39423 38804 39432
rect 38752 39389 38761 39423
rect 38761 39389 38795 39423
rect 38795 39389 38804 39423
rect 38752 39380 38804 39389
rect 42708 39380 42760 39432
rect 36084 39355 36136 39364
rect 36084 39321 36093 39355
rect 36093 39321 36127 39355
rect 36127 39321 36136 39355
rect 36084 39312 36136 39321
rect 19064 39287 19116 39296
rect 19064 39253 19073 39287
rect 19073 39253 19107 39287
rect 19107 39253 19116 39287
rect 19064 39244 19116 39253
rect 19432 39244 19484 39296
rect 21088 39244 21140 39296
rect 24952 39244 25004 39296
rect 25504 39244 25556 39296
rect 28632 39244 28684 39296
rect 29184 39287 29236 39296
rect 29184 39253 29193 39287
rect 29193 39253 29227 39287
rect 29227 39253 29236 39287
rect 29184 39244 29236 39253
rect 29460 39287 29512 39296
rect 29460 39253 29469 39287
rect 29469 39253 29503 39287
rect 29503 39253 29512 39287
rect 29460 39244 29512 39253
rect 30932 39244 30984 39296
rect 35348 39244 35400 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 16212 39083 16264 39092
rect 16212 39049 16221 39083
rect 16221 39049 16255 39083
rect 16255 39049 16264 39083
rect 16212 39040 16264 39049
rect 18052 39040 18104 39092
rect 18604 39040 18656 39092
rect 13912 38947 13964 38956
rect 13912 38913 13921 38947
rect 13921 38913 13955 38947
rect 13955 38913 13964 38947
rect 13912 38904 13964 38913
rect 15292 38947 15344 38956
rect 15292 38913 15301 38947
rect 15301 38913 15335 38947
rect 15335 38913 15344 38947
rect 15292 38904 15344 38913
rect 19064 38947 19116 38956
rect 13636 38836 13688 38888
rect 13820 38836 13872 38888
rect 19064 38913 19073 38947
rect 19073 38913 19107 38947
rect 19107 38913 19116 38947
rect 19064 38904 19116 38913
rect 23388 39040 23440 39092
rect 27160 39040 27212 39092
rect 28540 39040 28592 39092
rect 28724 39040 28776 39092
rect 29184 39040 29236 39092
rect 31024 39040 31076 39092
rect 32036 39040 32088 39092
rect 32864 39083 32916 39092
rect 32864 39049 32873 39083
rect 32873 39049 32907 39083
rect 32907 39049 32916 39083
rect 34612 39083 34664 39092
rect 32864 39040 32916 39049
rect 22008 39015 22060 39024
rect 22008 38981 22017 39015
rect 22017 38981 22051 39015
rect 22051 38981 22060 39015
rect 23296 39015 23348 39024
rect 22008 38972 22060 38981
rect 23296 38981 23305 39015
rect 23305 38981 23339 39015
rect 23339 38981 23348 39015
rect 23296 38972 23348 38981
rect 25136 39015 25188 39024
rect 25136 38981 25145 39015
rect 25145 38981 25179 39015
rect 25179 38981 25188 39015
rect 25136 38972 25188 38981
rect 27068 38972 27120 39024
rect 21456 38904 21508 38956
rect 23020 38904 23072 38956
rect 13544 38700 13596 38752
rect 16488 38836 16540 38888
rect 18788 38836 18840 38888
rect 18052 38768 18104 38820
rect 19156 38836 19208 38888
rect 19616 38879 19668 38888
rect 19616 38845 19625 38879
rect 19625 38845 19659 38879
rect 19659 38845 19668 38879
rect 19616 38836 19668 38845
rect 21364 38879 21416 38888
rect 21364 38845 21373 38879
rect 21373 38845 21407 38879
rect 21407 38845 21416 38879
rect 21364 38836 21416 38845
rect 22008 38768 22060 38820
rect 15752 38743 15804 38752
rect 15752 38709 15761 38743
rect 15761 38709 15795 38743
rect 15795 38709 15804 38743
rect 15752 38700 15804 38709
rect 16764 38700 16816 38752
rect 20352 38700 20404 38752
rect 25504 38904 25556 38956
rect 28356 38904 28408 38956
rect 29460 38904 29512 38956
rect 29644 38947 29696 38956
rect 29644 38913 29653 38947
rect 29653 38913 29687 38947
rect 29687 38913 29696 38947
rect 29644 38904 29696 38913
rect 24492 38836 24544 38888
rect 25964 38836 26016 38888
rect 27436 38836 27488 38888
rect 27896 38879 27948 38888
rect 27896 38845 27905 38879
rect 27905 38845 27939 38879
rect 27939 38845 27948 38879
rect 27896 38836 27948 38845
rect 28172 38879 28224 38888
rect 28172 38845 28181 38879
rect 28181 38845 28215 38879
rect 28215 38845 28224 38879
rect 28172 38836 28224 38845
rect 31484 38836 31536 38888
rect 33232 38836 33284 38888
rect 34612 39049 34621 39083
rect 34621 39049 34655 39083
rect 34655 39049 34664 39083
rect 34612 39040 34664 39049
rect 36636 39083 36688 39092
rect 36636 39049 36645 39083
rect 36645 39049 36679 39083
rect 36679 39049 36688 39083
rect 36636 39040 36688 39049
rect 36912 39083 36964 39092
rect 36912 39049 36921 39083
rect 36921 39049 36955 39083
rect 36955 39049 36964 39083
rect 36912 39040 36964 39049
rect 38108 39040 38160 39092
rect 40224 39083 40276 39092
rect 36084 38972 36136 39024
rect 33692 38947 33744 38956
rect 33692 38913 33701 38947
rect 33701 38913 33735 38947
rect 33735 38913 33744 38947
rect 33692 38904 33744 38913
rect 24124 38811 24176 38820
rect 24124 38777 24133 38811
rect 24133 38777 24167 38811
rect 24167 38777 24176 38811
rect 24124 38768 24176 38777
rect 24860 38768 24912 38820
rect 25136 38768 25188 38820
rect 27252 38768 27304 38820
rect 28540 38768 28592 38820
rect 24584 38700 24636 38752
rect 26148 38743 26200 38752
rect 26148 38709 26157 38743
rect 26157 38709 26191 38743
rect 26191 38709 26200 38743
rect 26148 38700 26200 38709
rect 29184 38700 29236 38752
rect 30288 38768 30340 38820
rect 33140 38768 33192 38820
rect 35256 38879 35308 38888
rect 35256 38845 35265 38879
rect 35265 38845 35299 38879
rect 35299 38845 35308 38879
rect 35256 38836 35308 38845
rect 40224 39049 40233 39083
rect 40233 39049 40267 39083
rect 40267 39049 40276 39083
rect 40224 39040 40276 39049
rect 40776 39040 40828 39092
rect 41420 39083 41472 39092
rect 41420 39049 41429 39083
rect 41429 39049 41463 39083
rect 41463 39049 41472 39083
rect 41420 39040 41472 39049
rect 42708 39040 42760 39092
rect 43444 39083 43496 39092
rect 43444 39049 43453 39083
rect 43453 39049 43487 39083
rect 43487 39049 43496 39083
rect 43444 39040 43496 39049
rect 39580 38947 39632 38956
rect 38844 38879 38896 38888
rect 38844 38845 38853 38879
rect 38853 38845 38887 38879
rect 38887 38845 38896 38879
rect 38844 38836 38896 38845
rect 39580 38913 39589 38947
rect 39589 38913 39623 38947
rect 39623 38913 39632 38947
rect 39580 38904 39632 38913
rect 41236 38836 41288 38888
rect 41420 38836 41472 38888
rect 41788 38836 41840 38888
rect 44272 38836 44324 38888
rect 39120 38768 39172 38820
rect 31760 38743 31812 38752
rect 31760 38709 31769 38743
rect 31769 38709 31803 38743
rect 31803 38709 31812 38743
rect 31760 38700 31812 38709
rect 32128 38700 32180 38752
rect 33324 38700 33376 38752
rect 33600 38700 33652 38752
rect 35532 38743 35584 38752
rect 35532 38709 35541 38743
rect 35541 38709 35575 38743
rect 35575 38709 35584 38743
rect 35532 38700 35584 38709
rect 37372 38700 37424 38752
rect 38016 38743 38068 38752
rect 38016 38709 38025 38743
rect 38025 38709 38059 38743
rect 38059 38709 38068 38743
rect 38016 38700 38068 38709
rect 40960 38700 41012 38752
rect 41972 38700 42024 38752
rect 42340 38743 42392 38752
rect 42340 38709 42349 38743
rect 42349 38709 42383 38743
rect 42383 38709 42392 38743
rect 42340 38700 42392 38709
rect 44180 38700 44232 38752
rect 44456 38700 44508 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 16488 38539 16540 38548
rect 16488 38505 16497 38539
rect 16497 38505 16531 38539
rect 16531 38505 16540 38539
rect 16488 38496 16540 38505
rect 16764 38539 16816 38548
rect 16764 38505 16773 38539
rect 16773 38505 16807 38539
rect 16807 38505 16816 38539
rect 16764 38496 16816 38505
rect 17960 38539 18012 38548
rect 17960 38505 17969 38539
rect 17969 38505 18003 38539
rect 18003 38505 18012 38539
rect 17960 38496 18012 38505
rect 19432 38496 19484 38548
rect 21180 38539 21232 38548
rect 21180 38505 21189 38539
rect 21189 38505 21223 38539
rect 21223 38505 21232 38539
rect 21180 38496 21232 38505
rect 22284 38496 22336 38548
rect 24492 38496 24544 38548
rect 25964 38539 26016 38548
rect 25964 38505 25973 38539
rect 25973 38505 26007 38539
rect 26007 38505 26016 38539
rect 25964 38496 26016 38505
rect 28264 38539 28316 38548
rect 28264 38505 28273 38539
rect 28273 38505 28307 38539
rect 28307 38505 28316 38539
rect 28264 38496 28316 38505
rect 31852 38539 31904 38548
rect 31852 38505 31861 38539
rect 31861 38505 31895 38539
rect 31895 38505 31904 38539
rect 31852 38496 31904 38505
rect 35256 38539 35308 38548
rect 13820 38428 13872 38480
rect 15568 38428 15620 38480
rect 16120 38471 16172 38480
rect 15660 38403 15712 38412
rect 15660 38369 15669 38403
rect 15669 38369 15703 38403
rect 15703 38369 15712 38403
rect 15660 38360 15712 38369
rect 16120 38437 16129 38471
rect 16129 38437 16163 38471
rect 16163 38437 16172 38471
rect 16120 38428 16172 38437
rect 18880 38471 18932 38480
rect 18880 38437 18889 38471
rect 18889 38437 18923 38471
rect 18923 38437 18932 38471
rect 18880 38428 18932 38437
rect 23020 38428 23072 38480
rect 24952 38471 25004 38480
rect 24952 38437 24961 38471
rect 24961 38437 24995 38471
rect 24995 38437 25004 38471
rect 24952 38428 25004 38437
rect 26148 38428 26200 38480
rect 26608 38428 26660 38480
rect 28724 38428 28776 38480
rect 30288 38428 30340 38480
rect 30380 38428 30432 38480
rect 31760 38428 31812 38480
rect 17868 38360 17920 38412
rect 19156 38360 19208 38412
rect 20536 38360 20588 38412
rect 20904 38403 20956 38412
rect 20904 38369 20913 38403
rect 20913 38369 20947 38403
rect 20947 38369 20956 38403
rect 20904 38360 20956 38369
rect 21364 38403 21416 38412
rect 21364 38369 21373 38403
rect 21373 38369 21407 38403
rect 21407 38369 21416 38403
rect 21364 38360 21416 38369
rect 32220 38360 32272 38412
rect 35256 38505 35265 38539
rect 35265 38505 35299 38539
rect 35299 38505 35308 38539
rect 35256 38496 35308 38505
rect 38016 38496 38068 38548
rect 38844 38539 38896 38548
rect 33324 38428 33376 38480
rect 38844 38505 38853 38539
rect 38853 38505 38887 38539
rect 38887 38505 38896 38539
rect 38844 38496 38896 38505
rect 38752 38428 38804 38480
rect 40960 38428 41012 38480
rect 41788 38471 41840 38480
rect 41788 38437 41797 38471
rect 41797 38437 41831 38471
rect 41831 38437 41840 38471
rect 41788 38428 41840 38437
rect 41880 38471 41932 38480
rect 41880 38437 41889 38471
rect 41889 38437 41923 38471
rect 41923 38437 41932 38471
rect 41880 38428 41932 38437
rect 44272 38428 44324 38480
rect 33600 38360 33652 38412
rect 33968 38403 34020 38412
rect 33968 38369 33977 38403
rect 33977 38369 34011 38403
rect 34011 38369 34020 38403
rect 33968 38360 34020 38369
rect 35256 38403 35308 38412
rect 35256 38369 35265 38403
rect 35265 38369 35299 38403
rect 35299 38369 35308 38403
rect 35256 38360 35308 38369
rect 35440 38403 35492 38412
rect 35440 38369 35449 38403
rect 35449 38369 35483 38403
rect 35483 38369 35492 38403
rect 35440 38360 35492 38369
rect 36912 38360 36964 38412
rect 37740 38403 37792 38412
rect 37740 38369 37749 38403
rect 37749 38369 37783 38403
rect 37783 38369 37792 38403
rect 37740 38360 37792 38369
rect 38016 38360 38068 38412
rect 39028 38360 39080 38412
rect 40316 38360 40368 38412
rect 17040 38199 17092 38208
rect 17040 38165 17049 38199
rect 17049 38165 17083 38199
rect 17083 38165 17092 38199
rect 17040 38156 17092 38165
rect 17776 38156 17828 38208
rect 20720 38156 20772 38208
rect 22744 38156 22796 38208
rect 24584 38292 24636 38344
rect 26976 38292 27028 38344
rect 28356 38292 28408 38344
rect 28540 38335 28592 38344
rect 28540 38301 28549 38335
rect 28549 38301 28583 38335
rect 28583 38301 28592 38335
rect 28540 38292 28592 38301
rect 26240 38224 26292 38276
rect 30472 38224 30524 38276
rect 31208 38292 31260 38344
rect 33508 38292 33560 38344
rect 39672 38292 39724 38344
rect 43996 38335 44048 38344
rect 43996 38301 44005 38335
rect 44005 38301 44039 38335
rect 44039 38301 44048 38335
rect 43996 38292 44048 38301
rect 31576 38224 31628 38276
rect 32864 38224 32916 38276
rect 43628 38224 43680 38276
rect 46204 38292 46256 38344
rect 23940 38199 23992 38208
rect 23940 38165 23949 38199
rect 23949 38165 23983 38199
rect 23983 38165 23992 38199
rect 23940 38156 23992 38165
rect 28172 38156 28224 38208
rect 29460 38199 29512 38208
rect 29460 38165 29469 38199
rect 29469 38165 29503 38199
rect 29503 38165 29512 38199
rect 29460 38156 29512 38165
rect 31484 38199 31536 38208
rect 31484 38165 31493 38199
rect 31493 38165 31527 38199
rect 31527 38165 31536 38199
rect 31484 38156 31536 38165
rect 33048 38199 33100 38208
rect 33048 38165 33057 38199
rect 33057 38165 33091 38199
rect 33091 38165 33100 38199
rect 33048 38156 33100 38165
rect 33140 38156 33192 38208
rect 35992 38199 36044 38208
rect 35992 38165 36001 38199
rect 36001 38165 36035 38199
rect 36035 38165 36044 38199
rect 35992 38156 36044 38165
rect 40592 38156 40644 38208
rect 40868 38156 40920 38208
rect 41052 38199 41104 38208
rect 41052 38165 41061 38199
rect 41061 38165 41095 38199
rect 41095 38165 41104 38199
rect 41052 38156 41104 38165
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 15660 37952 15712 38004
rect 18052 37952 18104 38004
rect 15200 37748 15252 37800
rect 15936 37884 15988 37936
rect 16580 37927 16632 37936
rect 16580 37893 16589 37927
rect 16589 37893 16623 37927
rect 16623 37893 16632 37927
rect 16580 37884 16632 37893
rect 20168 37952 20220 38004
rect 21364 37995 21416 38004
rect 21364 37961 21373 37995
rect 21373 37961 21407 37995
rect 21407 37961 21416 37995
rect 21364 37952 21416 37961
rect 26608 37995 26660 38004
rect 26608 37961 26617 37995
rect 26617 37961 26651 37995
rect 26651 37961 26660 37995
rect 26608 37952 26660 37961
rect 26976 37995 27028 38004
rect 26976 37961 26985 37995
rect 26985 37961 27019 37995
rect 27019 37961 27028 37995
rect 26976 37952 27028 37961
rect 27068 37952 27120 38004
rect 27620 37952 27672 38004
rect 28724 37995 28776 38004
rect 28724 37961 28733 37995
rect 28733 37961 28767 37995
rect 28767 37961 28776 37995
rect 28724 37952 28776 37961
rect 18696 37884 18748 37936
rect 20904 37927 20956 37936
rect 20904 37893 20913 37927
rect 20913 37893 20947 37927
rect 20947 37893 20956 37927
rect 20904 37884 20956 37893
rect 26792 37884 26844 37936
rect 29644 37952 29696 38004
rect 30380 37995 30432 38004
rect 30380 37961 30389 37995
rect 30389 37961 30423 37995
rect 30423 37961 30432 37995
rect 30380 37952 30432 37961
rect 32128 37995 32180 38004
rect 32128 37961 32137 37995
rect 32137 37961 32171 37995
rect 32171 37961 32180 37995
rect 32128 37952 32180 37961
rect 32220 37952 32272 38004
rect 33968 37995 34020 38004
rect 33968 37961 33977 37995
rect 33977 37961 34011 37995
rect 34011 37961 34020 37995
rect 33968 37952 34020 37961
rect 35440 37952 35492 38004
rect 35532 37995 35584 38004
rect 35532 37961 35541 37995
rect 35541 37961 35575 37995
rect 35575 37961 35584 37995
rect 35532 37952 35584 37961
rect 36452 37952 36504 38004
rect 39028 37995 39080 38004
rect 39028 37961 39037 37995
rect 39037 37961 39071 37995
rect 39071 37961 39080 37995
rect 39028 37952 39080 37961
rect 40316 37995 40368 38004
rect 40316 37961 40325 37995
rect 40325 37961 40359 37995
rect 40359 37961 40368 37995
rect 40316 37952 40368 37961
rect 43904 37952 43956 38004
rect 44088 37952 44140 38004
rect 44640 37952 44692 38004
rect 44732 37927 44784 37936
rect 44732 37893 44741 37927
rect 44741 37893 44775 37927
rect 44775 37893 44784 37927
rect 44732 37884 44784 37893
rect 19432 37816 19484 37868
rect 19892 37859 19944 37868
rect 19892 37825 19901 37859
rect 19901 37825 19935 37859
rect 19935 37825 19944 37859
rect 19892 37816 19944 37825
rect 22744 37859 22796 37868
rect 22744 37825 22753 37859
rect 22753 37825 22787 37859
rect 22787 37825 22796 37859
rect 22744 37816 22796 37825
rect 28264 37859 28316 37868
rect 28264 37825 28273 37859
rect 28273 37825 28307 37859
rect 28307 37825 28316 37859
rect 28264 37816 28316 37825
rect 31484 37859 31536 37868
rect 31484 37825 31493 37859
rect 31493 37825 31527 37859
rect 31527 37825 31536 37859
rect 31484 37816 31536 37825
rect 31576 37816 31628 37868
rect 35992 37816 36044 37868
rect 40592 37816 40644 37868
rect 44180 37859 44232 37868
rect 44180 37825 44189 37859
rect 44189 37825 44223 37859
rect 44223 37825 44232 37859
rect 44180 37816 44232 37825
rect 22008 37791 22060 37800
rect 22008 37757 22017 37791
rect 22017 37757 22051 37791
rect 22051 37757 22060 37791
rect 22008 37748 22060 37757
rect 23664 37791 23716 37800
rect 15476 37680 15528 37732
rect 16120 37723 16172 37732
rect 16120 37689 16129 37723
rect 16129 37689 16163 37723
rect 16163 37689 16172 37723
rect 16120 37680 16172 37689
rect 17868 37680 17920 37732
rect 23664 37757 23673 37791
rect 23673 37757 23707 37791
rect 23707 37757 23716 37791
rect 23664 37748 23716 37757
rect 27620 37791 27672 37800
rect 27620 37757 27629 37791
rect 27629 37757 27663 37791
rect 27663 37757 27672 37791
rect 27620 37748 27672 37757
rect 28172 37791 28224 37800
rect 28172 37757 28181 37791
rect 28181 37757 28215 37791
rect 28215 37757 28224 37791
rect 28172 37748 28224 37757
rect 29184 37748 29236 37800
rect 31208 37748 31260 37800
rect 31300 37748 31352 37800
rect 31852 37748 31904 37800
rect 38292 37791 38344 37800
rect 38292 37757 38301 37791
rect 38301 37757 38335 37791
rect 38335 37757 38344 37791
rect 38292 37748 38344 37757
rect 38476 37791 38528 37800
rect 38476 37757 38485 37791
rect 38485 37757 38519 37791
rect 38519 37757 38528 37791
rect 38476 37748 38528 37757
rect 15292 37612 15344 37664
rect 17040 37612 17092 37664
rect 18052 37612 18104 37664
rect 18420 37612 18472 37664
rect 19432 37655 19484 37664
rect 19432 37621 19441 37655
rect 19441 37621 19475 37655
rect 19475 37621 19484 37655
rect 20536 37655 20588 37664
rect 19432 37612 19484 37621
rect 20536 37621 20545 37655
rect 20545 37621 20579 37655
rect 20579 37621 20588 37655
rect 20536 37612 20588 37621
rect 21824 37655 21876 37664
rect 21824 37621 21833 37655
rect 21833 37621 21867 37655
rect 21867 37621 21876 37655
rect 21824 37612 21876 37621
rect 23020 37655 23072 37664
rect 23020 37621 23029 37655
rect 23029 37621 23063 37655
rect 23063 37621 23072 37655
rect 25688 37723 25740 37732
rect 25688 37689 25697 37723
rect 25697 37689 25731 37723
rect 25731 37689 25740 37723
rect 25688 37680 25740 37689
rect 23020 37612 23072 37621
rect 23848 37612 23900 37664
rect 26148 37680 26200 37732
rect 26884 37680 26936 37732
rect 29368 37723 29420 37732
rect 29368 37689 29377 37723
rect 29377 37689 29411 37723
rect 29411 37689 29420 37723
rect 29368 37680 29420 37689
rect 29460 37723 29512 37732
rect 29460 37689 29469 37723
rect 29469 37689 29503 37723
rect 29503 37689 29512 37723
rect 32680 37723 32732 37732
rect 29460 37680 29512 37689
rect 32680 37689 32689 37723
rect 32689 37689 32723 37723
rect 32723 37689 32732 37723
rect 32680 37680 32732 37689
rect 33048 37680 33100 37732
rect 35532 37680 35584 37732
rect 36636 37680 36688 37732
rect 30564 37612 30616 37664
rect 35256 37612 35308 37664
rect 36544 37612 36596 37664
rect 37740 37680 37792 37732
rect 38936 37680 38988 37732
rect 39764 37680 39816 37732
rect 41052 37680 41104 37732
rect 41512 37723 41564 37732
rect 41512 37689 41521 37723
rect 41521 37689 41555 37723
rect 41555 37689 41564 37723
rect 41512 37680 41564 37689
rect 42432 37723 42484 37732
rect 42432 37689 42441 37723
rect 42441 37689 42475 37723
rect 42475 37689 42484 37723
rect 42432 37680 42484 37689
rect 44272 37723 44324 37732
rect 36912 37655 36964 37664
rect 36912 37621 36921 37655
rect 36921 37621 36955 37655
rect 36955 37621 36964 37655
rect 36912 37612 36964 37621
rect 39672 37655 39724 37664
rect 39672 37621 39681 37655
rect 39681 37621 39715 37655
rect 39715 37621 39724 37655
rect 39672 37612 39724 37621
rect 41880 37612 41932 37664
rect 44272 37689 44281 37723
rect 44281 37689 44315 37723
rect 44315 37689 44324 37723
rect 44272 37680 44324 37689
rect 43996 37612 44048 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 15568 37451 15620 37460
rect 15568 37417 15577 37451
rect 15577 37417 15611 37451
rect 15611 37417 15620 37451
rect 15568 37408 15620 37417
rect 18420 37408 18472 37460
rect 20904 37408 20956 37460
rect 15292 37340 15344 37392
rect 16120 37383 16172 37392
rect 16120 37349 16129 37383
rect 16129 37349 16163 37383
rect 16163 37349 16172 37383
rect 16120 37340 16172 37349
rect 17776 37383 17828 37392
rect 17776 37349 17785 37383
rect 17785 37349 17819 37383
rect 17819 37349 17828 37383
rect 17776 37340 17828 37349
rect 17960 37340 18012 37392
rect 19432 37383 19484 37392
rect 19432 37349 19441 37383
rect 19441 37349 19475 37383
rect 19475 37349 19484 37383
rect 19432 37340 19484 37349
rect 21732 37340 21784 37392
rect 23664 37408 23716 37460
rect 24952 37451 25004 37460
rect 24952 37417 24961 37451
rect 24961 37417 24995 37451
rect 24995 37417 25004 37451
rect 24952 37408 25004 37417
rect 28172 37408 28224 37460
rect 28540 37408 28592 37460
rect 29276 37408 29328 37460
rect 31300 37408 31352 37460
rect 33048 37408 33100 37460
rect 28448 37340 28500 37392
rect 33784 37340 33836 37392
rect 35992 37340 36044 37392
rect 14004 37272 14056 37324
rect 22744 37315 22796 37324
rect 22744 37281 22753 37315
rect 22753 37281 22787 37315
rect 22787 37281 22796 37315
rect 22744 37272 22796 37281
rect 23204 37315 23256 37324
rect 23204 37281 23213 37315
rect 23213 37281 23247 37315
rect 23247 37281 23256 37315
rect 23204 37272 23256 37281
rect 24676 37272 24728 37324
rect 25320 37315 25372 37324
rect 25320 37281 25329 37315
rect 25329 37281 25363 37315
rect 25363 37281 25372 37315
rect 25320 37272 25372 37281
rect 26792 37272 26844 37324
rect 29828 37315 29880 37324
rect 29828 37281 29837 37315
rect 29837 37281 29871 37315
rect 29871 37281 29880 37315
rect 29828 37272 29880 37281
rect 31024 37315 31076 37324
rect 31024 37281 31033 37315
rect 31033 37281 31067 37315
rect 31067 37281 31076 37315
rect 31024 37272 31076 37281
rect 35348 37315 35400 37324
rect 35348 37281 35357 37315
rect 35357 37281 35391 37315
rect 35391 37281 35400 37315
rect 35348 37272 35400 37281
rect 35440 37272 35492 37324
rect 36268 37272 36320 37324
rect 39120 37408 39172 37460
rect 39764 37451 39816 37460
rect 39764 37417 39773 37451
rect 39773 37417 39807 37451
rect 39807 37417 39816 37451
rect 39764 37408 39816 37417
rect 41788 37451 41840 37460
rect 41788 37417 41797 37451
rect 41797 37417 41831 37451
rect 41831 37417 41840 37451
rect 41788 37408 41840 37417
rect 42432 37451 42484 37460
rect 42432 37417 42441 37451
rect 42441 37417 42475 37451
rect 42475 37417 42484 37451
rect 42432 37408 42484 37417
rect 43996 37451 44048 37460
rect 43996 37417 44005 37451
rect 44005 37417 44039 37451
rect 44039 37417 44048 37451
rect 43996 37408 44048 37417
rect 40684 37340 40736 37392
rect 45100 37340 45152 37392
rect 37832 37272 37884 37324
rect 19340 37247 19392 37256
rect 19340 37213 19349 37247
rect 19349 37213 19383 37247
rect 19383 37213 19392 37247
rect 19340 37204 19392 37213
rect 19616 37247 19668 37256
rect 19616 37213 19625 37247
rect 19625 37213 19659 37247
rect 19659 37213 19668 37247
rect 19616 37204 19668 37213
rect 20996 37247 21048 37256
rect 20996 37213 21005 37247
rect 21005 37213 21039 37247
rect 21039 37213 21048 37247
rect 20996 37204 21048 37213
rect 21364 37247 21416 37256
rect 21364 37213 21373 37247
rect 21373 37213 21407 37247
rect 21407 37213 21416 37247
rect 21364 37204 21416 37213
rect 25688 37204 25740 37256
rect 27712 37204 27764 37256
rect 28356 37204 28408 37256
rect 32220 37247 32272 37256
rect 32220 37213 32229 37247
rect 32229 37213 32263 37247
rect 32263 37213 32272 37247
rect 32220 37204 32272 37213
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 16396 37136 16448 37188
rect 19892 37136 19944 37188
rect 25228 37136 25280 37188
rect 31116 37136 31168 37188
rect 32680 37136 32732 37188
rect 34336 37204 34388 37256
rect 38936 37204 38988 37256
rect 40592 37247 40644 37256
rect 40592 37213 40601 37247
rect 40601 37213 40635 37247
rect 40635 37213 40644 37247
rect 40592 37204 40644 37213
rect 44364 37247 44416 37256
rect 44364 37213 44373 37247
rect 44373 37213 44407 37247
rect 44407 37213 44416 37247
rect 44364 37204 44416 37213
rect 44732 37247 44784 37256
rect 44732 37213 44741 37247
rect 44741 37213 44775 37247
rect 44775 37213 44784 37247
rect 44732 37204 44784 37213
rect 45928 37247 45980 37256
rect 45928 37213 45937 37247
rect 45937 37213 45971 37247
rect 45971 37213 45980 37247
rect 45928 37204 45980 37213
rect 46204 37247 46256 37256
rect 46204 37213 46213 37247
rect 46213 37213 46247 37247
rect 46247 37213 46256 37247
rect 46204 37204 46256 37213
rect 41052 37136 41104 37188
rect 44272 37136 44324 37188
rect 15384 37068 15436 37120
rect 16028 37068 16080 37120
rect 21824 37068 21876 37120
rect 22008 37111 22060 37120
rect 22008 37077 22017 37111
rect 22017 37077 22051 37111
rect 22051 37077 22060 37111
rect 22008 37068 22060 37077
rect 24124 37111 24176 37120
rect 24124 37077 24133 37111
rect 24133 37077 24167 37111
rect 24167 37077 24176 37111
rect 24124 37068 24176 37077
rect 26332 37068 26384 37120
rect 29368 37068 29420 37120
rect 30288 37068 30340 37120
rect 30472 37111 30524 37120
rect 30472 37077 30481 37111
rect 30481 37077 30515 37111
rect 30515 37077 30524 37111
rect 30472 37068 30524 37077
rect 31300 37068 31352 37120
rect 32404 37068 32456 37120
rect 37096 37111 37148 37120
rect 37096 37077 37105 37111
rect 37105 37077 37139 37111
rect 37139 37077 37148 37111
rect 37096 37068 37148 37077
rect 38200 37068 38252 37120
rect 38476 37068 38528 37120
rect 39028 37068 39080 37120
rect 43904 37068 43956 37120
rect 45744 37068 45796 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 16120 36864 16172 36916
rect 19340 36864 19392 36916
rect 20996 36864 21048 36916
rect 22744 36864 22796 36916
rect 24676 36907 24728 36916
rect 24676 36873 24685 36907
rect 24685 36873 24719 36907
rect 24719 36873 24728 36907
rect 24676 36864 24728 36873
rect 25320 36907 25372 36916
rect 25320 36873 25329 36907
rect 25329 36873 25363 36907
rect 25363 36873 25372 36907
rect 25320 36864 25372 36873
rect 26792 36907 26844 36916
rect 26792 36873 26801 36907
rect 26801 36873 26835 36907
rect 26835 36873 26844 36907
rect 26792 36864 26844 36873
rect 28080 36864 28132 36916
rect 29828 36864 29880 36916
rect 32220 36907 32272 36916
rect 32220 36873 32229 36907
rect 32229 36873 32263 36907
rect 32263 36873 32272 36907
rect 32220 36864 32272 36873
rect 35440 36864 35492 36916
rect 36636 36907 36688 36916
rect 36636 36873 36645 36907
rect 36645 36873 36679 36907
rect 36679 36873 36688 36907
rect 36636 36864 36688 36873
rect 41144 36864 41196 36916
rect 42432 36864 42484 36916
rect 44364 36864 44416 36916
rect 17684 36796 17736 36848
rect 19432 36839 19484 36848
rect 15384 36728 15436 36780
rect 16672 36728 16724 36780
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 19432 36805 19441 36839
rect 19441 36805 19475 36839
rect 19475 36805 19484 36839
rect 19432 36796 19484 36805
rect 21824 36796 21876 36848
rect 23204 36796 23256 36848
rect 24492 36796 24544 36848
rect 19616 36728 19668 36780
rect 19892 36728 19944 36780
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 24124 36728 24176 36780
rect 24216 36771 24268 36780
rect 24216 36737 24225 36771
rect 24225 36737 24259 36771
rect 24259 36737 24268 36771
rect 24216 36728 24268 36737
rect 26148 36728 26200 36780
rect 26240 36771 26292 36780
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 26240 36728 26292 36737
rect 26884 36728 26936 36780
rect 30472 36728 30524 36780
rect 14556 36703 14608 36712
rect 14556 36669 14565 36703
rect 14565 36669 14599 36703
rect 14599 36669 14608 36703
rect 14556 36660 14608 36669
rect 22652 36660 22704 36712
rect 28080 36660 28132 36712
rect 34152 36796 34204 36848
rect 35348 36796 35400 36848
rect 37832 36796 37884 36848
rect 39120 36796 39172 36848
rect 41052 36796 41104 36848
rect 41512 36839 41564 36848
rect 41512 36805 41521 36839
rect 41521 36805 41555 36839
rect 41555 36805 41564 36839
rect 41512 36796 41564 36805
rect 45100 36796 45152 36848
rect 32680 36771 32732 36780
rect 32680 36737 32689 36771
rect 32689 36737 32723 36771
rect 32723 36737 32732 36771
rect 32680 36728 32732 36737
rect 37096 36728 37148 36780
rect 38200 36728 38252 36780
rect 42340 36728 42392 36780
rect 38568 36703 38620 36712
rect 14648 36592 14700 36644
rect 14004 36567 14056 36576
rect 14004 36533 14013 36567
rect 14013 36533 14047 36567
rect 14047 36533 14056 36567
rect 14004 36524 14056 36533
rect 16120 36524 16172 36576
rect 17960 36592 18012 36644
rect 20812 36635 20864 36644
rect 20812 36601 20821 36635
rect 20821 36601 20855 36635
rect 20855 36601 20864 36635
rect 20812 36592 20864 36601
rect 21364 36635 21416 36644
rect 21364 36601 21373 36635
rect 21373 36601 21407 36635
rect 21407 36601 21416 36635
rect 21364 36592 21416 36601
rect 21732 36635 21784 36644
rect 21732 36601 21741 36635
rect 21741 36601 21775 36635
rect 21775 36601 21784 36635
rect 21732 36592 21784 36601
rect 23940 36592 23992 36644
rect 25964 36635 26016 36644
rect 25964 36601 25973 36635
rect 25973 36601 26007 36635
rect 26007 36601 26016 36635
rect 25964 36592 26016 36601
rect 29736 36635 29788 36644
rect 29736 36601 29745 36635
rect 29745 36601 29779 36635
rect 29779 36601 29788 36635
rect 29736 36592 29788 36601
rect 16580 36524 16632 36576
rect 22652 36567 22704 36576
rect 22652 36533 22661 36567
rect 22661 36533 22695 36567
rect 22695 36533 22704 36567
rect 22652 36524 22704 36533
rect 27712 36567 27764 36576
rect 27712 36533 27721 36567
rect 27721 36533 27755 36567
rect 27755 36533 27764 36567
rect 27712 36524 27764 36533
rect 27804 36524 27856 36576
rect 28448 36524 28500 36576
rect 30932 36592 30984 36644
rect 31024 36567 31076 36576
rect 31024 36533 31033 36567
rect 31033 36533 31067 36567
rect 31067 36533 31076 36567
rect 31024 36524 31076 36533
rect 31760 36567 31812 36576
rect 31760 36533 31769 36567
rect 31769 36533 31803 36567
rect 31803 36533 31812 36567
rect 31760 36524 31812 36533
rect 32496 36635 32548 36644
rect 32496 36601 32505 36635
rect 32505 36601 32539 36635
rect 32539 36601 32548 36635
rect 32496 36592 32548 36601
rect 33600 36592 33652 36644
rect 36636 36592 36688 36644
rect 33784 36524 33836 36576
rect 35532 36567 35584 36576
rect 35532 36533 35541 36567
rect 35541 36533 35575 36567
rect 35575 36533 35584 36567
rect 35532 36524 35584 36533
rect 36268 36567 36320 36576
rect 36268 36533 36277 36567
rect 36277 36533 36311 36567
rect 36311 36533 36320 36567
rect 36268 36524 36320 36533
rect 37832 36524 37884 36576
rect 38568 36669 38577 36703
rect 38577 36669 38611 36703
rect 38611 36669 38620 36703
rect 38568 36660 38620 36669
rect 39028 36703 39080 36712
rect 39028 36669 39037 36703
rect 39037 36669 39071 36703
rect 39071 36669 39080 36703
rect 39028 36660 39080 36669
rect 40684 36703 40736 36712
rect 40684 36669 40693 36703
rect 40693 36669 40727 36703
rect 40727 36669 40736 36703
rect 40684 36660 40736 36669
rect 42524 36703 42576 36712
rect 42524 36669 42542 36703
rect 42542 36669 42576 36703
rect 42524 36660 42576 36669
rect 40592 36592 40644 36644
rect 41052 36635 41104 36644
rect 41052 36601 41061 36635
rect 41061 36601 41095 36635
rect 41095 36601 41104 36635
rect 41052 36592 41104 36601
rect 40040 36524 40092 36576
rect 44272 36592 44324 36644
rect 45192 36635 45244 36644
rect 43904 36567 43956 36576
rect 43904 36533 43913 36567
rect 43913 36533 43947 36567
rect 43947 36533 43956 36567
rect 43904 36524 43956 36533
rect 45192 36601 45201 36635
rect 45201 36601 45235 36635
rect 45235 36601 45244 36635
rect 45192 36592 45244 36601
rect 46572 36567 46624 36576
rect 46572 36533 46581 36567
rect 46581 36533 46615 36567
rect 46615 36533 46624 36567
rect 46572 36524 46624 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 15292 36320 15344 36372
rect 15476 36363 15528 36372
rect 15476 36329 15485 36363
rect 15485 36329 15519 36363
rect 15519 36329 15528 36363
rect 15476 36320 15528 36329
rect 16120 36320 16172 36372
rect 17776 36363 17828 36372
rect 17776 36329 17785 36363
rect 17785 36329 17819 36363
rect 17819 36329 17828 36363
rect 17776 36320 17828 36329
rect 19340 36320 19392 36372
rect 20720 36363 20772 36372
rect 20720 36329 20729 36363
rect 20729 36329 20763 36363
rect 20763 36329 20772 36363
rect 20720 36320 20772 36329
rect 23940 36320 23992 36372
rect 25964 36320 26016 36372
rect 14556 36252 14608 36304
rect 16488 36295 16540 36304
rect 16488 36261 16497 36295
rect 16497 36261 16531 36295
rect 16531 36261 16540 36295
rect 16488 36252 16540 36261
rect 20812 36252 20864 36304
rect 23112 36252 23164 36304
rect 23848 36252 23900 36304
rect 26332 36252 26384 36304
rect 27804 36320 27856 36372
rect 29736 36363 29788 36372
rect 29736 36329 29745 36363
rect 29745 36329 29779 36363
rect 29779 36329 29788 36363
rect 29736 36320 29788 36329
rect 26792 36252 26844 36304
rect 28540 36295 28592 36304
rect 28540 36261 28549 36295
rect 28549 36261 28583 36295
rect 28583 36261 28592 36295
rect 28540 36252 28592 36261
rect 30288 36295 30340 36304
rect 30288 36261 30297 36295
rect 30297 36261 30331 36295
rect 30331 36261 30340 36295
rect 30288 36252 30340 36261
rect 30380 36295 30432 36304
rect 30380 36261 30389 36295
rect 30389 36261 30423 36295
rect 30423 36261 30432 36295
rect 32496 36320 32548 36372
rect 33140 36320 33192 36372
rect 38936 36363 38988 36372
rect 30380 36252 30432 36261
rect 13636 36227 13688 36236
rect 13636 36193 13645 36227
rect 13645 36193 13679 36227
rect 13679 36193 13688 36227
rect 13636 36184 13688 36193
rect 14188 36227 14240 36236
rect 14188 36193 14197 36227
rect 14197 36193 14231 36227
rect 14231 36193 14240 36227
rect 14188 36184 14240 36193
rect 14924 36184 14976 36236
rect 17868 36227 17920 36236
rect 17868 36193 17877 36227
rect 17877 36193 17911 36227
rect 17911 36193 17920 36227
rect 17868 36184 17920 36193
rect 18420 36227 18472 36236
rect 18420 36193 18429 36227
rect 18429 36193 18463 36227
rect 18463 36193 18472 36227
rect 18420 36184 18472 36193
rect 20260 36184 20312 36236
rect 21732 36227 21784 36236
rect 21732 36193 21741 36227
rect 21741 36193 21775 36227
rect 21775 36193 21784 36227
rect 21732 36184 21784 36193
rect 21916 36227 21968 36236
rect 21916 36193 21925 36227
rect 21925 36193 21959 36227
rect 21959 36193 21968 36227
rect 21916 36184 21968 36193
rect 24216 36184 24268 36236
rect 24492 36184 24544 36236
rect 30932 36184 30984 36236
rect 34060 36252 34112 36304
rect 34336 36295 34388 36304
rect 34336 36261 34345 36295
rect 34345 36261 34379 36295
rect 34379 36261 34388 36295
rect 34336 36252 34388 36261
rect 37096 36252 37148 36304
rect 36544 36184 36596 36236
rect 16396 36159 16448 36168
rect 16396 36125 16405 36159
rect 16405 36125 16439 36159
rect 16439 36125 16448 36159
rect 16396 36116 16448 36125
rect 17040 36159 17092 36168
rect 17040 36125 17049 36159
rect 17049 36125 17083 36159
rect 17083 36125 17092 36159
rect 17040 36116 17092 36125
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 18788 36116 18840 36168
rect 22192 36159 22244 36168
rect 22192 36125 22201 36159
rect 22201 36125 22235 36159
rect 22235 36125 22244 36159
rect 22192 36116 22244 36125
rect 23480 36116 23532 36168
rect 26884 36159 26936 36168
rect 26884 36125 26893 36159
rect 26893 36125 26927 36159
rect 26927 36125 26936 36159
rect 26884 36116 26936 36125
rect 28908 36116 28960 36168
rect 30472 36116 30524 36168
rect 32312 36116 32364 36168
rect 33692 36159 33744 36168
rect 33692 36125 33701 36159
rect 33701 36125 33735 36159
rect 33735 36125 33744 36159
rect 33692 36116 33744 36125
rect 21732 36048 21784 36100
rect 26240 36048 26292 36100
rect 29368 36048 29420 36100
rect 31392 36048 31444 36100
rect 36728 36184 36780 36236
rect 38936 36329 38945 36363
rect 38945 36329 38979 36363
rect 38979 36329 38988 36363
rect 38936 36320 38988 36329
rect 40592 36363 40644 36372
rect 40592 36329 40601 36363
rect 40601 36329 40635 36363
rect 40635 36329 40644 36363
rect 40592 36320 40644 36329
rect 45928 36320 45980 36372
rect 46572 36320 46624 36372
rect 40868 36252 40920 36304
rect 41144 36295 41196 36304
rect 41144 36261 41153 36295
rect 41153 36261 41187 36295
rect 41187 36261 41196 36295
rect 41144 36252 41196 36261
rect 45100 36252 45152 36304
rect 38844 36184 38896 36236
rect 39028 36116 39080 36168
rect 43720 36184 43772 36236
rect 46388 36227 46440 36236
rect 46388 36193 46397 36227
rect 46397 36193 46431 36227
rect 46431 36193 46440 36227
rect 46388 36184 46440 36193
rect 39856 36159 39908 36168
rect 39856 36125 39865 36159
rect 39865 36125 39899 36159
rect 39899 36125 39908 36159
rect 39856 36116 39908 36125
rect 41512 36159 41564 36168
rect 41512 36125 41521 36159
rect 41521 36125 41555 36159
rect 41555 36125 41564 36159
rect 41512 36116 41564 36125
rect 45192 36159 45244 36168
rect 19248 36023 19300 36032
rect 19248 35989 19257 36023
rect 19257 35989 19291 36023
rect 19291 35989 19300 36023
rect 19248 35980 19300 35989
rect 21272 36023 21324 36032
rect 21272 35989 21281 36023
rect 21281 35989 21315 36023
rect 21315 35989 21324 36023
rect 21272 35980 21324 35989
rect 26148 36023 26200 36032
rect 26148 35989 26157 36023
rect 26157 35989 26191 36023
rect 26191 35989 26200 36023
rect 26148 35980 26200 35989
rect 27160 35980 27212 36032
rect 29828 35980 29880 36032
rect 32864 35980 32916 36032
rect 37096 36023 37148 36032
rect 37096 35989 37105 36023
rect 37105 35989 37139 36023
rect 37139 35989 37148 36023
rect 37096 35980 37148 35989
rect 38568 36023 38620 36032
rect 38568 35989 38577 36023
rect 38577 35989 38611 36023
rect 38611 35989 38620 36023
rect 38568 35980 38620 35989
rect 44364 35980 44416 36032
rect 45192 36125 45201 36159
rect 45201 36125 45235 36159
rect 45235 36125 45244 36159
rect 45192 36116 45244 36125
rect 45652 35980 45704 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 14648 35819 14700 35828
rect 14648 35785 14657 35819
rect 14657 35785 14691 35819
rect 14691 35785 14700 35819
rect 14648 35776 14700 35785
rect 16488 35776 16540 35828
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 18604 35819 18656 35828
rect 18604 35785 18613 35819
rect 18613 35785 18647 35819
rect 18647 35785 18656 35819
rect 18604 35776 18656 35785
rect 20260 35819 20312 35828
rect 20260 35785 20269 35819
rect 20269 35785 20303 35819
rect 20303 35785 20312 35819
rect 20260 35776 20312 35785
rect 23112 35819 23164 35828
rect 23112 35785 23121 35819
rect 23121 35785 23155 35819
rect 23155 35785 23164 35819
rect 23112 35776 23164 35785
rect 23480 35819 23532 35828
rect 23480 35785 23489 35819
rect 23489 35785 23523 35819
rect 23523 35785 23532 35819
rect 23480 35776 23532 35785
rect 24124 35776 24176 35828
rect 24492 35776 24544 35828
rect 26148 35776 26200 35828
rect 26884 35819 26936 35828
rect 26884 35785 26893 35819
rect 26893 35785 26927 35819
rect 26927 35785 26936 35819
rect 26884 35776 26936 35785
rect 13268 35708 13320 35760
rect 15752 35708 15804 35760
rect 15844 35708 15896 35760
rect 18420 35708 18472 35760
rect 21916 35708 21968 35760
rect 13268 35615 13320 35624
rect 13268 35581 13277 35615
rect 13277 35581 13311 35615
rect 13311 35581 13320 35615
rect 13268 35572 13320 35581
rect 14188 35640 14240 35692
rect 19248 35683 19300 35692
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 19984 35640 20036 35692
rect 21272 35683 21324 35692
rect 21272 35649 21281 35683
rect 21281 35649 21315 35683
rect 21315 35649 21324 35683
rect 21272 35640 21324 35649
rect 21732 35640 21784 35692
rect 13820 35572 13872 35624
rect 14740 35615 14792 35624
rect 14740 35581 14749 35615
rect 14749 35581 14783 35615
rect 14783 35581 14792 35615
rect 14740 35572 14792 35581
rect 17500 35572 17552 35624
rect 18604 35572 18656 35624
rect 24308 35708 24360 35760
rect 29736 35776 29788 35828
rect 24584 35572 24636 35624
rect 14648 35504 14700 35556
rect 14924 35436 14976 35488
rect 17500 35479 17552 35488
rect 17500 35445 17509 35479
rect 17509 35445 17543 35479
rect 17543 35445 17552 35479
rect 17500 35436 17552 35445
rect 18420 35436 18472 35488
rect 19340 35547 19392 35556
rect 19340 35513 19349 35547
rect 19349 35513 19383 35547
rect 19383 35513 19392 35547
rect 19340 35504 19392 35513
rect 20628 35504 20680 35556
rect 24032 35504 24084 35556
rect 24216 35504 24268 35556
rect 25872 35547 25924 35556
rect 25872 35513 25881 35547
rect 25881 35513 25915 35547
rect 25915 35513 25924 35547
rect 25872 35504 25924 35513
rect 25964 35547 26016 35556
rect 25964 35513 25973 35547
rect 25973 35513 26007 35547
rect 26007 35513 26016 35547
rect 25964 35504 26016 35513
rect 28540 35708 28592 35760
rect 30380 35776 30432 35828
rect 32496 35776 32548 35828
rect 33692 35776 33744 35828
rect 36636 35819 36688 35828
rect 36636 35785 36645 35819
rect 36645 35785 36679 35819
rect 36679 35785 36688 35819
rect 36636 35776 36688 35785
rect 37648 35776 37700 35828
rect 38844 35776 38896 35828
rect 40868 35776 40920 35828
rect 41144 35776 41196 35828
rect 45100 35776 45152 35828
rect 45652 35819 45704 35828
rect 45652 35785 45661 35819
rect 45661 35785 45695 35819
rect 45695 35785 45704 35819
rect 45652 35776 45704 35785
rect 30472 35708 30524 35760
rect 27804 35640 27856 35692
rect 29736 35615 29788 35624
rect 29736 35581 29745 35615
rect 29745 35581 29779 35615
rect 29779 35581 29788 35615
rect 29736 35572 29788 35581
rect 30748 35572 30800 35624
rect 18972 35436 19024 35488
rect 22836 35436 22888 35488
rect 24952 35436 25004 35488
rect 28356 35547 28408 35556
rect 28356 35513 28365 35547
rect 28365 35513 28399 35547
rect 28399 35513 28408 35547
rect 28356 35504 28408 35513
rect 32128 35708 32180 35760
rect 34060 35751 34112 35760
rect 29000 35479 29052 35488
rect 29000 35445 29009 35479
rect 29009 35445 29043 35479
rect 29043 35445 29052 35479
rect 29000 35436 29052 35445
rect 34060 35717 34069 35751
rect 34069 35717 34103 35751
rect 34103 35717 34112 35751
rect 34060 35708 34112 35717
rect 37188 35708 37240 35760
rect 38660 35751 38712 35760
rect 38660 35717 38669 35751
rect 38669 35717 38703 35751
rect 38703 35717 38712 35751
rect 38660 35708 38712 35717
rect 39488 35708 39540 35760
rect 45008 35708 45060 35760
rect 46388 35751 46440 35760
rect 46388 35717 46397 35751
rect 46397 35717 46431 35751
rect 46431 35717 46440 35751
rect 46388 35708 46440 35717
rect 37096 35640 37148 35692
rect 32864 35615 32916 35624
rect 32864 35581 32873 35615
rect 32873 35581 32907 35615
rect 32907 35581 32916 35615
rect 32864 35572 32916 35581
rect 33784 35615 33836 35624
rect 33784 35581 33793 35615
rect 33793 35581 33827 35615
rect 33827 35581 33836 35615
rect 33784 35572 33836 35581
rect 36728 35572 36780 35624
rect 38108 35572 38160 35624
rect 41512 35640 41564 35692
rect 45192 35640 45244 35692
rect 33324 35504 33376 35556
rect 36636 35504 36688 35556
rect 38016 35504 38068 35556
rect 39948 35572 40000 35624
rect 42616 35572 42668 35624
rect 43260 35615 43312 35624
rect 43260 35581 43278 35615
rect 43278 35581 43312 35615
rect 43260 35572 43312 35581
rect 40408 35504 40460 35556
rect 41788 35547 41840 35556
rect 41788 35513 41797 35547
rect 41797 35513 41831 35547
rect 41831 35513 41840 35547
rect 41788 35504 41840 35513
rect 42800 35504 42852 35556
rect 44272 35547 44324 35556
rect 44272 35513 44281 35547
rect 44281 35513 44315 35547
rect 44315 35513 44324 35547
rect 44272 35504 44324 35513
rect 44364 35547 44416 35556
rect 44364 35513 44373 35547
rect 44373 35513 44407 35547
rect 44407 35513 44416 35547
rect 44364 35504 44416 35513
rect 32128 35436 32180 35488
rect 32312 35479 32364 35488
rect 32312 35445 32321 35479
rect 32321 35445 32355 35479
rect 32355 35445 32364 35479
rect 32312 35436 32364 35445
rect 36544 35436 36596 35488
rect 38200 35436 38252 35488
rect 38568 35436 38620 35488
rect 40868 35436 40920 35488
rect 43444 35436 43496 35488
rect 43720 35479 43772 35488
rect 43720 35445 43729 35479
rect 43729 35445 43763 35479
rect 43763 35445 43772 35479
rect 43720 35436 43772 35445
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 14740 35275 14792 35284
rect 14740 35241 14749 35275
rect 14749 35241 14783 35275
rect 14783 35241 14792 35275
rect 14740 35232 14792 35241
rect 15844 35232 15896 35284
rect 16396 35232 16448 35284
rect 18880 35275 18932 35284
rect 18880 35241 18889 35275
rect 18889 35241 18923 35275
rect 18923 35241 18932 35275
rect 18880 35232 18932 35241
rect 21272 35232 21324 35284
rect 22560 35275 22612 35284
rect 22560 35241 22569 35275
rect 22569 35241 22603 35275
rect 22603 35241 22612 35275
rect 22560 35232 22612 35241
rect 16488 35207 16540 35216
rect 16488 35173 16497 35207
rect 16497 35173 16531 35207
rect 16531 35173 16540 35207
rect 16488 35164 16540 35173
rect 26332 35232 26384 35284
rect 30288 35275 30340 35284
rect 30288 35241 30297 35275
rect 30297 35241 30331 35275
rect 30331 35241 30340 35275
rect 30288 35232 30340 35241
rect 30748 35275 30800 35284
rect 30748 35241 30757 35275
rect 30757 35241 30791 35275
rect 30791 35241 30800 35275
rect 30748 35232 30800 35241
rect 32404 35275 32456 35284
rect 32404 35241 32413 35275
rect 32413 35241 32447 35275
rect 32447 35241 32456 35275
rect 32404 35232 32456 35241
rect 33324 35275 33376 35284
rect 33324 35241 33333 35275
rect 33333 35241 33367 35275
rect 33367 35241 33376 35275
rect 33324 35232 33376 35241
rect 34060 35232 34112 35284
rect 38568 35232 38620 35284
rect 44272 35232 44324 35284
rect 24124 35207 24176 35216
rect 24124 35173 24133 35207
rect 24133 35173 24167 35207
rect 24167 35173 24176 35207
rect 24124 35164 24176 35173
rect 28448 35207 28500 35216
rect 28448 35173 28457 35207
rect 28457 35173 28491 35207
rect 28491 35173 28500 35207
rect 28448 35164 28500 35173
rect 29368 35164 29420 35216
rect 35624 35164 35676 35216
rect 37096 35164 37148 35216
rect 38016 35164 38068 35216
rect 40684 35164 40736 35216
rect 43536 35207 43588 35216
rect 43536 35173 43545 35207
rect 43545 35173 43579 35207
rect 43579 35173 43588 35207
rect 43536 35164 43588 35173
rect 45100 35207 45152 35216
rect 45100 35173 45109 35207
rect 45109 35173 45143 35207
rect 45143 35173 45152 35207
rect 45100 35164 45152 35173
rect 16028 35096 16080 35148
rect 18512 35139 18564 35148
rect 18512 35105 18521 35139
rect 18521 35105 18555 35139
rect 18555 35105 18564 35139
rect 18512 35096 18564 35105
rect 22192 35139 22244 35148
rect 22192 35105 22201 35139
rect 22201 35105 22235 35139
rect 22235 35105 22244 35139
rect 22192 35096 22244 35105
rect 27252 35139 27304 35148
rect 27252 35105 27261 35139
rect 27261 35105 27295 35139
rect 27295 35105 27304 35139
rect 27252 35096 27304 35105
rect 30748 35139 30800 35148
rect 30748 35105 30757 35139
rect 30757 35105 30791 35139
rect 30791 35105 30800 35139
rect 30748 35096 30800 35105
rect 31208 35096 31260 35148
rect 32220 35096 32272 35148
rect 34152 35096 34204 35148
rect 34796 35096 34848 35148
rect 36084 35139 36136 35148
rect 16580 35028 16632 35080
rect 17040 35071 17092 35080
rect 17040 35037 17049 35071
rect 17049 35037 17083 35071
rect 17083 35037 17092 35071
rect 17040 35028 17092 35037
rect 18604 35028 18656 35080
rect 24032 35071 24084 35080
rect 24032 35037 24041 35071
rect 24041 35037 24075 35071
rect 24075 35037 24084 35071
rect 24032 35028 24084 35037
rect 24308 35071 24360 35080
rect 24308 35037 24317 35071
rect 24317 35037 24351 35071
rect 24351 35037 24360 35071
rect 24308 35028 24360 35037
rect 32956 35071 33008 35080
rect 32956 35037 32965 35071
rect 32965 35037 32999 35071
rect 32999 35037 33008 35071
rect 32956 35028 33008 35037
rect 36084 35105 36093 35139
rect 36093 35105 36127 35139
rect 36127 35105 36136 35139
rect 36084 35096 36136 35105
rect 36728 35096 36780 35148
rect 39856 35096 39908 35148
rect 46940 35096 46992 35148
rect 36176 35028 36228 35080
rect 38016 35071 38068 35080
rect 38016 35037 38025 35071
rect 38025 35037 38059 35071
rect 38059 35037 38068 35071
rect 38016 35028 38068 35037
rect 43168 35028 43220 35080
rect 43628 35028 43680 35080
rect 29828 34960 29880 35012
rect 35808 34960 35860 35012
rect 41788 35003 41840 35012
rect 41788 34969 41797 35003
rect 41797 34969 41831 35003
rect 41831 34969 41840 35003
rect 41788 34960 41840 34969
rect 42800 34960 42852 35012
rect 45192 35028 45244 35080
rect 13268 34935 13320 34944
rect 13268 34901 13277 34935
rect 13277 34901 13311 34935
rect 13311 34901 13320 34935
rect 13268 34892 13320 34901
rect 13636 34935 13688 34944
rect 13636 34901 13645 34935
rect 13645 34901 13679 34935
rect 13679 34901 13688 34935
rect 13636 34892 13688 34901
rect 17224 34892 17276 34944
rect 17868 34935 17920 34944
rect 17868 34901 17877 34935
rect 17877 34901 17911 34935
rect 17911 34901 17920 34935
rect 17868 34892 17920 34901
rect 19340 34892 19392 34944
rect 20628 34892 20680 34944
rect 25596 34935 25648 34944
rect 25596 34901 25605 34935
rect 25605 34901 25639 34935
rect 25639 34901 25648 34935
rect 25596 34892 25648 34901
rect 25872 34935 25924 34944
rect 25872 34901 25881 34935
rect 25881 34901 25915 34935
rect 25915 34901 25924 34935
rect 25872 34892 25924 34901
rect 27804 34892 27856 34944
rect 35348 34892 35400 34944
rect 37188 34935 37240 34944
rect 37188 34901 37197 34935
rect 37197 34901 37231 34935
rect 37231 34901 37240 34935
rect 37188 34892 37240 34901
rect 45376 34892 45428 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 14648 34731 14700 34740
rect 14648 34697 14657 34731
rect 14657 34697 14691 34731
rect 14691 34697 14700 34731
rect 14648 34688 14700 34697
rect 16488 34731 16540 34740
rect 16488 34697 16497 34731
rect 16497 34697 16531 34731
rect 16531 34697 16540 34731
rect 16488 34688 16540 34697
rect 16580 34688 16632 34740
rect 18512 34688 18564 34740
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 22192 34688 22244 34740
rect 22836 34688 22888 34740
rect 24124 34731 24176 34740
rect 24124 34697 24133 34731
rect 24133 34697 24167 34731
rect 24167 34697 24176 34731
rect 24124 34688 24176 34697
rect 27804 34731 27856 34740
rect 27804 34697 27813 34731
rect 27813 34697 27847 34731
rect 27847 34697 27856 34731
rect 27804 34688 27856 34697
rect 29000 34688 29052 34740
rect 29828 34731 29880 34740
rect 29828 34697 29837 34731
rect 29837 34697 29871 34731
rect 29871 34697 29880 34731
rect 29828 34688 29880 34697
rect 30748 34688 30800 34740
rect 33416 34688 33468 34740
rect 33508 34688 33560 34740
rect 36084 34731 36136 34740
rect 16028 34663 16080 34672
rect 16028 34629 16037 34663
rect 16037 34629 16071 34663
rect 16071 34629 16080 34663
rect 16028 34620 16080 34629
rect 16396 34620 16448 34672
rect 18880 34620 18932 34672
rect 21364 34663 21416 34672
rect 21364 34629 21373 34663
rect 21373 34629 21407 34663
rect 21407 34629 21416 34663
rect 21364 34620 21416 34629
rect 22560 34620 22612 34672
rect 23112 34620 23164 34672
rect 24032 34620 24084 34672
rect 27712 34620 27764 34672
rect 29552 34620 29604 34672
rect 33324 34663 33376 34672
rect 13544 34527 13596 34536
rect 13544 34493 13553 34527
rect 13553 34493 13587 34527
rect 13587 34493 13596 34527
rect 13544 34484 13596 34493
rect 13820 34527 13872 34536
rect 13820 34493 13829 34527
rect 13829 34493 13863 34527
rect 13863 34493 13872 34527
rect 13820 34484 13872 34493
rect 14832 34527 14884 34536
rect 14832 34493 14841 34527
rect 14841 34493 14875 34527
rect 14875 34493 14884 34527
rect 14832 34484 14884 34493
rect 18052 34527 18104 34536
rect 18052 34493 18061 34527
rect 18061 34493 18095 34527
rect 18095 34493 18104 34527
rect 18052 34484 18104 34493
rect 14648 34416 14700 34468
rect 18420 34552 18472 34604
rect 19432 34552 19484 34604
rect 19892 34595 19944 34604
rect 19892 34561 19901 34595
rect 19901 34561 19935 34595
rect 19935 34561 19944 34595
rect 19892 34552 19944 34561
rect 20260 34552 20312 34604
rect 27252 34595 27304 34604
rect 27252 34561 27261 34595
rect 27261 34561 27295 34595
rect 27295 34561 27304 34595
rect 27252 34552 27304 34561
rect 28448 34595 28500 34604
rect 28448 34561 28457 34595
rect 28457 34561 28491 34595
rect 28491 34561 28500 34595
rect 28448 34552 28500 34561
rect 28540 34552 28592 34604
rect 31208 34552 31260 34604
rect 33324 34629 33333 34663
rect 33333 34629 33367 34663
rect 33367 34629 33376 34663
rect 33324 34620 33376 34629
rect 36084 34697 36093 34731
rect 36093 34697 36127 34731
rect 36127 34697 36136 34731
rect 36084 34688 36136 34697
rect 37924 34688 37976 34740
rect 39856 34731 39908 34740
rect 31760 34595 31812 34604
rect 22836 34484 22888 34536
rect 23572 34527 23624 34536
rect 23572 34493 23581 34527
rect 23581 34493 23615 34527
rect 23615 34493 23624 34527
rect 23572 34484 23624 34493
rect 24308 34484 24360 34536
rect 28632 34484 28684 34536
rect 29828 34484 29880 34536
rect 31760 34561 31769 34595
rect 31769 34561 31803 34595
rect 31803 34561 31812 34595
rect 31760 34552 31812 34561
rect 32956 34552 33008 34604
rect 19340 34459 19392 34468
rect 18144 34348 18196 34400
rect 18512 34348 18564 34400
rect 19064 34391 19116 34400
rect 19064 34357 19073 34391
rect 19073 34357 19107 34391
rect 19107 34357 19116 34391
rect 19064 34348 19116 34357
rect 19340 34425 19349 34459
rect 19349 34425 19383 34459
rect 19383 34425 19392 34459
rect 19340 34416 19392 34425
rect 20812 34459 20864 34468
rect 20812 34425 20821 34459
rect 20821 34425 20855 34459
rect 20855 34425 20864 34459
rect 20812 34416 20864 34425
rect 20352 34348 20404 34400
rect 20628 34348 20680 34400
rect 25596 34459 25648 34468
rect 25596 34425 25605 34459
rect 25605 34425 25639 34459
rect 25639 34425 25648 34459
rect 25596 34416 25648 34425
rect 22560 34348 22612 34400
rect 22928 34348 22980 34400
rect 25136 34348 25188 34400
rect 26884 34416 26936 34468
rect 26700 34348 26752 34400
rect 28080 34348 28132 34400
rect 31484 34484 31536 34536
rect 32404 34484 32456 34536
rect 35624 34527 35676 34536
rect 35624 34493 35633 34527
rect 35633 34493 35667 34527
rect 35667 34493 35676 34527
rect 35624 34484 35676 34493
rect 38016 34552 38068 34604
rect 39856 34697 39865 34731
rect 39865 34697 39899 34731
rect 39899 34697 39908 34731
rect 39856 34688 39908 34697
rect 40684 34688 40736 34740
rect 43536 34731 43588 34740
rect 43536 34697 43545 34731
rect 43545 34697 43579 34731
rect 43579 34697 43588 34731
rect 43536 34688 43588 34697
rect 45192 34688 45244 34740
rect 45100 34620 45152 34672
rect 37004 34484 37056 34536
rect 37188 34484 37240 34536
rect 38660 34527 38712 34536
rect 34796 34416 34848 34468
rect 35164 34416 35216 34468
rect 38660 34493 38669 34527
rect 38669 34493 38703 34527
rect 38703 34493 38712 34527
rect 38660 34484 38712 34493
rect 38568 34416 38620 34468
rect 40408 34552 40460 34604
rect 42800 34595 42852 34604
rect 42800 34561 42809 34595
rect 42809 34561 42843 34595
rect 42843 34561 42852 34595
rect 42800 34552 42852 34561
rect 43444 34552 43496 34604
rect 44548 34552 44600 34604
rect 40684 34416 40736 34468
rect 31208 34348 31260 34400
rect 35256 34391 35308 34400
rect 35256 34357 35265 34391
rect 35265 34357 35299 34391
rect 35299 34357 35308 34391
rect 35256 34348 35308 34357
rect 36728 34348 36780 34400
rect 44824 34484 44876 34536
rect 42524 34459 42576 34468
rect 42524 34425 42533 34459
rect 42533 34425 42567 34459
rect 42567 34425 42576 34459
rect 42524 34416 42576 34425
rect 43812 34416 43864 34468
rect 44364 34416 44416 34468
rect 44732 34459 44784 34468
rect 44732 34425 44741 34459
rect 44741 34425 44775 34459
rect 44775 34425 44784 34459
rect 44732 34416 44784 34425
rect 44272 34348 44324 34400
rect 45100 34348 45152 34400
rect 46940 34391 46992 34400
rect 46940 34357 46949 34391
rect 46949 34357 46983 34391
rect 46983 34357 46992 34391
rect 46940 34348 46992 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 13360 34187 13412 34196
rect 13360 34153 13369 34187
rect 13369 34153 13403 34187
rect 13403 34153 13412 34187
rect 13360 34144 13412 34153
rect 13544 34144 13596 34196
rect 14832 34187 14884 34196
rect 14832 34153 14841 34187
rect 14841 34153 14875 34187
rect 14875 34153 14884 34187
rect 14832 34144 14884 34153
rect 15660 34144 15712 34196
rect 16396 34187 16448 34196
rect 16396 34153 16405 34187
rect 16405 34153 16439 34187
rect 16439 34153 16448 34187
rect 16396 34144 16448 34153
rect 18052 34144 18104 34196
rect 19064 34144 19116 34196
rect 19340 34144 19392 34196
rect 19432 34144 19484 34196
rect 20812 34144 20864 34196
rect 22928 34144 22980 34196
rect 24124 34144 24176 34196
rect 32404 34144 32456 34196
rect 35624 34144 35676 34196
rect 36728 34187 36780 34196
rect 36728 34153 36737 34187
rect 36737 34153 36771 34187
rect 36771 34153 36780 34187
rect 36728 34144 36780 34153
rect 38016 34187 38068 34196
rect 38016 34153 38025 34187
rect 38025 34153 38059 34187
rect 38059 34153 38068 34187
rect 38016 34144 38068 34153
rect 38200 34144 38252 34196
rect 42524 34187 42576 34196
rect 17684 34119 17736 34128
rect 17684 34085 17693 34119
rect 17693 34085 17727 34119
rect 17727 34085 17736 34119
rect 17684 34076 17736 34085
rect 17960 34119 18012 34128
rect 17960 34085 17969 34119
rect 17969 34085 18003 34119
rect 18003 34085 18012 34119
rect 17960 34076 18012 34085
rect 18604 34076 18656 34128
rect 16028 33983 16080 33992
rect 16028 33949 16037 33983
rect 16037 33949 16071 33983
rect 16071 33949 16080 33983
rect 16028 33940 16080 33949
rect 20168 34008 20220 34060
rect 20720 34008 20772 34060
rect 22744 34051 22796 34060
rect 22744 34017 22753 34051
rect 22753 34017 22787 34051
rect 22787 34017 22796 34051
rect 22744 34008 22796 34017
rect 23204 34051 23256 34060
rect 23204 34017 23213 34051
rect 23213 34017 23247 34051
rect 23247 34017 23256 34051
rect 23204 34008 23256 34017
rect 23296 33983 23348 33992
rect 23296 33949 23305 33983
rect 23305 33949 23339 33983
rect 23339 33949 23348 33983
rect 23296 33940 23348 33949
rect 25136 34076 25188 34128
rect 26608 34076 26660 34128
rect 29736 34076 29788 34128
rect 32220 34051 32272 34060
rect 32220 34017 32229 34051
rect 32229 34017 32263 34051
rect 32263 34017 32272 34051
rect 32220 34008 32272 34017
rect 32864 34119 32916 34128
rect 32864 34085 32873 34119
rect 32873 34085 32907 34119
rect 32907 34085 32916 34119
rect 32864 34076 32916 34085
rect 35348 34076 35400 34128
rect 36452 34076 36504 34128
rect 38660 34076 38712 34128
rect 40408 34076 40460 34128
rect 40684 34119 40736 34128
rect 40684 34085 40693 34119
rect 40693 34085 40727 34119
rect 40727 34085 40736 34119
rect 40684 34076 40736 34085
rect 40868 34076 40920 34128
rect 42524 34153 42533 34187
rect 42533 34153 42567 34187
rect 42567 34153 42576 34187
rect 42524 34144 42576 34153
rect 44272 34144 44324 34196
rect 44548 34144 44600 34196
rect 41420 34076 41472 34128
rect 43168 34119 43220 34128
rect 43168 34085 43177 34119
rect 43177 34085 43211 34119
rect 43211 34085 43220 34119
rect 43168 34076 43220 34085
rect 43812 34119 43864 34128
rect 43812 34085 43821 34119
rect 43821 34085 43855 34119
rect 43855 34085 43864 34119
rect 43812 34076 43864 34085
rect 34612 34008 34664 34060
rect 37464 34008 37516 34060
rect 38476 34008 38528 34060
rect 38568 34051 38620 34060
rect 38568 34017 38577 34051
rect 38577 34017 38611 34051
rect 38611 34017 38620 34051
rect 39856 34051 39908 34060
rect 38568 34008 38620 34017
rect 39856 34017 39865 34051
rect 39865 34017 39899 34051
rect 39899 34017 39908 34051
rect 39856 34008 39908 34017
rect 45376 34008 45428 34060
rect 24676 33983 24728 33992
rect 24676 33949 24685 33983
rect 24685 33949 24719 33983
rect 24719 33949 24728 33983
rect 24676 33940 24728 33949
rect 24768 33940 24820 33992
rect 26700 33940 26752 33992
rect 26884 33983 26936 33992
rect 26884 33949 26893 33983
rect 26893 33949 26927 33983
rect 26927 33949 26936 33983
rect 26884 33940 26936 33949
rect 28172 33983 28224 33992
rect 28172 33949 28181 33983
rect 28181 33949 28215 33983
rect 28215 33949 28224 33983
rect 28172 33940 28224 33949
rect 31208 33940 31260 33992
rect 33876 33983 33928 33992
rect 33876 33949 33885 33983
rect 33885 33949 33919 33983
rect 33919 33949 33928 33983
rect 33876 33940 33928 33949
rect 29092 33872 29144 33924
rect 32956 33872 33008 33924
rect 34704 33872 34756 33924
rect 19800 33804 19852 33856
rect 21916 33804 21968 33856
rect 27528 33847 27580 33856
rect 27528 33813 27537 33847
rect 27537 33813 27571 33847
rect 27571 33813 27580 33847
rect 27528 33804 27580 33813
rect 31116 33847 31168 33856
rect 31116 33813 31125 33847
rect 31125 33813 31159 33847
rect 31159 33813 31168 33847
rect 31116 33804 31168 33813
rect 32404 33804 32456 33856
rect 34152 33847 34204 33856
rect 34152 33813 34161 33847
rect 34161 33813 34195 33847
rect 34195 33813 34204 33847
rect 34152 33804 34204 33813
rect 35164 33940 35216 33992
rect 35808 33940 35860 33992
rect 41512 33983 41564 33992
rect 41512 33949 41521 33983
rect 41521 33949 41555 33983
rect 41555 33949 41564 33983
rect 41512 33940 41564 33949
rect 44088 33940 44140 33992
rect 45100 33940 45152 33992
rect 35256 33915 35308 33924
rect 35256 33881 35265 33915
rect 35265 33881 35299 33915
rect 35299 33881 35308 33915
rect 35256 33872 35308 33881
rect 36728 33872 36780 33924
rect 43168 33872 43220 33924
rect 35624 33804 35676 33856
rect 40500 33804 40552 33856
rect 43628 33804 43680 33856
rect 44824 33804 44876 33856
rect 46020 33804 46072 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 14648 33600 14700 33652
rect 16396 33600 16448 33652
rect 17500 33643 17552 33652
rect 17500 33609 17509 33643
rect 17509 33609 17543 33643
rect 17543 33609 17552 33643
rect 17500 33600 17552 33609
rect 19432 33600 19484 33652
rect 20168 33600 20220 33652
rect 22744 33643 22796 33652
rect 22744 33609 22753 33643
rect 22753 33609 22787 33643
rect 22787 33609 22796 33643
rect 22744 33600 22796 33609
rect 23204 33643 23256 33652
rect 23204 33609 23213 33643
rect 23213 33609 23247 33643
rect 23247 33609 23256 33643
rect 23204 33600 23256 33609
rect 24676 33600 24728 33652
rect 25872 33600 25924 33652
rect 28172 33643 28224 33652
rect 28172 33609 28181 33643
rect 28181 33609 28215 33643
rect 28215 33609 28224 33643
rect 28172 33600 28224 33609
rect 31300 33643 31352 33652
rect 13820 33532 13872 33584
rect 24584 33532 24636 33584
rect 24860 33532 24912 33584
rect 29644 33532 29696 33584
rect 31300 33609 31309 33643
rect 31309 33609 31343 33643
rect 31343 33609 31352 33643
rect 31300 33600 31352 33609
rect 32404 33600 32456 33652
rect 35256 33600 35308 33652
rect 35532 33643 35584 33652
rect 35532 33609 35541 33643
rect 35541 33609 35575 33643
rect 35575 33609 35584 33643
rect 35532 33600 35584 33609
rect 36360 33600 36412 33652
rect 36728 33643 36780 33652
rect 36728 33609 36737 33643
rect 36737 33609 36771 33643
rect 36771 33609 36780 33643
rect 36728 33600 36780 33609
rect 36912 33643 36964 33652
rect 36912 33609 36921 33643
rect 36921 33609 36955 33643
rect 36955 33609 36964 33643
rect 36912 33600 36964 33609
rect 38476 33643 38528 33652
rect 38476 33609 38485 33643
rect 38485 33609 38519 33643
rect 38519 33609 38528 33643
rect 38476 33600 38528 33609
rect 40040 33600 40092 33652
rect 40868 33600 40920 33652
rect 35624 33532 35676 33584
rect 38568 33532 38620 33584
rect 39396 33532 39448 33584
rect 41236 33575 41288 33584
rect 16028 33507 16080 33516
rect 14740 33396 14792 33448
rect 15292 33396 15344 33448
rect 15660 33396 15712 33448
rect 16028 33473 16037 33507
rect 16037 33473 16071 33507
rect 16071 33473 16080 33507
rect 16028 33464 16080 33473
rect 18052 33464 18104 33516
rect 20076 33464 20128 33516
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 24768 33507 24820 33516
rect 24768 33473 24777 33507
rect 24777 33473 24811 33507
rect 24811 33473 24820 33507
rect 24768 33464 24820 33473
rect 26792 33507 26844 33516
rect 26792 33473 26801 33507
rect 26801 33473 26835 33507
rect 26835 33473 26844 33507
rect 26792 33464 26844 33473
rect 27528 33464 27580 33516
rect 31116 33464 31168 33516
rect 32312 33464 32364 33516
rect 35808 33464 35860 33516
rect 36820 33507 36872 33516
rect 36820 33473 36829 33507
rect 36829 33473 36863 33507
rect 36863 33473 36872 33507
rect 36820 33464 36872 33473
rect 39212 33464 39264 33516
rect 39856 33464 39908 33516
rect 17500 33396 17552 33448
rect 18604 33439 18656 33448
rect 18604 33405 18613 33439
rect 18613 33405 18647 33439
rect 18647 33405 18656 33439
rect 18604 33396 18656 33405
rect 16856 33328 16908 33380
rect 19800 33396 19852 33448
rect 21916 33439 21968 33448
rect 19064 33371 19116 33380
rect 19064 33337 19073 33371
rect 19073 33337 19107 33371
rect 19107 33337 19116 33371
rect 19064 33328 19116 33337
rect 17316 33260 17368 33312
rect 20076 33371 20128 33380
rect 20076 33337 20085 33371
rect 20085 33337 20119 33371
rect 20119 33337 20128 33371
rect 20076 33328 20128 33337
rect 21364 33328 21416 33380
rect 21916 33405 21925 33439
rect 21925 33405 21959 33439
rect 21959 33405 21968 33439
rect 21916 33396 21968 33405
rect 22376 33396 22428 33448
rect 26056 33439 26108 33448
rect 26056 33405 26065 33439
rect 26065 33405 26099 33439
rect 26099 33405 26108 33439
rect 26056 33396 26108 33405
rect 29736 33439 29788 33448
rect 29736 33405 29745 33439
rect 29745 33405 29779 33439
rect 29779 33405 29788 33439
rect 29736 33396 29788 33405
rect 31392 33396 31444 33448
rect 32220 33396 32272 33448
rect 34336 33396 34388 33448
rect 37280 33396 37332 33448
rect 40040 33396 40092 33448
rect 41236 33541 41245 33575
rect 41245 33541 41279 33575
rect 41279 33541 41288 33575
rect 41236 33532 41288 33541
rect 41420 33532 41472 33584
rect 43812 33600 43864 33652
rect 44088 33643 44140 33652
rect 44088 33609 44097 33643
rect 44097 33609 44131 33643
rect 44131 33609 44140 33643
rect 44088 33600 44140 33609
rect 45008 33643 45060 33652
rect 45008 33609 45017 33643
rect 45017 33609 45051 33643
rect 45051 33609 45060 33643
rect 45008 33600 45060 33609
rect 45376 33600 45428 33652
rect 22008 33328 22060 33380
rect 22836 33328 22888 33380
rect 24124 33328 24176 33380
rect 26608 33328 26660 33380
rect 27436 33371 27488 33380
rect 20260 33260 20312 33312
rect 20720 33260 20772 33312
rect 21732 33303 21784 33312
rect 21732 33269 21741 33303
rect 21741 33269 21775 33303
rect 21775 33269 21784 33303
rect 21732 33260 21784 33269
rect 25136 33303 25188 33312
rect 25136 33269 25145 33303
rect 25145 33269 25179 33303
rect 25179 33269 25188 33303
rect 25136 33260 25188 33269
rect 27436 33337 27445 33371
rect 27445 33337 27479 33371
rect 27479 33337 27488 33371
rect 27436 33328 27488 33337
rect 29828 33328 29880 33380
rect 30472 33328 30524 33380
rect 31760 33371 31812 33380
rect 31760 33337 31769 33371
rect 31769 33337 31803 33371
rect 31803 33337 31812 33371
rect 31760 33328 31812 33337
rect 33968 33371 34020 33380
rect 33968 33337 33977 33371
rect 33977 33337 34011 33371
rect 34011 33337 34020 33371
rect 33968 33328 34020 33337
rect 34612 33371 34664 33380
rect 34612 33337 34621 33371
rect 34621 33337 34655 33371
rect 34655 33337 34664 33371
rect 34612 33328 34664 33337
rect 34704 33328 34756 33380
rect 35256 33328 35308 33380
rect 36452 33371 36504 33380
rect 36452 33337 36461 33371
rect 36461 33337 36495 33371
rect 36495 33337 36504 33371
rect 36452 33328 36504 33337
rect 40592 33328 40644 33380
rect 42984 33396 43036 33448
rect 46940 33464 46992 33516
rect 45008 33396 45060 33448
rect 43628 33328 43680 33380
rect 38200 33303 38252 33312
rect 38200 33269 38209 33303
rect 38209 33269 38243 33303
rect 38243 33269 38252 33303
rect 38200 33260 38252 33269
rect 40960 33260 41012 33312
rect 42156 33260 42208 33312
rect 43168 33260 43220 33312
rect 44732 33260 44784 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 17960 33099 18012 33108
rect 17960 33065 17969 33099
rect 17969 33065 18003 33099
rect 18003 33065 18012 33099
rect 17960 33056 18012 33065
rect 20812 33056 20864 33108
rect 22652 33056 22704 33108
rect 13820 32988 13872 33040
rect 15384 33031 15436 33040
rect 15384 32997 15393 33031
rect 15393 32997 15427 33031
rect 15427 32997 15436 33031
rect 15384 32988 15436 32997
rect 15568 32988 15620 33040
rect 13636 32963 13688 32972
rect 13636 32929 13645 32963
rect 13645 32929 13679 32963
rect 13679 32929 13688 32963
rect 13636 32920 13688 32929
rect 13912 32920 13964 32972
rect 17224 32988 17276 33040
rect 19340 33031 19392 33040
rect 19340 32997 19349 33031
rect 19349 32997 19383 33031
rect 19383 32997 19392 33031
rect 19340 32988 19392 32997
rect 21088 33031 21140 33040
rect 21088 32997 21097 33031
rect 21097 32997 21131 33031
rect 21131 32997 21140 33031
rect 21088 32988 21140 32997
rect 23112 32988 23164 33040
rect 24124 33099 24176 33108
rect 24124 33065 24133 33099
rect 24133 33065 24167 33099
rect 24167 33065 24176 33099
rect 24124 33056 24176 33065
rect 26608 33056 26660 33108
rect 29644 33099 29696 33108
rect 29644 33065 29653 33099
rect 29653 33065 29687 33099
rect 29687 33065 29696 33099
rect 29644 33056 29696 33065
rect 29736 33056 29788 33108
rect 35440 33056 35492 33108
rect 36544 33056 36596 33108
rect 38108 33056 38160 33108
rect 38936 33056 38988 33108
rect 25136 32988 25188 33040
rect 27068 32988 27120 33040
rect 28632 33031 28684 33040
rect 28632 32997 28641 33031
rect 28641 32997 28675 33031
rect 28675 32997 28684 33031
rect 28632 32988 28684 32997
rect 32956 32988 33008 33040
rect 41052 33031 41104 33040
rect 41052 32997 41061 33031
rect 41061 32997 41095 33031
rect 41095 32997 41104 33031
rect 41052 32988 41104 32997
rect 44824 33031 44876 33040
rect 44824 32997 44833 33031
rect 44833 32997 44867 33031
rect 44867 32997 44876 33031
rect 44824 32988 44876 32997
rect 17132 32920 17184 32972
rect 18144 32920 18196 32972
rect 14372 32895 14424 32904
rect 14372 32861 14381 32895
rect 14381 32861 14415 32895
rect 14415 32861 14424 32895
rect 14372 32852 14424 32861
rect 15844 32895 15896 32904
rect 15844 32861 15853 32895
rect 15853 32861 15887 32895
rect 15887 32861 15896 32895
rect 15844 32852 15896 32861
rect 18052 32852 18104 32904
rect 19064 32895 19116 32904
rect 19064 32861 19073 32895
rect 19073 32861 19107 32895
rect 19107 32861 19116 32895
rect 19064 32852 19116 32861
rect 19892 32920 19944 32972
rect 20076 32920 20128 32972
rect 23296 32920 23348 32972
rect 25320 32920 25372 32972
rect 30288 32963 30340 32972
rect 30288 32929 30297 32963
rect 30297 32929 30331 32963
rect 30331 32929 30340 32963
rect 30288 32920 30340 32929
rect 30564 32963 30616 32972
rect 30564 32929 30573 32963
rect 30573 32929 30607 32963
rect 30607 32929 30616 32963
rect 30564 32920 30616 32929
rect 32312 32920 32364 32972
rect 34244 32963 34296 32972
rect 22652 32852 22704 32904
rect 21640 32784 21692 32836
rect 27436 32852 27488 32904
rect 27712 32852 27764 32904
rect 28540 32895 28592 32904
rect 28540 32861 28549 32895
rect 28549 32861 28583 32895
rect 28583 32861 28592 32895
rect 28540 32852 28592 32861
rect 32496 32895 32548 32904
rect 32496 32861 32505 32895
rect 32505 32861 32539 32895
rect 32539 32861 32548 32895
rect 32496 32852 32548 32861
rect 32588 32895 32640 32904
rect 32588 32861 32597 32895
rect 32597 32861 32631 32895
rect 32631 32861 32640 32895
rect 32588 32852 32640 32861
rect 29092 32827 29144 32836
rect 29092 32793 29101 32827
rect 29101 32793 29135 32827
rect 29135 32793 29144 32827
rect 29092 32784 29144 32793
rect 31116 32784 31168 32836
rect 31852 32784 31904 32836
rect 33692 32784 33744 32836
rect 34244 32929 34253 32963
rect 34253 32929 34287 32963
rect 34287 32929 34296 32963
rect 34244 32920 34296 32929
rect 35256 32963 35308 32972
rect 35256 32929 35265 32963
rect 35265 32929 35299 32963
rect 35299 32929 35308 32963
rect 35256 32920 35308 32929
rect 35440 32920 35492 32972
rect 36084 32920 36136 32972
rect 37464 32920 37516 32972
rect 38200 32963 38252 32972
rect 38200 32929 38209 32963
rect 38209 32929 38243 32963
rect 38243 32929 38252 32963
rect 38200 32920 38252 32929
rect 39764 32920 39816 32972
rect 43812 32920 43864 32972
rect 45744 32920 45796 32972
rect 35716 32852 35768 32904
rect 38108 32852 38160 32904
rect 40316 32852 40368 32904
rect 41880 32852 41932 32904
rect 44732 32895 44784 32904
rect 44732 32861 44741 32895
rect 44741 32861 44775 32895
rect 44775 32861 44784 32895
rect 44732 32852 44784 32861
rect 45008 32895 45060 32904
rect 45008 32861 45017 32895
rect 45017 32861 45051 32895
rect 45051 32861 45060 32895
rect 45008 32852 45060 32861
rect 18604 32716 18656 32768
rect 19248 32716 19300 32768
rect 20260 32759 20312 32768
rect 20260 32725 20269 32759
rect 20269 32725 20303 32759
rect 20303 32725 20312 32759
rect 20260 32716 20312 32725
rect 20628 32716 20680 32768
rect 25412 32716 25464 32768
rect 26148 32716 26200 32768
rect 27528 32759 27580 32768
rect 27528 32725 27537 32759
rect 27537 32725 27571 32759
rect 27571 32725 27580 32759
rect 27528 32716 27580 32725
rect 31944 32759 31996 32768
rect 31944 32725 31953 32759
rect 31953 32725 31987 32759
rect 31987 32725 31996 32759
rect 31944 32716 31996 32725
rect 32404 32759 32456 32768
rect 32404 32725 32413 32759
rect 32413 32725 32447 32759
rect 32447 32725 32456 32759
rect 32404 32716 32456 32725
rect 33600 32716 33652 32768
rect 33784 32759 33836 32768
rect 33784 32725 33793 32759
rect 33793 32725 33827 32759
rect 33827 32725 33836 32759
rect 33784 32716 33836 32725
rect 33968 32784 34020 32836
rect 35808 32784 35860 32836
rect 36360 32784 36412 32836
rect 34704 32716 34756 32768
rect 35900 32759 35952 32768
rect 35900 32725 35909 32759
rect 35909 32725 35943 32759
rect 35943 32725 35952 32759
rect 35900 32716 35952 32725
rect 38016 32716 38068 32768
rect 44456 32716 44508 32768
rect 45836 32716 45888 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 13820 32512 13872 32564
rect 13820 32376 13872 32428
rect 13544 32308 13596 32360
rect 14004 32512 14056 32564
rect 14556 32512 14608 32564
rect 15384 32512 15436 32564
rect 16856 32555 16908 32564
rect 16856 32521 16865 32555
rect 16865 32521 16899 32555
rect 16899 32521 16908 32555
rect 16856 32512 16908 32521
rect 17224 32512 17276 32564
rect 19064 32512 19116 32564
rect 22652 32555 22704 32564
rect 22652 32521 22661 32555
rect 22661 32521 22695 32555
rect 22695 32521 22704 32555
rect 22652 32512 22704 32521
rect 23296 32512 23348 32564
rect 24584 32512 24636 32564
rect 26148 32555 26200 32564
rect 26148 32521 26157 32555
rect 26157 32521 26191 32555
rect 26191 32521 26200 32555
rect 26148 32512 26200 32521
rect 26792 32512 26844 32564
rect 27068 32512 27120 32564
rect 15568 32487 15620 32496
rect 15568 32453 15577 32487
rect 15577 32453 15611 32487
rect 15611 32453 15620 32487
rect 15568 32444 15620 32453
rect 16396 32444 16448 32496
rect 14372 32419 14424 32428
rect 14372 32385 14381 32419
rect 14381 32385 14415 32419
rect 14415 32385 14424 32419
rect 14372 32376 14424 32385
rect 16856 32308 16908 32360
rect 14556 32240 14608 32292
rect 20536 32444 20588 32496
rect 20720 32444 20772 32496
rect 25320 32444 25372 32496
rect 28632 32444 28684 32496
rect 18052 32419 18104 32428
rect 18052 32385 18061 32419
rect 18061 32385 18095 32419
rect 18095 32385 18104 32419
rect 18052 32376 18104 32385
rect 24492 32419 24544 32428
rect 24492 32385 24501 32419
rect 24501 32385 24535 32419
rect 24535 32385 24544 32419
rect 24492 32376 24544 32385
rect 24768 32419 24820 32428
rect 24768 32385 24777 32419
rect 24777 32385 24811 32419
rect 24811 32385 24820 32419
rect 24768 32376 24820 32385
rect 20352 32308 20404 32360
rect 20536 32351 20588 32360
rect 20536 32317 20545 32351
rect 20545 32317 20579 32351
rect 20579 32317 20588 32351
rect 20536 32308 20588 32317
rect 21732 32308 21784 32360
rect 21916 32308 21968 32360
rect 25412 32308 25464 32360
rect 29276 32351 29328 32360
rect 19340 32240 19392 32292
rect 23112 32240 23164 32292
rect 24584 32283 24636 32292
rect 24584 32249 24593 32283
rect 24593 32249 24627 32283
rect 24627 32249 24636 32283
rect 24584 32240 24636 32249
rect 13636 32172 13688 32224
rect 16396 32215 16448 32224
rect 16396 32181 16405 32215
rect 16405 32181 16439 32215
rect 16439 32181 16448 32215
rect 17132 32215 17184 32224
rect 16396 32172 16448 32181
rect 17132 32181 17141 32215
rect 17141 32181 17175 32215
rect 17175 32181 17184 32215
rect 17132 32172 17184 32181
rect 18972 32215 19024 32224
rect 18972 32181 18981 32215
rect 18981 32181 19015 32215
rect 19015 32181 19024 32215
rect 18972 32172 19024 32181
rect 20444 32172 20496 32224
rect 21088 32172 21140 32224
rect 29276 32317 29285 32351
rect 29285 32317 29319 32351
rect 29319 32317 29328 32351
rect 29276 32308 29328 32317
rect 31668 32308 31720 32360
rect 31852 32444 31904 32496
rect 32128 32487 32180 32496
rect 32128 32453 32137 32487
rect 32137 32453 32171 32487
rect 32171 32453 32180 32487
rect 32128 32444 32180 32453
rect 33140 32512 33192 32564
rect 34244 32512 34296 32564
rect 34704 32555 34756 32564
rect 34704 32521 34713 32555
rect 34713 32521 34747 32555
rect 34747 32521 34756 32555
rect 34704 32512 34756 32521
rect 35440 32512 35492 32564
rect 36268 32512 36320 32564
rect 37464 32555 37516 32564
rect 37464 32521 37473 32555
rect 37473 32521 37507 32555
rect 37507 32521 37516 32555
rect 37464 32512 37516 32521
rect 38200 32512 38252 32564
rect 40316 32555 40368 32564
rect 40316 32521 40325 32555
rect 40325 32521 40359 32555
rect 40359 32521 40368 32555
rect 40316 32512 40368 32521
rect 41052 32512 41104 32564
rect 32956 32487 33008 32496
rect 32956 32453 32965 32487
rect 32965 32453 32999 32487
rect 32999 32453 33008 32487
rect 32956 32444 33008 32453
rect 33876 32419 33928 32428
rect 31944 32308 31996 32360
rect 33876 32385 33885 32419
rect 33885 32385 33919 32419
rect 33919 32385 33928 32419
rect 33876 32376 33928 32385
rect 33600 32351 33652 32360
rect 33600 32317 33609 32351
rect 33609 32317 33643 32351
rect 33643 32317 33652 32351
rect 33600 32308 33652 32317
rect 34612 32444 34664 32496
rect 35716 32444 35768 32496
rect 35348 32376 35400 32428
rect 27436 32283 27488 32292
rect 27436 32249 27445 32283
rect 27445 32249 27479 32283
rect 27479 32249 27488 32283
rect 27436 32240 27488 32249
rect 27528 32283 27580 32292
rect 27528 32249 27537 32283
rect 27537 32249 27571 32283
rect 27571 32249 27580 32283
rect 27528 32240 27580 32249
rect 27712 32240 27764 32292
rect 28448 32240 28500 32292
rect 27068 32172 27120 32224
rect 28632 32172 28684 32224
rect 28724 32172 28776 32224
rect 29828 32240 29880 32292
rect 34796 32308 34848 32360
rect 35992 32308 36044 32360
rect 34888 32283 34940 32292
rect 34888 32249 34897 32283
rect 34897 32249 34931 32283
rect 34931 32249 34940 32283
rect 36544 32376 36596 32428
rect 38016 32419 38068 32428
rect 38016 32385 38025 32419
rect 38025 32385 38059 32419
rect 38059 32385 38068 32419
rect 38016 32376 38068 32385
rect 40960 32376 41012 32428
rect 42156 32376 42208 32428
rect 42892 32376 42944 32428
rect 36268 32283 36320 32292
rect 34888 32240 34940 32249
rect 36268 32249 36277 32283
rect 36277 32249 36311 32283
rect 36311 32249 36320 32283
rect 36636 32308 36688 32360
rect 36912 32308 36964 32360
rect 38200 32308 38252 32360
rect 41788 32351 41840 32360
rect 41788 32317 41797 32351
rect 41797 32317 41831 32351
rect 41831 32317 41840 32351
rect 41788 32308 41840 32317
rect 36268 32240 36320 32249
rect 38660 32240 38712 32292
rect 41144 32240 41196 32292
rect 42892 32283 42944 32292
rect 42892 32249 42901 32283
rect 42901 32249 42935 32283
rect 42935 32249 42944 32283
rect 42892 32240 42944 32249
rect 44456 32419 44508 32428
rect 44456 32385 44465 32419
rect 44465 32385 44499 32419
rect 44499 32385 44508 32419
rect 44456 32376 44508 32385
rect 46664 32376 46716 32428
rect 45560 32308 45612 32360
rect 30656 32215 30708 32224
rect 30656 32181 30665 32215
rect 30665 32181 30699 32215
rect 30699 32181 30708 32215
rect 30656 32172 30708 32181
rect 32404 32172 32456 32224
rect 35440 32172 35492 32224
rect 37924 32172 37976 32224
rect 39764 32172 39816 32224
rect 42616 32215 42668 32224
rect 42616 32181 42625 32215
rect 42625 32181 42659 32215
rect 42659 32181 42668 32215
rect 44824 32240 44876 32292
rect 43812 32215 43864 32224
rect 42616 32172 42668 32181
rect 43812 32181 43821 32215
rect 43821 32181 43855 32215
rect 43855 32181 43864 32215
rect 43812 32172 43864 32181
rect 45192 32172 45244 32224
rect 46848 32283 46900 32292
rect 46848 32249 46857 32283
rect 46857 32249 46891 32283
rect 46891 32249 46900 32283
rect 46848 32240 46900 32249
rect 45744 32172 45796 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 14372 31968 14424 32020
rect 14740 31968 14792 32020
rect 15568 31900 15620 31952
rect 18052 31943 18104 31952
rect 18052 31909 18061 31943
rect 18061 31909 18095 31943
rect 18095 31909 18104 31943
rect 18052 31900 18104 31909
rect 18972 31900 19024 31952
rect 16856 31875 16908 31884
rect 16856 31841 16865 31875
rect 16865 31841 16899 31875
rect 16899 31841 16908 31875
rect 16856 31832 16908 31841
rect 13728 31807 13780 31816
rect 13728 31773 13737 31807
rect 13737 31773 13771 31807
rect 13771 31773 13780 31807
rect 13728 31764 13780 31773
rect 14372 31807 14424 31816
rect 14372 31773 14381 31807
rect 14381 31773 14415 31807
rect 14415 31773 14424 31807
rect 14372 31764 14424 31773
rect 15384 31807 15436 31816
rect 15384 31773 15393 31807
rect 15393 31773 15427 31807
rect 15427 31773 15436 31807
rect 15384 31764 15436 31773
rect 17684 31764 17736 31816
rect 18236 31807 18288 31816
rect 18236 31773 18245 31807
rect 18245 31773 18279 31807
rect 18279 31773 18288 31807
rect 18236 31764 18288 31773
rect 18880 31764 18932 31816
rect 20260 31968 20312 32020
rect 21916 32011 21968 32020
rect 21916 31977 21925 32011
rect 21925 31977 21959 32011
rect 21959 31977 21968 32011
rect 21916 31968 21968 31977
rect 27436 31968 27488 32020
rect 29276 32011 29328 32020
rect 29276 31977 29285 32011
rect 29285 31977 29319 32011
rect 29319 31977 29328 32011
rect 29276 31968 29328 31977
rect 30564 32011 30616 32020
rect 30564 31977 30573 32011
rect 30573 31977 30607 32011
rect 30607 31977 30616 32011
rect 30564 31968 30616 31977
rect 31760 31968 31812 32020
rect 19892 31900 19944 31952
rect 21640 31943 21692 31952
rect 21640 31909 21649 31943
rect 21649 31909 21683 31943
rect 21683 31909 21692 31943
rect 21640 31900 21692 31909
rect 24584 31900 24636 31952
rect 25412 31900 25464 31952
rect 19432 31832 19484 31884
rect 19984 31832 20036 31884
rect 23020 31875 23072 31884
rect 23020 31841 23029 31875
rect 23029 31841 23063 31875
rect 23063 31841 23072 31875
rect 23020 31832 23072 31841
rect 23204 31875 23256 31884
rect 23204 31841 23213 31875
rect 23213 31841 23247 31875
rect 23247 31841 23256 31875
rect 23204 31832 23256 31841
rect 28080 31900 28132 31952
rect 28540 31900 28592 31952
rect 32128 31943 32180 31952
rect 32128 31909 32137 31943
rect 32137 31909 32171 31943
rect 32171 31909 32180 31943
rect 32128 31900 32180 31909
rect 32312 31900 32364 31952
rect 33784 31968 33836 32020
rect 33692 31943 33744 31952
rect 33692 31909 33701 31943
rect 33701 31909 33735 31943
rect 33735 31909 33744 31943
rect 33692 31900 33744 31909
rect 27528 31832 27580 31884
rect 28632 31832 28684 31884
rect 30012 31832 30064 31884
rect 30564 31832 30616 31884
rect 30748 31875 30800 31884
rect 30748 31841 30757 31875
rect 30757 31841 30791 31875
rect 30791 31841 30800 31875
rect 30748 31832 30800 31841
rect 32036 31832 32088 31884
rect 21732 31764 21784 31816
rect 23296 31807 23348 31816
rect 23296 31773 23305 31807
rect 23305 31773 23339 31807
rect 23339 31773 23348 31807
rect 23296 31764 23348 31773
rect 24032 31764 24084 31816
rect 26884 31764 26936 31816
rect 31024 31764 31076 31816
rect 32312 31807 32364 31816
rect 32312 31773 32318 31807
rect 32318 31773 32364 31807
rect 32312 31764 32364 31773
rect 32404 31764 32456 31816
rect 34888 31968 34940 32020
rect 35808 31968 35860 32020
rect 35992 31968 36044 32020
rect 41052 32011 41104 32020
rect 41052 31977 41061 32011
rect 41061 31977 41095 32011
rect 41095 31977 41104 32011
rect 41052 31968 41104 31977
rect 42892 32011 42944 32020
rect 42892 31977 42901 32011
rect 42901 31977 42935 32011
rect 42935 31977 42944 32011
rect 42892 31968 42944 31977
rect 44732 32011 44784 32020
rect 44732 31977 44741 32011
rect 44741 31977 44775 32011
rect 44775 31977 44784 32011
rect 44732 31968 44784 31977
rect 46664 32011 46716 32020
rect 46664 31977 46673 32011
rect 46673 31977 46707 32011
rect 46707 31977 46716 32011
rect 46664 31968 46716 31977
rect 36912 31943 36964 31952
rect 36912 31909 36921 31943
rect 36921 31909 36955 31943
rect 36955 31909 36964 31943
rect 36912 31900 36964 31909
rect 38660 31900 38712 31952
rect 40408 31900 40460 31952
rect 40500 31900 40552 31952
rect 41604 31943 41656 31952
rect 41604 31909 41613 31943
rect 41613 31909 41647 31943
rect 41647 31909 41656 31943
rect 41604 31900 41656 31909
rect 41696 31943 41748 31952
rect 41696 31909 41705 31943
rect 41705 31909 41739 31943
rect 41739 31909 41748 31943
rect 41696 31900 41748 31909
rect 42616 31900 42668 31952
rect 45008 31900 45060 31952
rect 45192 31900 45244 31952
rect 34704 31764 34756 31816
rect 35900 31832 35952 31884
rect 36268 31832 36320 31884
rect 38108 31832 38160 31884
rect 46388 31875 46440 31884
rect 46388 31841 46397 31875
rect 46397 31841 46431 31875
rect 46431 31841 46440 31875
rect 46388 31832 46440 31841
rect 35072 31764 35124 31816
rect 15660 31696 15712 31748
rect 14648 31628 14700 31680
rect 15292 31628 15344 31680
rect 16304 31671 16356 31680
rect 16304 31637 16313 31671
rect 16313 31637 16347 31671
rect 16347 31637 16356 31671
rect 16304 31628 16356 31637
rect 31944 31696 31996 31748
rect 32036 31696 32088 31748
rect 33600 31696 33652 31748
rect 34060 31696 34112 31748
rect 37280 31764 37332 31816
rect 39764 31807 39816 31816
rect 39764 31773 39773 31807
rect 39773 31773 39807 31807
rect 39807 31773 39816 31807
rect 39764 31764 39816 31773
rect 41880 31807 41932 31816
rect 41880 31773 41889 31807
rect 41889 31773 41923 31807
rect 41923 31773 41932 31807
rect 41880 31764 41932 31773
rect 35440 31696 35492 31748
rect 18788 31628 18840 31680
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 28356 31628 28408 31680
rect 29736 31628 29788 31680
rect 30288 31671 30340 31680
rect 30288 31637 30297 31671
rect 30297 31637 30331 31671
rect 30331 31637 30340 31671
rect 30288 31628 30340 31637
rect 32496 31628 32548 31680
rect 35532 31671 35584 31680
rect 35532 31637 35541 31671
rect 35541 31637 35575 31671
rect 35575 31637 35584 31671
rect 35532 31628 35584 31637
rect 36912 31696 36964 31748
rect 41696 31696 41748 31748
rect 43168 31764 43220 31816
rect 45836 31764 45888 31816
rect 44916 31696 44968 31748
rect 37740 31628 37792 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 13728 31424 13780 31476
rect 15384 31424 15436 31476
rect 15568 31424 15620 31476
rect 18052 31424 18104 31476
rect 19892 31424 19944 31476
rect 21732 31467 21784 31476
rect 21732 31433 21741 31467
rect 21741 31433 21775 31467
rect 21775 31433 21784 31467
rect 21732 31424 21784 31433
rect 24400 31424 24452 31476
rect 25412 31424 25464 31476
rect 27436 31424 27488 31476
rect 16856 31356 16908 31408
rect 19432 31356 19484 31408
rect 20444 31356 20496 31408
rect 24032 31399 24084 31408
rect 24032 31365 24041 31399
rect 24041 31365 24075 31399
rect 24075 31365 24084 31399
rect 24032 31356 24084 31365
rect 28264 31399 28316 31408
rect 28264 31365 28273 31399
rect 28273 31365 28307 31399
rect 28307 31365 28316 31399
rect 28264 31356 28316 31365
rect 30196 31356 30248 31408
rect 34336 31424 34388 31476
rect 34704 31424 34756 31476
rect 34796 31424 34848 31476
rect 35348 31424 35400 31476
rect 36268 31467 36320 31476
rect 36268 31433 36277 31467
rect 36277 31433 36311 31467
rect 36311 31433 36320 31467
rect 36268 31424 36320 31433
rect 38108 31424 38160 31476
rect 41052 31424 41104 31476
rect 41696 31424 41748 31476
rect 32588 31356 32640 31408
rect 43168 31424 43220 31476
rect 45192 31424 45244 31476
rect 45836 31467 45888 31476
rect 45836 31433 45845 31467
rect 45845 31433 45879 31467
rect 45879 31433 45888 31467
rect 45836 31424 45888 31433
rect 42616 31356 42668 31408
rect 15016 31288 15068 31340
rect 15200 31288 15252 31340
rect 15660 31331 15712 31340
rect 15660 31297 15669 31331
rect 15669 31297 15703 31331
rect 15703 31297 15712 31331
rect 15660 31288 15712 31297
rect 17316 31288 17368 31340
rect 18788 31263 18840 31272
rect 18788 31229 18797 31263
rect 18797 31229 18831 31263
rect 18831 31229 18840 31263
rect 21640 31288 21692 31340
rect 23204 31288 23256 31340
rect 24768 31288 24820 31340
rect 24952 31288 25004 31340
rect 31944 31331 31996 31340
rect 18788 31220 18840 31229
rect 22284 31220 22336 31272
rect 16120 31152 16172 31204
rect 16488 31152 16540 31204
rect 14740 31084 14792 31136
rect 18052 31084 18104 31136
rect 20260 31152 20312 31204
rect 19984 31084 20036 31136
rect 21272 31152 21324 31204
rect 23020 31220 23072 31272
rect 23940 31220 23992 31272
rect 31944 31297 31953 31331
rect 31953 31297 31987 31331
rect 31987 31297 31996 31331
rect 31944 31288 31996 31297
rect 37832 31288 37884 31340
rect 39764 31288 39816 31340
rect 40592 31288 40644 31340
rect 41144 31331 41196 31340
rect 41144 31297 41153 31331
rect 41153 31297 41187 31331
rect 41187 31297 41196 31331
rect 41144 31288 41196 31297
rect 29736 31263 29788 31272
rect 29736 31229 29745 31263
rect 29745 31229 29779 31263
rect 29779 31229 29788 31263
rect 29736 31220 29788 31229
rect 24584 31195 24636 31204
rect 24584 31161 24593 31195
rect 24593 31161 24627 31195
rect 24627 31161 24636 31195
rect 24584 31152 24636 31161
rect 25688 31152 25740 31204
rect 26240 31195 26292 31204
rect 21180 31084 21232 31136
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 26240 31161 26249 31195
rect 26249 31161 26283 31195
rect 26283 31161 26292 31195
rect 26240 31152 26292 31161
rect 28448 31152 28500 31204
rect 31852 31220 31904 31272
rect 31576 31195 31628 31204
rect 31576 31161 31585 31195
rect 31585 31161 31619 31195
rect 31619 31161 31628 31195
rect 31576 31152 31628 31161
rect 26700 31084 26752 31136
rect 28632 31127 28684 31136
rect 28632 31093 28641 31127
rect 28641 31093 28675 31127
rect 28675 31093 28684 31127
rect 28632 31084 28684 31093
rect 29368 31127 29420 31136
rect 29368 31093 29377 31127
rect 29377 31093 29411 31127
rect 29411 31093 29420 31127
rect 29368 31084 29420 31093
rect 30472 31127 30524 31136
rect 30472 31093 30481 31127
rect 30481 31093 30515 31127
rect 30515 31093 30524 31127
rect 30472 31084 30524 31093
rect 30840 31127 30892 31136
rect 30840 31093 30849 31127
rect 30849 31093 30883 31127
rect 30883 31093 30892 31127
rect 30840 31084 30892 31093
rect 32220 31127 32272 31136
rect 32220 31093 32229 31127
rect 32229 31093 32263 31127
rect 32263 31093 32272 31127
rect 32220 31084 32272 31093
rect 32588 31127 32640 31136
rect 32588 31093 32597 31127
rect 32597 31093 32631 31127
rect 32631 31093 32640 31127
rect 34152 31220 34204 31272
rect 34704 31220 34756 31272
rect 37188 31220 37240 31272
rect 37464 31220 37516 31272
rect 38292 31220 38344 31272
rect 38844 31263 38896 31272
rect 38844 31229 38853 31263
rect 38853 31229 38887 31263
rect 38887 31229 38896 31263
rect 38844 31220 38896 31229
rect 35900 31152 35952 31204
rect 37556 31195 37608 31204
rect 37556 31161 37565 31195
rect 37565 31161 37599 31195
rect 37599 31161 37608 31195
rect 37556 31152 37608 31161
rect 32588 31084 32640 31093
rect 34704 31084 34756 31136
rect 38660 31084 38712 31136
rect 41052 31084 41104 31136
rect 42064 31152 42116 31204
rect 43904 31288 43956 31340
rect 45284 31288 45336 31340
rect 45652 31220 45704 31272
rect 46112 31263 46164 31272
rect 46112 31229 46121 31263
rect 46121 31229 46155 31263
rect 46155 31229 46164 31263
rect 46112 31220 46164 31229
rect 43076 31195 43128 31204
rect 43076 31161 43085 31195
rect 43085 31161 43119 31195
rect 43119 31161 43128 31195
rect 43076 31152 43128 31161
rect 43720 31195 43772 31204
rect 43720 31161 43729 31195
rect 43729 31161 43763 31195
rect 43763 31161 43772 31195
rect 43720 31152 43772 31161
rect 45100 31152 45152 31204
rect 45284 31152 45336 31204
rect 46388 31152 46440 31204
rect 44824 31084 44876 31136
rect 46296 31127 46348 31136
rect 46296 31093 46305 31127
rect 46305 31093 46339 31127
rect 46339 31093 46348 31127
rect 46296 31084 46348 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 15384 30880 15436 30932
rect 16304 30880 16356 30932
rect 17684 30923 17736 30932
rect 17684 30889 17693 30923
rect 17693 30889 17727 30923
rect 17727 30889 17736 30923
rect 17684 30880 17736 30889
rect 20168 30880 20220 30932
rect 22284 30880 22336 30932
rect 14556 30812 14608 30864
rect 15292 30812 15344 30864
rect 18052 30855 18104 30864
rect 18052 30821 18061 30855
rect 18061 30821 18095 30855
rect 18095 30821 18104 30855
rect 18052 30812 18104 30821
rect 21180 30812 21232 30864
rect 12716 30744 12768 30796
rect 13268 30744 13320 30796
rect 13912 30744 13964 30796
rect 20444 30744 20496 30796
rect 20720 30744 20772 30796
rect 23296 30880 23348 30932
rect 16580 30676 16632 30728
rect 20352 30676 20404 30728
rect 18420 30608 18472 30660
rect 23112 30676 23164 30728
rect 24584 30923 24636 30932
rect 24584 30889 24593 30923
rect 24593 30889 24627 30923
rect 24627 30889 24636 30923
rect 24584 30880 24636 30889
rect 30012 30923 30064 30932
rect 30012 30889 30021 30923
rect 30021 30889 30055 30923
rect 30055 30889 30064 30923
rect 30012 30880 30064 30889
rect 31392 30880 31444 30932
rect 31668 30923 31720 30932
rect 31668 30889 31677 30923
rect 31677 30889 31711 30923
rect 31711 30889 31720 30923
rect 31668 30880 31720 30889
rect 31760 30880 31812 30932
rect 32404 30880 32456 30932
rect 34060 30923 34112 30932
rect 34060 30889 34069 30923
rect 34069 30889 34103 30923
rect 34103 30889 34112 30923
rect 34060 30880 34112 30889
rect 26700 30855 26752 30864
rect 26700 30821 26709 30855
rect 26709 30821 26743 30855
rect 26743 30821 26752 30855
rect 26700 30812 26752 30821
rect 26884 30812 26936 30864
rect 29184 30855 29236 30864
rect 29184 30821 29193 30855
rect 29193 30821 29227 30855
rect 29227 30821 29236 30855
rect 29184 30812 29236 30821
rect 32128 30855 32180 30864
rect 32128 30821 32137 30855
rect 32137 30821 32171 30855
rect 32171 30821 32180 30855
rect 32128 30812 32180 30821
rect 34704 30880 34756 30932
rect 35900 30923 35952 30932
rect 35900 30889 35909 30923
rect 35909 30889 35943 30923
rect 35943 30889 35952 30923
rect 35900 30880 35952 30889
rect 39396 30880 39448 30932
rect 40592 30880 40644 30932
rect 41144 30923 41196 30932
rect 41144 30889 41153 30923
rect 41153 30889 41187 30923
rect 41187 30889 41196 30923
rect 41144 30880 41196 30889
rect 41604 30880 41656 30932
rect 43076 30923 43128 30932
rect 43076 30889 43085 30923
rect 43085 30889 43119 30923
rect 43119 30889 43128 30923
rect 43076 30880 43128 30889
rect 41512 30855 41564 30864
rect 41512 30821 41521 30855
rect 41521 30821 41555 30855
rect 41555 30821 41564 30855
rect 41512 30812 41564 30821
rect 44640 30812 44692 30864
rect 45100 30855 45152 30864
rect 45100 30821 45109 30855
rect 45109 30821 45143 30855
rect 45143 30821 45152 30855
rect 45100 30812 45152 30821
rect 46848 30812 46900 30864
rect 24952 30787 25004 30796
rect 24952 30753 24961 30787
rect 24961 30753 24995 30787
rect 24995 30753 25004 30787
rect 24952 30744 25004 30753
rect 31116 30744 31168 30796
rect 31852 30744 31904 30796
rect 34520 30787 34572 30796
rect 34520 30753 34529 30787
rect 34529 30753 34563 30787
rect 34563 30753 34572 30787
rect 34520 30744 34572 30753
rect 36176 30744 36228 30796
rect 36912 30744 36964 30796
rect 38016 30744 38068 30796
rect 38936 30744 38988 30796
rect 39396 30744 39448 30796
rect 27436 30676 27488 30728
rect 29092 30719 29144 30728
rect 29092 30685 29101 30719
rect 29101 30685 29135 30719
rect 29135 30685 29144 30719
rect 29092 30676 29144 30685
rect 30656 30676 30708 30728
rect 31760 30676 31812 30728
rect 31944 30676 31996 30728
rect 33232 30676 33284 30728
rect 34888 30719 34940 30728
rect 34888 30685 34897 30719
rect 34897 30685 34931 30719
rect 34931 30685 34940 30719
rect 34888 30676 34940 30685
rect 38844 30719 38896 30728
rect 15476 30540 15528 30592
rect 21364 30608 21416 30660
rect 29644 30651 29696 30660
rect 29644 30617 29653 30651
rect 29653 30617 29687 30651
rect 29687 30617 29696 30651
rect 29644 30608 29696 30617
rect 29736 30608 29788 30660
rect 33140 30608 33192 30660
rect 20260 30540 20312 30592
rect 24124 30583 24176 30592
rect 24124 30549 24133 30583
rect 24133 30549 24167 30583
rect 24167 30549 24176 30583
rect 24124 30540 24176 30549
rect 26240 30583 26292 30592
rect 26240 30549 26249 30583
rect 26249 30549 26283 30583
rect 26283 30549 26292 30583
rect 26240 30540 26292 30549
rect 32496 30540 32548 30592
rect 33416 30540 33468 30592
rect 34612 30608 34664 30660
rect 37464 30608 37516 30660
rect 38844 30685 38853 30719
rect 38853 30685 38887 30719
rect 38887 30685 38896 30719
rect 39580 30744 39632 30796
rect 43260 30744 43312 30796
rect 45928 30787 45980 30796
rect 45928 30753 45937 30787
rect 45937 30753 45971 30787
rect 45971 30753 45980 30787
rect 45928 30744 45980 30753
rect 39672 30719 39724 30728
rect 38844 30676 38896 30685
rect 39672 30685 39681 30719
rect 39681 30685 39715 30719
rect 39715 30685 39724 30719
rect 39672 30676 39724 30685
rect 41880 30676 41932 30728
rect 43076 30676 43128 30728
rect 45468 30676 45520 30728
rect 35624 30583 35676 30592
rect 35624 30549 35633 30583
rect 35633 30549 35667 30583
rect 35667 30549 35676 30583
rect 35624 30540 35676 30549
rect 36268 30583 36320 30592
rect 36268 30549 36277 30583
rect 36277 30549 36311 30583
rect 36311 30549 36320 30583
rect 36268 30540 36320 30549
rect 38292 30540 38344 30592
rect 40500 30583 40552 30592
rect 40500 30549 40509 30583
rect 40509 30549 40543 30583
rect 40543 30549 40552 30583
rect 40500 30540 40552 30549
rect 47032 30540 47084 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 13268 30336 13320 30388
rect 15108 30336 15160 30388
rect 15292 30379 15344 30388
rect 15292 30345 15301 30379
rect 15301 30345 15335 30379
rect 15335 30345 15344 30379
rect 15292 30336 15344 30345
rect 16580 30379 16632 30388
rect 16580 30345 16589 30379
rect 16589 30345 16623 30379
rect 16623 30345 16632 30379
rect 16580 30336 16632 30345
rect 18052 30336 18104 30388
rect 18420 30336 18472 30388
rect 20168 30379 20220 30388
rect 20168 30345 20177 30379
rect 20177 30345 20211 30379
rect 20211 30345 20220 30379
rect 20168 30336 20220 30345
rect 21180 30336 21232 30388
rect 22376 30379 22428 30388
rect 22376 30345 22385 30379
rect 22385 30345 22419 30379
rect 22419 30345 22428 30379
rect 22376 30336 22428 30345
rect 23112 30336 23164 30388
rect 23756 30336 23808 30388
rect 24400 30336 24452 30388
rect 25688 30379 25740 30388
rect 25688 30345 25697 30379
rect 25697 30345 25731 30379
rect 25731 30345 25740 30379
rect 25688 30336 25740 30345
rect 27436 30379 27488 30388
rect 27436 30345 27445 30379
rect 27445 30345 27479 30379
rect 27479 30345 27488 30379
rect 27436 30336 27488 30345
rect 31024 30336 31076 30388
rect 32588 30336 32640 30388
rect 20260 30268 20312 30320
rect 21272 30311 21324 30320
rect 21272 30277 21281 30311
rect 21281 30277 21315 30311
rect 21315 30277 21324 30311
rect 21272 30268 21324 30277
rect 22836 30268 22888 30320
rect 28632 30268 28684 30320
rect 31944 30268 31996 30320
rect 33784 30336 33836 30388
rect 34796 30336 34848 30388
rect 35532 30336 35584 30388
rect 35900 30336 35952 30388
rect 37464 30379 37516 30388
rect 37464 30345 37473 30379
rect 37473 30345 37507 30379
rect 37507 30345 37516 30379
rect 37464 30336 37516 30345
rect 37740 30379 37792 30388
rect 37740 30345 37749 30379
rect 37749 30345 37783 30379
rect 37783 30345 37792 30379
rect 37740 30336 37792 30345
rect 38016 30379 38068 30388
rect 38016 30345 38025 30379
rect 38025 30345 38059 30379
rect 38059 30345 38068 30379
rect 38016 30336 38068 30345
rect 38476 30379 38528 30388
rect 38476 30345 38485 30379
rect 38485 30345 38519 30379
rect 38519 30345 38528 30379
rect 38476 30336 38528 30345
rect 41880 30336 41932 30388
rect 43260 30336 43312 30388
rect 44364 30336 44416 30388
rect 45100 30336 45152 30388
rect 45468 30379 45520 30388
rect 34612 30268 34664 30320
rect 29368 30200 29420 30252
rect 31852 30243 31904 30252
rect 31852 30209 31861 30243
rect 31861 30209 31895 30243
rect 31895 30209 31904 30243
rect 31852 30200 31904 30209
rect 34060 30200 34112 30252
rect 34520 30200 34572 30252
rect 36176 30268 36228 30320
rect 45468 30345 45477 30379
rect 45477 30345 45511 30379
rect 45511 30345 45520 30379
rect 45468 30336 45520 30345
rect 47584 30379 47636 30388
rect 47584 30345 47593 30379
rect 47593 30345 47627 30379
rect 47627 30345 47636 30379
rect 47584 30336 47636 30345
rect 45928 30268 45980 30320
rect 12716 30039 12768 30048
rect 12716 30005 12725 30039
rect 12725 30005 12759 30039
rect 12759 30005 12768 30039
rect 12716 29996 12768 30005
rect 13084 30039 13136 30048
rect 13084 30005 13093 30039
rect 13093 30005 13127 30039
rect 13127 30005 13136 30039
rect 13084 29996 13136 30005
rect 14096 30039 14148 30048
rect 14096 30005 14105 30039
rect 14105 30005 14139 30039
rect 14139 30005 14148 30039
rect 14096 29996 14148 30005
rect 20168 30132 20220 30184
rect 15476 30064 15528 30116
rect 15752 30107 15804 30116
rect 15752 30073 15761 30107
rect 15761 30073 15795 30107
rect 15795 30073 15804 30107
rect 15752 30064 15804 30073
rect 16488 30064 16540 30116
rect 16580 29996 16632 30048
rect 16948 30039 17000 30048
rect 16948 30005 16957 30039
rect 16957 30005 16991 30039
rect 16991 30005 17000 30039
rect 16948 29996 17000 30005
rect 17776 30039 17828 30048
rect 17776 30005 17785 30039
rect 17785 30005 17819 30039
rect 17819 30005 17828 30039
rect 18236 30107 18288 30116
rect 18236 30073 18245 30107
rect 18245 30073 18279 30107
rect 18279 30073 18288 30107
rect 18788 30107 18840 30116
rect 18236 30064 18288 30073
rect 18788 30073 18797 30107
rect 18797 30073 18831 30107
rect 18831 30073 18840 30107
rect 18788 30064 18840 30073
rect 22744 30175 22796 30184
rect 22744 30141 22753 30175
rect 22753 30141 22787 30175
rect 22787 30141 22796 30175
rect 22744 30132 22796 30141
rect 23664 30175 23716 30184
rect 23664 30141 23673 30175
rect 23673 30141 23707 30175
rect 23707 30141 23716 30175
rect 23664 30132 23716 30141
rect 26332 30132 26384 30184
rect 20720 30064 20772 30116
rect 21088 30064 21140 30116
rect 23756 30064 23808 30116
rect 26148 30107 26200 30116
rect 26148 30073 26157 30107
rect 26157 30073 26191 30107
rect 26191 30073 26200 30107
rect 26148 30064 26200 30073
rect 29184 30132 29236 30184
rect 31116 30132 31168 30184
rect 32496 30132 32548 30184
rect 33416 30175 33468 30184
rect 33416 30141 33422 30175
rect 33422 30141 33468 30175
rect 36360 30243 36412 30252
rect 36360 30209 36369 30243
rect 36369 30209 36403 30243
rect 36403 30209 36412 30243
rect 36360 30200 36412 30209
rect 39304 30200 39356 30252
rect 41512 30200 41564 30252
rect 42800 30243 42852 30252
rect 42800 30209 42809 30243
rect 42809 30209 42843 30243
rect 42843 30209 42852 30243
rect 43076 30243 43128 30252
rect 42800 30200 42852 30209
rect 43076 30209 43085 30243
rect 43085 30209 43119 30243
rect 43119 30209 43128 30243
rect 43076 30200 43128 30209
rect 45008 30243 45060 30252
rect 45008 30209 45017 30243
rect 45017 30209 45051 30243
rect 45051 30209 45060 30243
rect 45008 30200 45060 30209
rect 33416 30132 33468 30141
rect 36268 30132 36320 30184
rect 37556 30175 37608 30184
rect 37556 30141 37565 30175
rect 37565 30141 37599 30175
rect 37599 30141 37608 30175
rect 37556 30132 37608 30141
rect 38476 30132 38528 30184
rect 39580 30132 39632 30184
rect 39764 30132 39816 30184
rect 40500 30175 40552 30184
rect 40500 30141 40509 30175
rect 40509 30141 40543 30175
rect 40543 30141 40552 30175
rect 40500 30132 40552 30141
rect 46940 30200 46992 30252
rect 47032 30132 47084 30184
rect 17776 29996 17828 30005
rect 19984 29996 20036 30048
rect 20444 30039 20496 30048
rect 20444 30005 20453 30039
rect 20453 30005 20487 30039
rect 20487 30005 20496 30039
rect 20444 29996 20496 30005
rect 24952 30039 25004 30048
rect 24952 30005 24961 30039
rect 24961 30005 24995 30039
rect 24995 30005 25004 30039
rect 24952 29996 25004 30005
rect 27160 30039 27212 30048
rect 27160 30005 27169 30039
rect 27169 30005 27203 30039
rect 27203 30005 27212 30039
rect 27160 29996 27212 30005
rect 29092 30064 29144 30116
rect 28724 29996 28776 30048
rect 31668 30064 31720 30116
rect 32956 30064 33008 30116
rect 34704 30064 34756 30116
rect 35624 30064 35676 30116
rect 37280 30064 37332 30116
rect 40684 30064 40736 30116
rect 44548 30107 44600 30116
rect 31392 29996 31444 30048
rect 32588 30039 32640 30048
rect 32588 30005 32597 30039
rect 32597 30005 32631 30039
rect 32631 30005 32640 30039
rect 32588 29996 32640 30005
rect 35808 29996 35860 30048
rect 37096 30039 37148 30048
rect 37096 30005 37105 30039
rect 37105 30005 37139 30039
rect 37139 30005 37148 30039
rect 37096 29996 37148 30005
rect 39488 29996 39540 30048
rect 40224 30039 40276 30048
rect 40224 30005 40233 30039
rect 40233 30005 40267 30039
rect 40267 30005 40276 30039
rect 41420 30039 41472 30048
rect 40224 29996 40276 30005
rect 41420 30005 41429 30039
rect 41429 30005 41463 30039
rect 41463 30005 41472 30039
rect 41420 29996 41472 30005
rect 42432 29996 42484 30048
rect 44548 30073 44557 30107
rect 44557 30073 44591 30107
rect 44591 30073 44600 30107
rect 44548 30064 44600 30073
rect 44640 30107 44692 30116
rect 44640 30073 44649 30107
rect 44649 30073 44683 30107
rect 44683 30073 44692 30107
rect 44640 30064 44692 30073
rect 46388 29996 46440 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 14372 29792 14424 29844
rect 15476 29792 15528 29844
rect 15752 29792 15804 29844
rect 16948 29792 17000 29844
rect 17776 29792 17828 29844
rect 18052 29835 18104 29844
rect 18052 29801 18061 29835
rect 18061 29801 18095 29835
rect 18095 29801 18104 29835
rect 18052 29792 18104 29801
rect 20352 29835 20404 29844
rect 20352 29801 20361 29835
rect 20361 29801 20395 29835
rect 20395 29801 20404 29835
rect 20352 29792 20404 29801
rect 23756 29835 23808 29844
rect 23756 29801 23765 29835
rect 23765 29801 23799 29835
rect 23799 29801 23808 29835
rect 23756 29792 23808 29801
rect 28724 29792 28776 29844
rect 29368 29792 29420 29844
rect 30472 29792 30524 29844
rect 31484 29792 31536 29844
rect 31668 29792 31720 29844
rect 32128 29792 32180 29844
rect 33232 29792 33284 29844
rect 34520 29835 34572 29844
rect 34520 29801 34529 29835
rect 34529 29801 34563 29835
rect 34563 29801 34572 29835
rect 34520 29792 34572 29801
rect 35624 29792 35676 29844
rect 35900 29792 35952 29844
rect 36176 29835 36228 29844
rect 36176 29801 36185 29835
rect 36185 29801 36219 29835
rect 36219 29801 36228 29835
rect 36176 29792 36228 29801
rect 36268 29792 36320 29844
rect 37004 29792 37056 29844
rect 38660 29792 38712 29844
rect 39304 29835 39356 29844
rect 39304 29801 39313 29835
rect 39313 29801 39347 29835
rect 39347 29801 39356 29835
rect 39304 29792 39356 29801
rect 39672 29792 39724 29844
rect 40500 29792 40552 29844
rect 42432 29835 42484 29844
rect 42432 29801 42441 29835
rect 42441 29801 42475 29835
rect 42475 29801 42484 29835
rect 42432 29792 42484 29801
rect 14556 29724 14608 29776
rect 15292 29724 15344 29776
rect 18420 29767 18472 29776
rect 18420 29733 18429 29767
rect 18429 29733 18463 29767
rect 18463 29733 18472 29767
rect 18420 29724 18472 29733
rect 21088 29767 21140 29776
rect 21088 29733 21097 29767
rect 21097 29733 21131 29767
rect 21131 29733 21140 29767
rect 21088 29724 21140 29733
rect 23664 29724 23716 29776
rect 24124 29724 24176 29776
rect 27160 29724 27212 29776
rect 29184 29724 29236 29776
rect 31852 29724 31904 29776
rect 34336 29724 34388 29776
rect 13912 29656 13964 29708
rect 19892 29656 19944 29708
rect 20812 29656 20864 29708
rect 22928 29699 22980 29708
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 23204 29699 23256 29708
rect 23204 29665 23213 29699
rect 23213 29665 23247 29699
rect 23247 29665 23256 29699
rect 23204 29656 23256 29665
rect 31024 29699 31076 29708
rect 31024 29665 31033 29699
rect 31033 29665 31067 29699
rect 31067 29665 31076 29699
rect 31024 29656 31076 29665
rect 13728 29588 13780 29640
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 15292 29631 15344 29640
rect 15292 29597 15301 29631
rect 15301 29597 15335 29631
rect 15335 29597 15344 29631
rect 15292 29588 15344 29597
rect 18788 29588 18840 29640
rect 19984 29588 20036 29640
rect 16488 29520 16540 29572
rect 18972 29520 19024 29572
rect 24768 29588 24820 29640
rect 26884 29588 26936 29640
rect 28264 29588 28316 29640
rect 33692 29656 33744 29708
rect 34704 29656 34756 29708
rect 33324 29588 33376 29640
rect 35348 29588 35400 29640
rect 24676 29520 24728 29572
rect 29644 29520 29696 29572
rect 33048 29520 33100 29572
rect 33968 29520 34020 29572
rect 37556 29724 37608 29776
rect 42524 29724 42576 29776
rect 44640 29835 44692 29844
rect 44640 29801 44649 29835
rect 44649 29801 44683 29835
rect 44683 29801 44692 29835
rect 44640 29792 44692 29801
rect 36636 29699 36688 29708
rect 36636 29665 36645 29699
rect 36645 29665 36679 29699
rect 36679 29665 36688 29699
rect 36636 29656 36688 29665
rect 40132 29699 40184 29708
rect 40132 29665 40141 29699
rect 40141 29665 40175 29699
rect 40175 29665 40184 29699
rect 40132 29656 40184 29665
rect 40684 29656 40736 29708
rect 41512 29699 41564 29708
rect 41512 29665 41521 29699
rect 41521 29665 41555 29699
rect 41555 29665 41564 29699
rect 41512 29656 41564 29665
rect 42800 29699 42852 29708
rect 42800 29665 42809 29699
rect 42809 29665 42843 29699
rect 42843 29665 42852 29699
rect 43352 29699 43404 29708
rect 42800 29656 42852 29665
rect 43352 29665 43361 29699
rect 43361 29665 43395 29699
rect 43395 29665 43404 29699
rect 43352 29656 43404 29665
rect 46940 29699 46992 29708
rect 46940 29665 46949 29699
rect 46949 29665 46983 29699
rect 46983 29665 46992 29699
rect 46940 29656 46992 29665
rect 47216 29656 47268 29708
rect 38384 29631 38436 29640
rect 38384 29597 38393 29631
rect 38393 29597 38427 29631
rect 38427 29597 38436 29631
rect 38384 29588 38436 29597
rect 45376 29588 45428 29640
rect 45560 29631 45612 29640
rect 45560 29597 45569 29631
rect 45569 29597 45603 29631
rect 45603 29597 45612 29631
rect 45560 29588 45612 29597
rect 20168 29452 20220 29504
rect 26332 29495 26384 29504
rect 26332 29461 26341 29495
rect 26341 29461 26375 29495
rect 26375 29461 26384 29495
rect 26332 29452 26384 29461
rect 29460 29452 29512 29504
rect 33232 29452 33284 29504
rect 34336 29452 34388 29504
rect 34520 29452 34572 29504
rect 37740 29520 37792 29572
rect 40316 29563 40368 29572
rect 40316 29529 40325 29563
rect 40325 29529 40359 29563
rect 40359 29529 40368 29563
rect 40316 29520 40368 29529
rect 36360 29452 36412 29504
rect 37464 29452 37516 29504
rect 38016 29495 38068 29504
rect 38016 29461 38025 29495
rect 38025 29461 38059 29495
rect 38059 29461 38068 29495
rect 38016 29452 38068 29461
rect 39580 29495 39632 29504
rect 39580 29461 39589 29495
rect 39589 29461 39623 29495
rect 39623 29461 39632 29495
rect 39580 29452 39632 29461
rect 46848 29495 46900 29504
rect 46848 29461 46857 29495
rect 46857 29461 46891 29495
rect 46891 29461 46900 29495
rect 46848 29452 46900 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 13360 29248 13412 29300
rect 15200 29248 15252 29300
rect 16672 29180 16724 29232
rect 17224 29180 17276 29232
rect 14372 29112 14424 29164
rect 13360 29087 13412 29096
rect 13360 29053 13369 29087
rect 13369 29053 13403 29087
rect 13403 29053 13412 29087
rect 13360 29044 13412 29053
rect 13820 29087 13872 29096
rect 13820 29053 13829 29087
rect 13829 29053 13863 29087
rect 13863 29053 13872 29087
rect 13820 29044 13872 29053
rect 15292 29044 15344 29096
rect 14556 28908 14608 28960
rect 15200 28951 15252 28960
rect 15200 28917 15209 28951
rect 15209 28917 15243 28951
rect 15243 28917 15252 28951
rect 15200 28908 15252 28917
rect 15936 28908 15988 28960
rect 18420 29248 18472 29300
rect 19984 29248 20036 29300
rect 21088 29248 21140 29300
rect 23204 29248 23256 29300
rect 24124 29248 24176 29300
rect 24676 29291 24728 29300
rect 24676 29257 24685 29291
rect 24685 29257 24719 29291
rect 24719 29257 24728 29291
rect 24676 29248 24728 29257
rect 24768 29248 24820 29300
rect 27160 29248 27212 29300
rect 28356 29291 28408 29300
rect 28356 29257 28365 29291
rect 28365 29257 28399 29291
rect 28399 29257 28408 29291
rect 28356 29248 28408 29257
rect 18788 29180 18840 29232
rect 21364 29223 21416 29232
rect 21364 29189 21373 29223
rect 21373 29189 21407 29223
rect 21407 29189 21416 29223
rect 21364 29180 21416 29189
rect 20168 29112 20220 29164
rect 21272 29112 21324 29164
rect 26332 29155 26384 29164
rect 26332 29121 26341 29155
rect 26341 29121 26375 29155
rect 26375 29121 26384 29155
rect 26332 29112 26384 29121
rect 26884 29112 26936 29164
rect 18052 29087 18104 29096
rect 18052 29053 18061 29087
rect 18061 29053 18095 29087
rect 18095 29053 18104 29087
rect 18052 29044 18104 29053
rect 19892 29019 19944 29028
rect 19892 28985 19901 29019
rect 19901 28985 19935 29019
rect 19935 28985 19944 29019
rect 19892 28976 19944 28985
rect 21088 28976 21140 29028
rect 21824 28976 21876 29028
rect 22928 28976 22980 29028
rect 24676 29044 24728 29096
rect 30012 29248 30064 29300
rect 32588 29248 32640 29300
rect 35900 29248 35952 29300
rect 37004 29248 37056 29300
rect 33508 29223 33560 29232
rect 33508 29189 33517 29223
rect 33517 29189 33551 29223
rect 33551 29189 33560 29223
rect 33508 29180 33560 29189
rect 37280 29180 37332 29232
rect 29644 29155 29696 29164
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 33784 29112 33836 29164
rect 34520 29112 34572 29164
rect 35256 29112 35308 29164
rect 36268 29112 36320 29164
rect 36360 29155 36412 29164
rect 36360 29121 36369 29155
rect 36369 29121 36403 29155
rect 36403 29121 36412 29155
rect 36360 29112 36412 29121
rect 36636 29112 36688 29164
rect 37004 29155 37056 29164
rect 37004 29121 37013 29155
rect 37013 29121 37047 29155
rect 37047 29121 37056 29155
rect 37004 29112 37056 29121
rect 31668 29087 31720 29096
rect 17592 28908 17644 28960
rect 22652 28908 22704 28960
rect 23480 28951 23532 28960
rect 23480 28917 23489 28951
rect 23489 28917 23523 28951
rect 23523 28917 23532 28951
rect 23480 28908 23532 28917
rect 24124 28908 24176 28960
rect 25872 28976 25924 29028
rect 28356 28976 28408 29028
rect 28448 28976 28500 29028
rect 29368 29019 29420 29028
rect 29368 28985 29377 29019
rect 29377 28985 29411 29019
rect 29411 28985 29420 29019
rect 29368 28976 29420 28985
rect 29460 29019 29512 29028
rect 29460 28985 29469 29019
rect 29469 28985 29503 29019
rect 29503 28985 29512 29019
rect 29460 28976 29512 28985
rect 31024 28976 31076 29028
rect 31668 29053 31677 29087
rect 31677 29053 31711 29087
rect 31711 29053 31720 29087
rect 31668 29044 31720 29053
rect 33692 29044 33744 29096
rect 31576 28976 31628 29028
rect 32956 28976 33008 29028
rect 43352 29248 43404 29300
rect 44640 29248 44692 29300
rect 47032 29291 47084 29300
rect 47032 29257 47041 29291
rect 47041 29257 47075 29291
rect 47075 29257 47084 29291
rect 47032 29248 47084 29257
rect 39028 29180 39080 29232
rect 40132 29180 40184 29232
rect 42524 29180 42576 29232
rect 46940 29180 46992 29232
rect 38016 29112 38068 29164
rect 39580 29112 39632 29164
rect 40500 29155 40552 29164
rect 40500 29121 40509 29155
rect 40509 29121 40543 29155
rect 40543 29121 40552 29155
rect 40500 29112 40552 29121
rect 42156 29112 42208 29164
rect 42340 29155 42392 29164
rect 42340 29121 42349 29155
rect 42349 29121 42383 29155
rect 42383 29121 42392 29155
rect 42340 29112 42392 29121
rect 43076 29112 43128 29164
rect 44824 29112 44876 29164
rect 44916 29155 44968 29164
rect 44916 29121 44925 29155
rect 44925 29121 44959 29155
rect 44959 29121 44968 29155
rect 44916 29112 44968 29121
rect 38384 29087 38436 29096
rect 38384 29053 38393 29087
rect 38393 29053 38427 29087
rect 38427 29053 38436 29087
rect 38384 29044 38436 29053
rect 47216 29087 47268 29096
rect 34336 28976 34388 29028
rect 34520 28976 34572 29028
rect 34704 28976 34756 29028
rect 36084 28976 36136 29028
rect 26424 28908 26476 28960
rect 28264 28908 28316 28960
rect 28724 28951 28776 28960
rect 28724 28917 28733 28951
rect 28733 28917 28767 28951
rect 28767 28917 28776 28951
rect 28724 28908 28776 28917
rect 31484 28951 31536 28960
rect 31484 28917 31493 28951
rect 31493 28917 31527 28951
rect 31527 28917 31536 28951
rect 31484 28908 31536 28917
rect 31760 28908 31812 28960
rect 34244 28951 34296 28960
rect 34244 28917 34253 28951
rect 34253 28917 34287 28951
rect 34287 28917 34296 28951
rect 34244 28908 34296 28917
rect 38660 28908 38712 28960
rect 38936 28908 38988 28960
rect 39396 28951 39448 28960
rect 39396 28917 39405 28951
rect 39405 28917 39439 28951
rect 39439 28917 39448 28951
rect 39396 28908 39448 28917
rect 40224 28951 40276 28960
rect 40224 28917 40233 28951
rect 40233 28917 40267 28951
rect 40267 28917 40276 28951
rect 40224 28908 40276 28917
rect 47216 29053 47225 29087
rect 47225 29053 47259 29087
rect 47259 29053 47268 29087
rect 47216 29044 47268 29053
rect 44640 29019 44692 29028
rect 44640 28985 44649 29019
rect 44649 28985 44683 29019
rect 44683 28985 44692 29019
rect 44640 28976 44692 28985
rect 42524 28908 42576 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 13084 28704 13136 28756
rect 13728 28704 13780 28756
rect 15292 28704 15344 28756
rect 13820 28636 13872 28688
rect 16396 28704 16448 28756
rect 18420 28747 18472 28756
rect 15936 28679 15988 28688
rect 15936 28645 15945 28679
rect 15945 28645 15979 28679
rect 15979 28645 15988 28679
rect 15936 28636 15988 28645
rect 18420 28713 18429 28747
rect 18429 28713 18463 28747
rect 18463 28713 18472 28747
rect 18420 28704 18472 28713
rect 19156 28747 19208 28756
rect 19156 28713 19165 28747
rect 19165 28713 19199 28747
rect 19199 28713 19208 28747
rect 19156 28704 19208 28713
rect 21272 28704 21324 28756
rect 18052 28679 18104 28688
rect 18052 28645 18061 28679
rect 18061 28645 18095 28679
rect 18095 28645 18104 28679
rect 18052 28636 18104 28645
rect 17224 28568 17276 28620
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 19248 28568 19300 28620
rect 19340 28568 19392 28620
rect 20904 28611 20956 28620
rect 14372 28500 14424 28552
rect 15476 28500 15528 28552
rect 15844 28543 15896 28552
rect 15844 28509 15853 28543
rect 15853 28509 15887 28543
rect 15887 28509 15896 28543
rect 15844 28500 15896 28509
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 17224 28364 17276 28416
rect 20904 28577 20913 28611
rect 20913 28577 20947 28611
rect 20947 28577 20956 28611
rect 20904 28568 20956 28577
rect 22836 28704 22888 28756
rect 24216 28704 24268 28756
rect 25872 28747 25924 28756
rect 25872 28713 25881 28747
rect 25881 28713 25915 28747
rect 25915 28713 25924 28747
rect 25872 28704 25924 28713
rect 26240 28704 26292 28756
rect 28264 28747 28316 28756
rect 28264 28713 28273 28747
rect 28273 28713 28307 28747
rect 28307 28713 28316 28747
rect 28264 28704 28316 28713
rect 29460 28704 29512 28756
rect 30012 28704 30064 28756
rect 32220 28747 32272 28756
rect 32220 28713 32229 28747
rect 32229 28713 32263 28747
rect 32263 28713 32272 28747
rect 32220 28704 32272 28713
rect 33508 28704 33560 28756
rect 34520 28704 34572 28756
rect 35348 28747 35400 28756
rect 35348 28713 35357 28747
rect 35357 28713 35391 28747
rect 35391 28713 35400 28747
rect 35348 28704 35400 28713
rect 37648 28704 37700 28756
rect 38292 28704 38344 28756
rect 38384 28704 38436 28756
rect 38936 28704 38988 28756
rect 40224 28704 40276 28756
rect 41512 28747 41564 28756
rect 41512 28713 41521 28747
rect 41521 28713 41555 28747
rect 41555 28713 41564 28747
rect 41512 28704 41564 28713
rect 42340 28704 42392 28756
rect 44548 28747 44600 28756
rect 44548 28713 44557 28747
rect 44557 28713 44591 28747
rect 44591 28713 44600 28747
rect 44548 28704 44600 28713
rect 44824 28704 44876 28756
rect 26148 28636 26200 28688
rect 23480 28568 23532 28620
rect 22744 28543 22796 28552
rect 22744 28509 22753 28543
rect 22753 28509 22787 28543
rect 22787 28509 22796 28543
rect 22744 28500 22796 28509
rect 26700 28568 26752 28620
rect 26976 28568 27028 28620
rect 28172 28611 28224 28620
rect 28172 28577 28181 28611
rect 28181 28577 28215 28611
rect 28215 28577 28224 28611
rect 28172 28568 28224 28577
rect 28356 28568 28408 28620
rect 29368 28568 29420 28620
rect 30104 28636 30156 28688
rect 32036 28636 32088 28688
rect 33692 28679 33744 28688
rect 33692 28645 33701 28679
rect 33701 28645 33735 28679
rect 33735 28645 33744 28679
rect 39764 28679 39816 28688
rect 33692 28636 33744 28645
rect 31024 28611 31076 28620
rect 31024 28577 31033 28611
rect 31033 28577 31067 28611
rect 31067 28577 31076 28611
rect 31024 28568 31076 28577
rect 31392 28568 31444 28620
rect 32496 28568 32548 28620
rect 32680 28611 32732 28620
rect 32680 28577 32689 28611
rect 32689 28577 32723 28611
rect 32723 28577 32732 28611
rect 32680 28568 32732 28577
rect 34336 28611 34388 28620
rect 34336 28577 34345 28611
rect 34345 28577 34379 28611
rect 34379 28577 34388 28611
rect 34336 28568 34388 28577
rect 35256 28568 35308 28620
rect 36084 28611 36136 28620
rect 36084 28577 36093 28611
rect 36093 28577 36127 28611
rect 36127 28577 36136 28611
rect 36084 28568 36136 28577
rect 37096 28568 37148 28620
rect 37740 28611 37792 28620
rect 37740 28577 37749 28611
rect 37749 28577 37783 28611
rect 37783 28577 37792 28611
rect 37740 28568 37792 28577
rect 39764 28645 39773 28679
rect 39773 28645 39807 28679
rect 39807 28645 39816 28679
rect 39764 28636 39816 28645
rect 41420 28636 41472 28688
rect 42064 28636 42116 28688
rect 39304 28568 39356 28620
rect 39580 28611 39632 28620
rect 39580 28577 39589 28611
rect 39589 28577 39623 28611
rect 39623 28577 39632 28611
rect 39580 28568 39632 28577
rect 40592 28611 40644 28620
rect 40592 28577 40601 28611
rect 40601 28577 40635 28611
rect 40635 28577 40644 28611
rect 40592 28568 40644 28577
rect 43076 28568 43128 28620
rect 45744 28568 45796 28620
rect 47124 28568 47176 28620
rect 24492 28543 24544 28552
rect 24492 28509 24501 28543
rect 24501 28509 24535 28543
rect 24535 28509 24544 28543
rect 24492 28500 24544 28509
rect 30472 28500 30524 28552
rect 31668 28500 31720 28552
rect 34060 28500 34112 28552
rect 41788 28500 41840 28552
rect 23204 28432 23256 28484
rect 24216 28432 24268 28484
rect 24308 28432 24360 28484
rect 34612 28475 34664 28484
rect 34612 28441 34621 28475
rect 34621 28441 34655 28475
rect 34655 28441 34664 28475
rect 34612 28432 34664 28441
rect 21088 28407 21140 28416
rect 21088 28373 21097 28407
rect 21097 28373 21131 28407
rect 21131 28373 21140 28407
rect 21088 28364 21140 28373
rect 21456 28364 21508 28416
rect 25412 28407 25464 28416
rect 25412 28373 25421 28407
rect 25421 28373 25455 28407
rect 25455 28373 25464 28407
rect 25412 28364 25464 28373
rect 34704 28364 34756 28416
rect 38476 28407 38528 28416
rect 38476 28373 38485 28407
rect 38485 28373 38519 28407
rect 38519 28373 38528 28407
rect 38476 28364 38528 28373
rect 40960 28364 41012 28416
rect 41144 28407 41196 28416
rect 41144 28373 41153 28407
rect 41153 28373 41187 28407
rect 41187 28373 41196 28407
rect 41144 28364 41196 28373
rect 43168 28364 43220 28416
rect 45376 28407 45428 28416
rect 45376 28373 45385 28407
rect 45385 28373 45419 28407
rect 45419 28373 45428 28407
rect 45376 28364 45428 28373
rect 46204 28364 46256 28416
rect 46756 28407 46808 28416
rect 46756 28373 46765 28407
rect 46765 28373 46799 28407
rect 46799 28373 46808 28407
rect 46756 28364 46808 28373
rect 47216 28364 47268 28416
rect 48228 28364 48280 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 14372 28160 14424 28212
rect 15476 28203 15528 28212
rect 15476 28169 15485 28203
rect 15485 28169 15519 28203
rect 15519 28169 15528 28203
rect 15476 28160 15528 28169
rect 15936 28160 15988 28212
rect 17776 28203 17828 28212
rect 17776 28169 17785 28203
rect 17785 28169 17819 28203
rect 17819 28169 17828 28203
rect 17776 28160 17828 28169
rect 19340 28203 19392 28212
rect 13636 27999 13688 28008
rect 13636 27965 13645 27999
rect 13645 27965 13679 27999
rect 13679 27965 13688 27999
rect 13636 27956 13688 27965
rect 16672 27999 16724 28008
rect 13728 27888 13780 27940
rect 16672 27965 16681 27999
rect 16681 27965 16715 27999
rect 16715 27965 16724 27999
rect 16672 27956 16724 27965
rect 17500 27956 17552 28008
rect 17132 27931 17184 27940
rect 17132 27897 17141 27931
rect 17141 27897 17175 27931
rect 17175 27897 17184 27931
rect 17132 27888 17184 27897
rect 19340 28169 19349 28203
rect 19349 28169 19383 28203
rect 19383 28169 19392 28203
rect 19340 28160 19392 28169
rect 20904 28203 20956 28212
rect 20904 28169 20913 28203
rect 20913 28169 20947 28203
rect 20947 28169 20956 28203
rect 20904 28160 20956 28169
rect 22836 28203 22888 28212
rect 22836 28169 22845 28203
rect 22845 28169 22879 28203
rect 22879 28169 22888 28203
rect 22836 28160 22888 28169
rect 28172 28160 28224 28212
rect 30104 28203 30156 28212
rect 30104 28169 30113 28203
rect 30113 28169 30147 28203
rect 30147 28169 30156 28203
rect 30104 28160 30156 28169
rect 31024 28203 31076 28212
rect 31024 28169 31033 28203
rect 31033 28169 31067 28203
rect 31067 28169 31076 28203
rect 31024 28160 31076 28169
rect 31852 28160 31904 28212
rect 32404 28160 32456 28212
rect 32680 28160 32732 28212
rect 34060 28203 34112 28212
rect 34060 28169 34069 28203
rect 34069 28169 34103 28203
rect 34103 28169 34112 28203
rect 34060 28160 34112 28169
rect 34612 28160 34664 28212
rect 35256 28160 35308 28212
rect 36360 28160 36412 28212
rect 37188 28160 37240 28212
rect 39304 28160 39356 28212
rect 39580 28160 39632 28212
rect 40224 28160 40276 28212
rect 40592 28160 40644 28212
rect 42064 28203 42116 28212
rect 42064 28169 42073 28203
rect 42073 28169 42107 28203
rect 42107 28169 42116 28203
rect 42064 28160 42116 28169
rect 43076 28160 43128 28212
rect 45376 28160 45428 28212
rect 19248 28092 19300 28144
rect 28264 28092 28316 28144
rect 33324 28092 33376 28144
rect 39488 28092 39540 28144
rect 41880 28092 41932 28144
rect 24492 28067 24544 28076
rect 24492 28033 24501 28067
rect 24501 28033 24535 28067
rect 24535 28033 24544 28067
rect 24492 28024 24544 28033
rect 26056 28024 26108 28076
rect 26332 28024 26384 28076
rect 21088 27956 21140 28008
rect 21824 27999 21876 28008
rect 21824 27965 21833 27999
rect 21833 27965 21867 27999
rect 21867 27965 21876 27999
rect 21824 27956 21876 27965
rect 21456 27888 21508 27940
rect 22652 27956 22704 28008
rect 23480 27999 23532 28008
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 24124 27956 24176 28008
rect 24308 27999 24360 28008
rect 24308 27965 24317 27999
rect 24317 27965 24351 27999
rect 24351 27965 24360 27999
rect 24308 27956 24360 27965
rect 25688 27999 25740 28008
rect 25688 27965 25697 27999
rect 25697 27965 25731 27999
rect 25731 27965 25740 27999
rect 25688 27956 25740 27965
rect 28356 28024 28408 28076
rect 31484 28067 31536 28076
rect 31484 28033 31493 28067
rect 31493 28033 31527 28067
rect 31527 28033 31536 28067
rect 31484 28024 31536 28033
rect 29184 27956 29236 28008
rect 30472 27999 30524 28008
rect 30472 27965 30481 27999
rect 30481 27965 30515 27999
rect 30515 27965 30524 27999
rect 30472 27956 30524 27965
rect 30840 27956 30892 28008
rect 33048 27956 33100 28008
rect 26148 27888 26200 27940
rect 30932 27888 30984 27940
rect 31852 27888 31904 27940
rect 32036 27888 32088 27940
rect 14464 27863 14516 27872
rect 14464 27829 14473 27863
rect 14473 27829 14507 27863
rect 14507 27829 14516 27863
rect 14464 27820 14516 27829
rect 17224 27820 17276 27872
rect 18236 27863 18288 27872
rect 18236 27829 18245 27863
rect 18245 27829 18279 27863
rect 18279 27829 18288 27863
rect 18236 27820 18288 27829
rect 19984 27863 20036 27872
rect 19984 27829 19993 27863
rect 19993 27829 20027 27863
rect 20027 27829 20036 27863
rect 19984 27820 20036 27829
rect 21916 27863 21968 27872
rect 21916 27829 21925 27863
rect 21925 27829 21959 27863
rect 21959 27829 21968 27863
rect 21916 27820 21968 27829
rect 26608 27863 26660 27872
rect 26608 27829 26617 27863
rect 26617 27829 26651 27863
rect 26651 27829 26660 27863
rect 26608 27820 26660 27829
rect 26700 27820 26752 27872
rect 28080 27820 28132 27872
rect 29276 27820 29328 27872
rect 30564 27820 30616 27872
rect 32496 27820 32548 27872
rect 32956 27820 33008 27872
rect 35624 27820 35676 27872
rect 37188 27956 37240 28008
rect 37556 27956 37608 28008
rect 38476 27999 38528 28008
rect 38476 27965 38485 27999
rect 38485 27965 38519 27999
rect 38519 27965 38528 27999
rect 39028 28024 39080 28076
rect 44364 28024 44416 28076
rect 46204 28067 46256 28076
rect 46204 28033 46213 28067
rect 46213 28033 46247 28067
rect 46247 28033 46256 28067
rect 46204 28024 46256 28033
rect 46480 28067 46532 28076
rect 46480 28033 46489 28067
rect 46489 28033 46523 28067
rect 46523 28033 46532 28067
rect 46480 28024 46532 28033
rect 38476 27956 38528 27965
rect 38752 27956 38804 28008
rect 39396 27956 39448 28008
rect 41144 27931 41196 27940
rect 41144 27897 41153 27931
rect 41153 27897 41187 27931
rect 41187 27897 41196 27931
rect 41144 27888 41196 27897
rect 41236 27931 41288 27940
rect 41236 27897 41245 27931
rect 41245 27897 41279 27931
rect 41279 27897 41288 27931
rect 41236 27888 41288 27897
rect 36176 27820 36228 27872
rect 37096 27863 37148 27872
rect 37096 27829 37105 27863
rect 37105 27829 37139 27863
rect 37139 27829 37148 27863
rect 37096 27820 37148 27829
rect 37740 27820 37792 27872
rect 38844 27820 38896 27872
rect 40040 27820 40092 27872
rect 44456 27956 44508 28008
rect 44640 27956 44692 28008
rect 42064 27888 42116 27940
rect 42524 27820 42576 27872
rect 44640 27863 44692 27872
rect 44640 27829 44649 27863
rect 44649 27829 44683 27863
rect 44683 27829 44692 27863
rect 44640 27820 44692 27829
rect 45744 27820 45796 27872
rect 46204 27888 46256 27940
rect 46480 27820 46532 27872
rect 47124 27863 47176 27872
rect 47124 27829 47133 27863
rect 47133 27829 47167 27863
rect 47167 27829 47176 27863
rect 47124 27820 47176 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 15384 27659 15436 27668
rect 15384 27625 15393 27659
rect 15393 27625 15427 27659
rect 15427 27625 15436 27659
rect 15384 27616 15436 27625
rect 16672 27616 16724 27668
rect 19340 27591 19392 27600
rect 19340 27557 19349 27591
rect 19349 27557 19383 27591
rect 19383 27557 19392 27591
rect 19340 27548 19392 27557
rect 14188 27523 14240 27532
rect 14188 27489 14197 27523
rect 14197 27489 14231 27523
rect 14231 27489 14240 27523
rect 14188 27480 14240 27489
rect 14556 27480 14608 27532
rect 15752 27480 15804 27532
rect 17224 27523 17276 27532
rect 17224 27489 17233 27523
rect 17233 27489 17267 27523
rect 17267 27489 17276 27523
rect 17224 27480 17276 27489
rect 17500 27480 17552 27532
rect 18236 27480 18288 27532
rect 19156 27480 19208 27532
rect 24308 27616 24360 27668
rect 26516 27616 26568 27668
rect 29276 27616 29328 27668
rect 31484 27659 31536 27668
rect 31484 27625 31493 27659
rect 31493 27625 31527 27659
rect 31527 27625 31536 27659
rect 31484 27616 31536 27625
rect 31668 27616 31720 27668
rect 32496 27659 32548 27668
rect 32496 27625 32505 27659
rect 32505 27625 32539 27659
rect 32539 27625 32548 27659
rect 32496 27616 32548 27625
rect 33048 27616 33100 27668
rect 34428 27616 34480 27668
rect 23020 27548 23072 27600
rect 25688 27548 25740 27600
rect 28724 27548 28776 27600
rect 30564 27591 30616 27600
rect 30564 27557 30573 27591
rect 30573 27557 30607 27591
rect 30607 27557 30616 27591
rect 30564 27548 30616 27557
rect 38476 27616 38528 27668
rect 38752 27659 38804 27668
rect 38752 27625 38761 27659
rect 38761 27625 38795 27659
rect 38795 27625 38804 27659
rect 38752 27616 38804 27625
rect 38936 27616 38988 27668
rect 39488 27616 39540 27668
rect 41236 27616 41288 27668
rect 35900 27548 35952 27600
rect 21088 27480 21140 27532
rect 21456 27523 21508 27532
rect 21456 27489 21465 27523
rect 21465 27489 21499 27523
rect 21499 27489 21508 27523
rect 21456 27480 21508 27489
rect 22744 27480 22796 27532
rect 24860 27523 24912 27532
rect 24860 27489 24869 27523
rect 24869 27489 24903 27523
rect 24903 27489 24912 27523
rect 24860 27480 24912 27489
rect 16396 27412 16448 27464
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 21732 27455 21784 27464
rect 21732 27421 21741 27455
rect 21741 27421 21775 27455
rect 21775 27421 21784 27455
rect 21732 27412 21784 27421
rect 22652 27412 22704 27464
rect 26424 27480 26476 27532
rect 25504 27412 25556 27464
rect 32220 27480 32272 27532
rect 34152 27523 34204 27532
rect 34152 27489 34161 27523
rect 34161 27489 34195 27523
rect 34195 27489 34204 27523
rect 34152 27480 34204 27489
rect 34336 27523 34388 27532
rect 34336 27489 34345 27523
rect 34345 27489 34379 27523
rect 34379 27489 34388 27523
rect 34336 27480 34388 27489
rect 38108 27480 38160 27532
rect 40960 27548 41012 27600
rect 41788 27591 41840 27600
rect 41788 27557 41797 27591
rect 41797 27557 41831 27591
rect 41831 27557 41840 27591
rect 41788 27548 41840 27557
rect 43904 27616 43956 27668
rect 41972 27548 42024 27600
rect 44456 27548 44508 27600
rect 43260 27480 43312 27532
rect 44364 27480 44416 27532
rect 28356 27412 28408 27464
rect 30472 27455 30524 27464
rect 30472 27421 30481 27455
rect 30481 27421 30515 27455
rect 30515 27421 30524 27455
rect 30472 27412 30524 27421
rect 34428 27455 34480 27464
rect 34428 27421 34437 27455
rect 34437 27421 34471 27455
rect 34471 27421 34480 27455
rect 34428 27412 34480 27421
rect 35716 27455 35768 27464
rect 35716 27421 35725 27455
rect 35725 27421 35759 27455
rect 35759 27421 35768 27455
rect 35716 27412 35768 27421
rect 36360 27455 36412 27464
rect 36360 27421 36369 27455
rect 36369 27421 36403 27455
rect 36403 27421 36412 27455
rect 36360 27412 36412 27421
rect 39580 27412 39632 27464
rect 43720 27412 43772 27464
rect 23848 27344 23900 27396
rect 29184 27344 29236 27396
rect 31024 27387 31076 27396
rect 31024 27353 31033 27387
rect 31033 27353 31067 27387
rect 31067 27353 31076 27387
rect 31024 27344 31076 27353
rect 13360 27276 13412 27328
rect 14372 27319 14424 27328
rect 14372 27285 14381 27319
rect 14381 27285 14415 27319
rect 14415 27285 14424 27319
rect 14372 27276 14424 27285
rect 19892 27276 19944 27328
rect 23480 27319 23532 27328
rect 23480 27285 23489 27319
rect 23489 27285 23523 27319
rect 23523 27285 23532 27319
rect 29092 27319 29144 27328
rect 23480 27276 23532 27285
rect 29092 27285 29101 27319
rect 29101 27285 29135 27319
rect 29135 27285 29144 27319
rect 29092 27276 29144 27285
rect 31116 27276 31168 27328
rect 35256 27319 35308 27328
rect 35256 27285 35265 27319
rect 35265 27285 35299 27319
rect 35299 27285 35308 27319
rect 35256 27276 35308 27285
rect 36728 27319 36780 27328
rect 36728 27285 36737 27319
rect 36737 27285 36771 27319
rect 36771 27285 36780 27319
rect 36728 27276 36780 27285
rect 39396 27276 39448 27328
rect 40132 27319 40184 27328
rect 40132 27285 40141 27319
rect 40141 27285 40175 27319
rect 40175 27285 40184 27319
rect 40132 27276 40184 27285
rect 40500 27319 40552 27328
rect 40500 27285 40509 27319
rect 40509 27285 40543 27319
rect 40543 27285 40552 27319
rect 40500 27276 40552 27285
rect 43260 27276 43312 27328
rect 45836 27276 45888 27328
rect 46204 27548 46256 27600
rect 46388 27455 46440 27464
rect 46388 27421 46397 27455
rect 46397 27421 46431 27455
rect 46431 27421 46440 27455
rect 46388 27412 46440 27421
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 13728 27115 13780 27124
rect 13728 27081 13737 27115
rect 13737 27081 13771 27115
rect 13771 27081 13780 27115
rect 13728 27072 13780 27081
rect 14740 27072 14792 27124
rect 17500 27115 17552 27124
rect 17500 27081 17509 27115
rect 17509 27081 17543 27115
rect 17543 27081 17552 27115
rect 17500 27072 17552 27081
rect 21088 27115 21140 27124
rect 21088 27081 21097 27115
rect 21097 27081 21131 27115
rect 21131 27081 21140 27115
rect 21088 27072 21140 27081
rect 22744 27072 22796 27124
rect 26424 27115 26476 27124
rect 26424 27081 26433 27115
rect 26433 27081 26467 27115
rect 26467 27081 26476 27115
rect 26424 27072 26476 27081
rect 28724 27115 28776 27124
rect 28724 27081 28733 27115
rect 28733 27081 28767 27115
rect 28767 27081 28776 27115
rect 28724 27072 28776 27081
rect 30564 27072 30616 27124
rect 38108 27115 38160 27124
rect 38108 27081 38117 27115
rect 38117 27081 38151 27115
rect 38151 27081 38160 27115
rect 38108 27072 38160 27081
rect 41788 27072 41840 27124
rect 43076 27072 43128 27124
rect 43352 27072 43404 27124
rect 46388 27072 46440 27124
rect 22928 27004 22980 27056
rect 29092 27047 29144 27056
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 17224 26936 17276 26988
rect 18052 26979 18104 26988
rect 18052 26945 18061 26979
rect 18061 26945 18095 26979
rect 18095 26945 18104 26979
rect 18052 26936 18104 26945
rect 19984 26936 20036 26988
rect 21916 26936 21968 26988
rect 14372 26911 14424 26920
rect 14372 26877 14381 26911
rect 14381 26877 14415 26911
rect 14415 26877 14424 26911
rect 14372 26868 14424 26877
rect 14740 26911 14792 26920
rect 14740 26877 14749 26911
rect 14749 26877 14783 26911
rect 14783 26877 14792 26911
rect 14740 26868 14792 26877
rect 15108 26868 15160 26920
rect 16120 26911 16172 26920
rect 16120 26877 16129 26911
rect 16129 26877 16163 26911
rect 16163 26877 16172 26911
rect 16120 26868 16172 26877
rect 16396 26911 16448 26920
rect 16396 26877 16405 26911
rect 16405 26877 16439 26911
rect 16439 26877 16448 26911
rect 16396 26868 16448 26877
rect 16580 26868 16632 26920
rect 21088 26868 21140 26920
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 25044 26911 25096 26920
rect 25044 26877 25053 26911
rect 25053 26877 25087 26911
rect 25087 26877 25096 26911
rect 25044 26868 25096 26877
rect 25504 26911 25556 26920
rect 25504 26877 25513 26911
rect 25513 26877 25547 26911
rect 25547 26877 25556 26911
rect 25504 26868 25556 26877
rect 29092 27013 29101 27047
rect 29101 27013 29135 27047
rect 29135 27013 29144 27047
rect 29092 27004 29144 27013
rect 29276 27004 29328 27056
rect 31024 27004 31076 27056
rect 29828 26979 29880 26988
rect 29828 26945 29837 26979
rect 29837 26945 29871 26979
rect 29871 26945 29880 26979
rect 29828 26936 29880 26945
rect 30932 26979 30984 26988
rect 30932 26945 30941 26979
rect 30941 26945 30975 26979
rect 30975 26945 30984 26979
rect 30932 26936 30984 26945
rect 31576 27004 31628 27056
rect 32404 27004 32456 27056
rect 34152 27004 34204 27056
rect 37464 27004 37516 27056
rect 14188 26775 14240 26784
rect 14188 26741 14197 26775
rect 14197 26741 14231 26775
rect 14231 26741 14240 26775
rect 14188 26732 14240 26741
rect 15752 26732 15804 26784
rect 15936 26775 15988 26784
rect 15936 26741 15945 26775
rect 15945 26741 15979 26775
rect 15979 26741 15988 26775
rect 15936 26732 15988 26741
rect 17776 26775 17828 26784
rect 17776 26741 17785 26775
rect 17785 26741 17819 26775
rect 17819 26741 17828 26775
rect 19340 26800 19392 26852
rect 22008 26800 22060 26852
rect 23020 26843 23072 26852
rect 23020 26809 23029 26843
rect 23029 26809 23063 26843
rect 23063 26809 23072 26843
rect 23020 26800 23072 26809
rect 26976 26800 27028 26852
rect 27896 26911 27948 26920
rect 27896 26877 27905 26911
rect 27905 26877 27939 26911
rect 27939 26877 27948 26911
rect 27896 26868 27948 26877
rect 28264 26868 28316 26920
rect 32956 26868 33008 26920
rect 33600 26936 33652 26988
rect 35256 26936 35308 26988
rect 36728 26979 36780 26988
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 38384 26936 38436 26988
rect 43260 26979 43312 26988
rect 43260 26945 43269 26979
rect 43269 26945 43303 26979
rect 43303 26945 43312 26979
rect 43260 26936 43312 26945
rect 43904 26979 43956 26988
rect 43904 26945 43913 26979
rect 43913 26945 43947 26979
rect 43947 26945 43956 26979
rect 43904 26936 43956 26945
rect 28356 26843 28408 26852
rect 28356 26809 28365 26843
rect 28365 26809 28399 26843
rect 28399 26809 28408 26843
rect 28356 26800 28408 26809
rect 29092 26800 29144 26852
rect 31116 26800 31168 26852
rect 33876 26868 33928 26920
rect 34336 26868 34388 26920
rect 39672 26868 39724 26920
rect 40500 26911 40552 26920
rect 40500 26877 40509 26911
rect 40509 26877 40543 26911
rect 40543 26877 40552 26911
rect 40500 26868 40552 26877
rect 45284 27004 45336 27056
rect 46756 27047 46808 27056
rect 46756 27013 46765 27047
rect 46765 27013 46799 27047
rect 46799 27013 46808 27047
rect 46756 27004 46808 27013
rect 18972 26775 19024 26784
rect 17776 26732 17828 26741
rect 18972 26741 18981 26775
rect 18981 26741 19015 26775
rect 19015 26741 19024 26775
rect 18972 26732 19024 26741
rect 20260 26732 20312 26784
rect 22744 26775 22796 26784
rect 22744 26741 22753 26775
rect 22753 26741 22787 26775
rect 22787 26741 22796 26775
rect 22744 26732 22796 26741
rect 27068 26775 27120 26784
rect 27068 26741 27077 26775
rect 27077 26741 27111 26775
rect 27111 26741 27120 26775
rect 27068 26732 27120 26741
rect 32496 26732 32548 26784
rect 35992 26800 36044 26852
rect 35900 26732 35952 26784
rect 39488 26800 39540 26852
rect 43536 26800 43588 26852
rect 43628 26800 43680 26852
rect 44732 26800 44784 26852
rect 46204 26843 46256 26852
rect 46204 26809 46213 26843
rect 46213 26809 46247 26843
rect 46247 26809 46256 26843
rect 46204 26800 46256 26809
rect 39580 26775 39632 26784
rect 39580 26741 39589 26775
rect 39589 26741 39623 26775
rect 39623 26741 39632 26775
rect 39580 26732 39632 26741
rect 41972 26732 42024 26784
rect 44456 26732 44508 26784
rect 45284 26732 45336 26784
rect 45836 26775 45888 26784
rect 45836 26741 45845 26775
rect 45845 26741 45879 26775
rect 45879 26741 45888 26775
rect 45836 26732 45888 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 14740 26528 14792 26580
rect 16396 26528 16448 26580
rect 17132 26528 17184 26580
rect 18052 26571 18104 26580
rect 18052 26537 18061 26571
rect 18061 26537 18095 26571
rect 18095 26537 18104 26571
rect 18052 26528 18104 26537
rect 19156 26528 19208 26580
rect 19984 26528 20036 26580
rect 21456 26571 21508 26580
rect 21456 26537 21465 26571
rect 21465 26537 21499 26571
rect 21499 26537 21508 26571
rect 21456 26528 21508 26537
rect 21916 26571 21968 26580
rect 21916 26537 21925 26571
rect 21925 26537 21959 26571
rect 21959 26537 21968 26571
rect 21916 26528 21968 26537
rect 28264 26528 28316 26580
rect 28356 26528 28408 26580
rect 29092 26528 29144 26580
rect 29460 26571 29512 26580
rect 29460 26537 29469 26571
rect 29469 26537 29503 26571
rect 29503 26537 29512 26571
rect 29460 26528 29512 26537
rect 30472 26571 30524 26580
rect 30472 26537 30481 26571
rect 30481 26537 30515 26571
rect 30515 26537 30524 26571
rect 30472 26528 30524 26537
rect 30932 26571 30984 26580
rect 30932 26537 30941 26571
rect 30941 26537 30975 26571
rect 30975 26537 30984 26571
rect 30932 26528 30984 26537
rect 32220 26528 32272 26580
rect 14096 26460 14148 26512
rect 15384 26392 15436 26444
rect 15568 26503 15620 26512
rect 15568 26469 15577 26503
rect 15577 26469 15611 26503
rect 15611 26469 15620 26503
rect 15568 26460 15620 26469
rect 18880 26460 18932 26512
rect 22008 26460 22060 26512
rect 33876 26571 33928 26580
rect 33876 26537 33885 26571
rect 33885 26537 33919 26571
rect 33919 26537 33928 26571
rect 33876 26528 33928 26537
rect 34520 26528 34572 26580
rect 35992 26528 36044 26580
rect 17224 26392 17276 26444
rect 21088 26392 21140 26444
rect 21732 26392 21784 26444
rect 22928 26392 22980 26444
rect 23940 26392 23992 26444
rect 24768 26435 24820 26444
rect 24768 26401 24777 26435
rect 24777 26401 24811 26435
rect 24811 26401 24820 26435
rect 24768 26392 24820 26401
rect 25504 26392 25556 26444
rect 27160 26392 27212 26444
rect 28908 26392 28960 26444
rect 30012 26435 30064 26444
rect 18420 26367 18472 26376
rect 18420 26333 18429 26367
rect 18429 26333 18463 26367
rect 18463 26333 18472 26367
rect 18420 26324 18472 26333
rect 18512 26324 18564 26376
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 28080 26324 28132 26376
rect 30012 26401 30021 26435
rect 30021 26401 30055 26435
rect 30055 26401 30064 26435
rect 30012 26392 30064 26401
rect 30932 26392 30984 26444
rect 32036 26392 32088 26444
rect 32128 26392 32180 26444
rect 35624 26460 35676 26512
rect 36084 26503 36136 26512
rect 36084 26469 36093 26503
rect 36093 26469 36127 26503
rect 36127 26469 36136 26503
rect 36084 26460 36136 26469
rect 41144 26528 41196 26580
rect 39672 26503 39724 26512
rect 39672 26469 39681 26503
rect 39681 26469 39715 26503
rect 39715 26469 39724 26503
rect 39672 26460 39724 26469
rect 41972 26460 42024 26512
rect 43904 26528 43956 26580
rect 44364 26528 44416 26580
rect 46204 26528 46256 26580
rect 46848 26528 46900 26580
rect 49516 26528 49568 26580
rect 43536 26503 43588 26512
rect 43536 26469 43545 26503
rect 43545 26469 43579 26503
rect 43579 26469 43588 26503
rect 43536 26460 43588 26469
rect 45836 26503 45888 26512
rect 45836 26469 45845 26503
rect 45845 26469 45879 26503
rect 45879 26469 45888 26503
rect 45836 26460 45888 26469
rect 33324 26392 33376 26444
rect 33968 26392 34020 26444
rect 34428 26392 34480 26444
rect 38016 26392 38068 26444
rect 38844 26392 38896 26444
rect 39396 26435 39448 26444
rect 39396 26401 39405 26435
rect 39405 26401 39439 26435
rect 39439 26401 39448 26435
rect 39396 26392 39448 26401
rect 29552 26324 29604 26376
rect 33048 26324 33100 26376
rect 36360 26367 36412 26376
rect 36360 26333 36369 26367
rect 36369 26333 36403 26367
rect 36403 26333 36412 26367
rect 36360 26324 36412 26333
rect 39212 26324 39264 26376
rect 47124 26392 47176 26444
rect 40684 26324 40736 26376
rect 42524 26324 42576 26376
rect 43628 26324 43680 26376
rect 43720 26367 43772 26376
rect 43720 26333 43729 26367
rect 43729 26333 43763 26367
rect 43763 26333 43772 26367
rect 43720 26324 43772 26333
rect 44824 26324 44876 26376
rect 34152 26256 34204 26308
rect 35992 26256 36044 26308
rect 45560 26256 45612 26308
rect 14372 26231 14424 26240
rect 14372 26197 14381 26231
rect 14381 26197 14415 26231
rect 14415 26197 14424 26231
rect 14372 26188 14424 26197
rect 16396 26188 16448 26240
rect 17960 26188 18012 26240
rect 20076 26188 20128 26240
rect 22192 26231 22244 26240
rect 22192 26197 22201 26231
rect 22201 26197 22235 26231
rect 22235 26197 22244 26231
rect 22192 26188 22244 26197
rect 23296 26231 23348 26240
rect 23296 26197 23305 26231
rect 23305 26197 23339 26231
rect 23339 26197 23348 26231
rect 23296 26188 23348 26197
rect 27528 26188 27580 26240
rect 29000 26188 29052 26240
rect 29276 26188 29328 26240
rect 33232 26188 33284 26240
rect 35624 26231 35676 26240
rect 35624 26197 35633 26231
rect 35633 26197 35667 26231
rect 35667 26197 35676 26231
rect 35624 26188 35676 26197
rect 38384 26231 38436 26240
rect 38384 26197 38393 26231
rect 38393 26197 38427 26231
rect 38427 26197 38436 26231
rect 38384 26188 38436 26197
rect 41052 26188 41104 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 15384 25984 15436 26036
rect 18420 25984 18472 26036
rect 18972 25984 19024 26036
rect 19892 25984 19944 26036
rect 21732 25984 21784 26036
rect 22928 26027 22980 26036
rect 22928 25993 22937 26027
rect 22937 25993 22971 26027
rect 22971 25993 22980 26027
rect 22928 25984 22980 25993
rect 24768 26027 24820 26036
rect 24768 25993 24777 26027
rect 24777 25993 24811 26027
rect 24811 25993 24820 26027
rect 24768 25984 24820 25993
rect 28080 26027 28132 26036
rect 28080 25993 28089 26027
rect 28089 25993 28123 26027
rect 28123 25993 28132 26027
rect 28080 25984 28132 25993
rect 31852 25984 31904 26036
rect 32128 26027 32180 26036
rect 32128 25993 32137 26027
rect 32137 25993 32171 26027
rect 32171 25993 32180 26027
rect 32128 25984 32180 25993
rect 33324 26027 33376 26036
rect 33324 25993 33333 26027
rect 33333 25993 33367 26027
rect 33367 25993 33376 26027
rect 33324 25984 33376 25993
rect 35624 25984 35676 26036
rect 36728 25984 36780 26036
rect 39396 25984 39448 26036
rect 40684 26027 40736 26036
rect 40684 25993 40693 26027
rect 40693 25993 40727 26027
rect 40727 25993 40736 26027
rect 40684 25984 40736 25993
rect 41972 26027 42024 26036
rect 41972 25993 41981 26027
rect 41981 25993 42015 26027
rect 42015 25993 42024 26027
rect 41972 25984 42024 25993
rect 17960 25916 18012 25968
rect 14832 25891 14884 25900
rect 14832 25857 14841 25891
rect 14841 25857 14875 25891
rect 14875 25857 14884 25891
rect 14832 25848 14884 25857
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 20076 25891 20128 25900
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 22192 25916 22244 25968
rect 22008 25848 22060 25900
rect 17776 25823 17828 25832
rect 17776 25789 17785 25823
rect 17785 25789 17819 25823
rect 17819 25789 17828 25823
rect 17776 25780 17828 25789
rect 23664 25780 23716 25832
rect 25596 25891 25648 25900
rect 25596 25857 25605 25891
rect 25605 25857 25639 25891
rect 25639 25857 25648 25891
rect 25596 25848 25648 25857
rect 26056 25848 26108 25900
rect 28908 25916 28960 25968
rect 30012 25916 30064 25968
rect 33692 25916 33744 25968
rect 43536 25984 43588 26036
rect 44824 26027 44876 26036
rect 44824 25993 44833 26027
rect 44833 25993 44867 26027
rect 44867 25993 44876 26027
rect 44824 25984 44876 25993
rect 45836 26027 45888 26036
rect 45836 25993 45845 26027
rect 45845 25993 45879 26027
rect 45879 25993 45888 26027
rect 45836 25984 45888 25993
rect 46204 25984 46256 26036
rect 29000 25848 29052 25900
rect 29736 25848 29788 25900
rect 27160 25780 27212 25832
rect 27988 25780 28040 25832
rect 28724 25823 28776 25832
rect 28724 25789 28733 25823
rect 28733 25789 28767 25823
rect 28767 25789 28776 25823
rect 28724 25780 28776 25789
rect 30196 25780 30248 25832
rect 32036 25780 32088 25832
rect 32680 25823 32732 25832
rect 32680 25789 32689 25823
rect 32689 25789 32723 25823
rect 32723 25789 32732 25823
rect 32680 25780 32732 25789
rect 33048 25780 33100 25832
rect 34796 25848 34848 25900
rect 43628 25916 43680 25968
rect 39580 25848 39632 25900
rect 41052 25891 41104 25900
rect 41052 25857 41061 25891
rect 41061 25857 41095 25891
rect 41095 25857 41104 25891
rect 41052 25848 41104 25857
rect 41696 25891 41748 25900
rect 41696 25857 41705 25891
rect 41705 25857 41739 25891
rect 41739 25857 41748 25891
rect 41696 25848 41748 25857
rect 42064 25848 42116 25900
rect 17224 25712 17276 25764
rect 20260 25712 20312 25764
rect 20352 25712 20404 25764
rect 21732 25755 21784 25764
rect 15476 25644 15528 25696
rect 15752 25687 15804 25696
rect 15752 25653 15761 25687
rect 15761 25653 15795 25687
rect 15795 25653 15804 25687
rect 15752 25644 15804 25653
rect 17316 25644 17368 25696
rect 18972 25687 19024 25696
rect 18972 25653 18981 25687
rect 18981 25653 19015 25687
rect 19015 25653 19024 25687
rect 18972 25644 19024 25653
rect 21088 25687 21140 25696
rect 21088 25653 21097 25687
rect 21097 25653 21131 25687
rect 21131 25653 21140 25687
rect 21088 25644 21140 25653
rect 21732 25721 21741 25755
rect 21741 25721 21775 25755
rect 21775 25721 21784 25755
rect 21732 25712 21784 25721
rect 22468 25712 22520 25764
rect 25136 25712 25188 25764
rect 26884 25712 26936 25764
rect 28816 25712 28868 25764
rect 28908 25712 28960 25764
rect 29460 25755 29512 25764
rect 29460 25721 29469 25755
rect 29469 25721 29503 25755
rect 29503 25721 29512 25755
rect 29460 25712 29512 25721
rect 30012 25755 30064 25764
rect 30012 25721 30021 25755
rect 30021 25721 30055 25755
rect 30055 25721 30064 25755
rect 30012 25712 30064 25721
rect 38476 25823 38528 25832
rect 26700 25644 26752 25696
rect 30932 25644 30984 25696
rect 31668 25644 31720 25696
rect 32128 25644 32180 25696
rect 34520 25644 34572 25696
rect 34796 25644 34848 25696
rect 35348 25687 35400 25696
rect 35348 25653 35357 25687
rect 35357 25653 35391 25687
rect 35391 25653 35400 25687
rect 35348 25644 35400 25653
rect 35992 25687 36044 25696
rect 35992 25653 36001 25687
rect 36001 25653 36035 25687
rect 36035 25653 36044 25687
rect 35992 25644 36044 25653
rect 38476 25789 38485 25823
rect 38485 25789 38519 25823
rect 38519 25789 38528 25823
rect 38476 25780 38528 25789
rect 38752 25823 38804 25832
rect 38752 25789 38761 25823
rect 38761 25789 38795 25823
rect 38795 25789 38804 25823
rect 38752 25780 38804 25789
rect 40132 25712 40184 25764
rect 41052 25712 41104 25764
rect 43536 25755 43588 25764
rect 43536 25721 43545 25755
rect 43545 25721 43579 25755
rect 43579 25721 43588 25755
rect 43536 25712 43588 25721
rect 44732 25780 44784 25832
rect 45376 25823 45428 25832
rect 45376 25789 45385 25823
rect 45385 25789 45419 25823
rect 45419 25789 45428 25823
rect 45376 25780 45428 25789
rect 45468 25780 45520 25832
rect 47032 25780 47084 25832
rect 37280 25644 37332 25696
rect 38016 25687 38068 25696
rect 38016 25653 38025 25687
rect 38025 25653 38059 25687
rect 38059 25653 38068 25687
rect 38016 25644 38068 25653
rect 38844 25644 38896 25696
rect 43352 25644 43404 25696
rect 46572 25644 46624 25696
rect 46664 25644 46716 25696
rect 47124 25644 47176 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 14832 25483 14884 25492
rect 14832 25449 14841 25483
rect 14841 25449 14875 25483
rect 14875 25449 14884 25483
rect 14832 25440 14884 25449
rect 15752 25440 15804 25492
rect 16212 25440 16264 25492
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 23756 25440 23808 25492
rect 25504 25440 25556 25492
rect 25596 25440 25648 25492
rect 26884 25483 26936 25492
rect 26884 25449 26893 25483
rect 26893 25449 26927 25483
rect 26927 25449 26936 25483
rect 26884 25440 26936 25449
rect 29736 25483 29788 25492
rect 29736 25449 29745 25483
rect 29745 25449 29779 25483
rect 29779 25449 29788 25483
rect 29736 25440 29788 25449
rect 31668 25440 31720 25492
rect 15476 25372 15528 25424
rect 16396 25372 16448 25424
rect 17132 25372 17184 25424
rect 17316 25372 17368 25424
rect 18696 25415 18748 25424
rect 18696 25381 18705 25415
rect 18705 25381 18739 25415
rect 18739 25381 18748 25415
rect 18696 25372 18748 25381
rect 18972 25372 19024 25424
rect 21088 25372 21140 25424
rect 21916 25372 21968 25424
rect 22192 25372 22244 25424
rect 22744 25415 22796 25424
rect 22744 25381 22753 25415
rect 22753 25381 22787 25415
rect 22787 25381 22796 25415
rect 22744 25372 22796 25381
rect 25044 25415 25096 25424
rect 25044 25381 25053 25415
rect 25053 25381 25087 25415
rect 25087 25381 25096 25415
rect 25044 25372 25096 25381
rect 28908 25415 28960 25424
rect 28908 25381 28917 25415
rect 28917 25381 28951 25415
rect 28951 25381 28960 25415
rect 28908 25372 28960 25381
rect 30564 25372 30616 25424
rect 14924 25304 14976 25356
rect 15936 25304 15988 25356
rect 17868 25304 17920 25356
rect 18512 25304 18564 25356
rect 19432 25304 19484 25356
rect 21548 25304 21600 25356
rect 26516 25347 26568 25356
rect 26516 25313 26525 25347
rect 26525 25313 26559 25347
rect 26559 25313 26568 25347
rect 26516 25304 26568 25313
rect 17408 25236 17460 25288
rect 18420 25236 18472 25288
rect 20352 25236 20404 25288
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 23940 25236 23992 25288
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 28816 25279 28868 25288
rect 28816 25245 28825 25279
rect 28825 25245 28859 25279
rect 28859 25245 28868 25279
rect 28816 25236 28868 25245
rect 30380 25236 30432 25288
rect 30564 25279 30616 25288
rect 30564 25245 30573 25279
rect 30573 25245 30607 25279
rect 30607 25245 30616 25279
rect 30564 25236 30616 25245
rect 34428 25440 34480 25492
rect 34796 25440 34848 25492
rect 36084 25483 36136 25492
rect 36084 25449 36093 25483
rect 36093 25449 36127 25483
rect 36127 25449 36136 25483
rect 36084 25440 36136 25449
rect 38384 25440 38436 25492
rect 41052 25483 41104 25492
rect 41052 25449 41061 25483
rect 41061 25449 41095 25483
rect 41095 25449 41104 25483
rect 41052 25440 41104 25449
rect 32312 25415 32364 25424
rect 32312 25381 32321 25415
rect 32321 25381 32355 25415
rect 32355 25381 32364 25415
rect 32312 25372 32364 25381
rect 34612 25372 34664 25424
rect 35900 25372 35952 25424
rect 37188 25372 37240 25424
rect 38292 25372 38344 25424
rect 41788 25415 41840 25424
rect 34244 25304 34296 25356
rect 36268 25304 36320 25356
rect 37832 25304 37884 25356
rect 41788 25381 41797 25415
rect 41797 25381 41831 25415
rect 41831 25381 41840 25415
rect 41788 25372 41840 25381
rect 43536 25415 43588 25424
rect 43536 25381 43545 25415
rect 43545 25381 43579 25415
rect 43579 25381 43588 25415
rect 43536 25372 43588 25381
rect 46296 25372 46348 25424
rect 39304 25304 39356 25356
rect 39396 25304 39448 25356
rect 32496 25279 32548 25288
rect 16120 25168 16172 25220
rect 32496 25245 32505 25279
rect 32505 25245 32539 25279
rect 32539 25245 32548 25279
rect 32496 25236 32548 25245
rect 35532 25236 35584 25288
rect 38108 25236 38160 25288
rect 38476 25236 38528 25288
rect 39948 25279 40000 25288
rect 39948 25245 39957 25279
rect 39957 25245 39991 25279
rect 39991 25245 40000 25279
rect 39948 25236 40000 25245
rect 41696 25279 41748 25288
rect 41696 25245 41705 25279
rect 41705 25245 41739 25279
rect 41739 25245 41748 25279
rect 41696 25236 41748 25245
rect 41972 25279 42024 25288
rect 41972 25245 41981 25279
rect 41981 25245 42015 25279
rect 42015 25245 42024 25279
rect 43444 25279 43496 25288
rect 41972 25236 42024 25245
rect 35440 25211 35492 25220
rect 35440 25177 35449 25211
rect 35449 25177 35483 25211
rect 35483 25177 35492 25211
rect 35440 25168 35492 25177
rect 38384 25168 38436 25220
rect 43444 25245 43453 25279
rect 43453 25245 43487 25279
rect 43487 25245 43496 25279
rect 43444 25236 43496 25245
rect 45284 25279 45336 25288
rect 43628 25168 43680 25220
rect 45284 25245 45293 25279
rect 45293 25245 45327 25279
rect 45327 25245 45336 25279
rect 45284 25236 45336 25245
rect 45560 25279 45612 25288
rect 45560 25245 45569 25279
rect 45569 25245 45603 25279
rect 45603 25245 45612 25279
rect 45560 25236 45612 25245
rect 46204 25236 46256 25288
rect 16304 25100 16356 25152
rect 18420 25143 18472 25152
rect 18420 25109 18429 25143
rect 18429 25109 18463 25143
rect 18463 25109 18472 25143
rect 18420 25100 18472 25109
rect 19984 25100 20036 25152
rect 27436 25143 27488 25152
rect 27436 25109 27445 25143
rect 27445 25109 27479 25143
rect 27479 25109 27488 25143
rect 27436 25100 27488 25109
rect 30656 25100 30708 25152
rect 32312 25100 32364 25152
rect 36912 25143 36964 25152
rect 36912 25109 36921 25143
rect 36921 25109 36955 25143
rect 36955 25109 36964 25143
rect 36912 25100 36964 25109
rect 44548 25143 44600 25152
rect 44548 25109 44557 25143
rect 44557 25109 44591 25143
rect 44591 25109 44600 25143
rect 44548 25100 44600 25109
rect 46296 25143 46348 25152
rect 46296 25109 46305 25143
rect 46305 25109 46339 25143
rect 46339 25109 46348 25143
rect 46296 25100 46348 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 14924 24939 14976 24948
rect 14924 24905 14933 24939
rect 14933 24905 14967 24939
rect 14967 24905 14976 24939
rect 14924 24896 14976 24905
rect 17132 24939 17184 24948
rect 17132 24905 17141 24939
rect 17141 24905 17175 24939
rect 17175 24905 17184 24939
rect 17132 24896 17184 24905
rect 17408 24939 17460 24948
rect 17408 24905 17417 24939
rect 17417 24905 17451 24939
rect 17451 24905 17460 24939
rect 17408 24896 17460 24905
rect 18604 24896 18656 24948
rect 18696 24896 18748 24948
rect 19892 24896 19944 24948
rect 20076 24896 20128 24948
rect 23296 24896 23348 24948
rect 25136 24939 25188 24948
rect 25136 24905 25145 24939
rect 25145 24905 25179 24939
rect 25179 24905 25188 24939
rect 25136 24896 25188 24905
rect 26516 24896 26568 24948
rect 28908 24896 28960 24948
rect 30656 24896 30708 24948
rect 31116 24896 31168 24948
rect 32312 24896 32364 24948
rect 33324 24896 33376 24948
rect 34612 24939 34664 24948
rect 34612 24905 34621 24939
rect 34621 24905 34655 24939
rect 34655 24905 34664 24939
rect 34612 24896 34664 24905
rect 37832 24939 37884 24948
rect 37832 24905 37841 24939
rect 37841 24905 37875 24939
rect 37875 24905 37884 24939
rect 37832 24896 37884 24905
rect 39304 24939 39356 24948
rect 39304 24905 39313 24939
rect 39313 24905 39347 24939
rect 39347 24905 39356 24939
rect 39304 24896 39356 24905
rect 39396 24896 39448 24948
rect 43444 24896 43496 24948
rect 45560 24896 45612 24948
rect 16764 24828 16816 24880
rect 17868 24828 17920 24880
rect 18880 24828 18932 24880
rect 18604 24760 18656 24812
rect 19156 24760 19208 24812
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 23756 24803 23808 24812
rect 22376 24760 22428 24769
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 23940 24760 23992 24812
rect 25044 24828 25096 24880
rect 30012 24828 30064 24880
rect 32496 24828 32548 24880
rect 32680 24828 32732 24880
rect 36268 24828 36320 24880
rect 39212 24828 39264 24880
rect 25320 24803 25372 24812
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 25320 24760 25372 24769
rect 25596 24760 25648 24812
rect 27252 24760 27304 24812
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 30380 24760 30432 24769
rect 31668 24803 31720 24812
rect 31668 24769 31677 24803
rect 31677 24769 31711 24803
rect 31711 24769 31720 24803
rect 31668 24760 31720 24769
rect 32128 24760 32180 24812
rect 33232 24803 33284 24812
rect 33232 24769 33241 24803
rect 33241 24769 33275 24803
rect 33275 24769 33284 24803
rect 33232 24760 33284 24769
rect 33508 24803 33560 24812
rect 33508 24769 33517 24803
rect 33517 24769 33551 24803
rect 33551 24769 33560 24803
rect 33508 24760 33560 24769
rect 34796 24760 34848 24812
rect 35440 24803 35492 24812
rect 35440 24769 35449 24803
rect 35449 24769 35483 24803
rect 35483 24769 35492 24803
rect 35440 24760 35492 24769
rect 37464 24803 37516 24812
rect 37464 24769 37473 24803
rect 37473 24769 37507 24803
rect 37507 24769 37516 24803
rect 37464 24760 37516 24769
rect 37648 24760 37700 24812
rect 38384 24803 38436 24812
rect 38384 24769 38393 24803
rect 38393 24769 38427 24803
rect 38427 24769 38436 24803
rect 38384 24760 38436 24769
rect 38476 24760 38528 24812
rect 43996 24828 44048 24880
rect 46756 24871 46808 24880
rect 41972 24760 42024 24812
rect 44548 24803 44600 24812
rect 44548 24769 44557 24803
rect 44557 24769 44591 24803
rect 44591 24769 44600 24803
rect 44548 24760 44600 24769
rect 46756 24837 46765 24871
rect 46765 24837 46799 24871
rect 46799 24837 46808 24871
rect 46756 24828 46808 24837
rect 46204 24803 46256 24812
rect 46204 24769 46213 24803
rect 46213 24769 46247 24803
rect 46247 24769 46256 24803
rect 46204 24760 46256 24769
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 16120 24667 16172 24676
rect 16120 24633 16129 24667
rect 16129 24633 16163 24667
rect 16163 24633 16172 24667
rect 16120 24624 16172 24633
rect 16212 24667 16264 24676
rect 16212 24633 16221 24667
rect 16221 24633 16255 24667
rect 16255 24633 16264 24667
rect 16212 24624 16264 24633
rect 18420 24624 18472 24676
rect 19340 24624 19392 24676
rect 19984 24667 20036 24676
rect 16028 24556 16080 24608
rect 18144 24556 18196 24608
rect 19984 24633 19993 24667
rect 19993 24633 20027 24667
rect 20027 24633 20036 24667
rect 19984 24624 20036 24633
rect 20076 24667 20128 24676
rect 20076 24633 20085 24667
rect 20085 24633 20119 24667
rect 20119 24633 20128 24667
rect 20628 24667 20680 24676
rect 20076 24624 20128 24633
rect 20628 24633 20637 24667
rect 20637 24633 20671 24667
rect 20671 24633 20680 24667
rect 20628 24624 20680 24633
rect 21456 24624 21508 24676
rect 22192 24667 22244 24676
rect 22192 24633 22201 24667
rect 22201 24633 22235 24667
rect 22235 24633 22244 24667
rect 22192 24624 22244 24633
rect 23296 24624 23348 24676
rect 21548 24599 21600 24608
rect 21548 24565 21557 24599
rect 21557 24565 21591 24599
rect 21591 24565 21600 24599
rect 21548 24556 21600 24565
rect 25136 24624 25188 24676
rect 42432 24692 42484 24744
rect 27160 24667 27212 24676
rect 27160 24633 27169 24667
rect 27169 24633 27203 24667
rect 27203 24633 27212 24667
rect 27160 24624 27212 24633
rect 26884 24556 26936 24608
rect 27436 24624 27488 24676
rect 30104 24667 30156 24676
rect 30104 24633 30113 24667
rect 30113 24633 30147 24667
rect 30147 24633 30156 24667
rect 30104 24624 30156 24633
rect 32312 24624 32364 24676
rect 33324 24667 33376 24676
rect 33324 24633 33333 24667
rect 33333 24633 33367 24667
rect 33367 24633 33376 24667
rect 33324 24624 33376 24633
rect 34244 24667 34296 24676
rect 34244 24633 34253 24667
rect 34253 24633 34287 24667
rect 34287 24633 34296 24667
rect 34244 24624 34296 24633
rect 35992 24667 36044 24676
rect 35992 24633 36001 24667
rect 36001 24633 36035 24667
rect 36035 24633 36044 24667
rect 35992 24624 36044 24633
rect 36636 24624 36688 24676
rect 36912 24667 36964 24676
rect 36912 24633 36921 24667
rect 36921 24633 36955 24667
rect 36955 24633 36964 24667
rect 36912 24624 36964 24633
rect 40960 24667 41012 24676
rect 40960 24633 40969 24667
rect 40969 24633 41003 24667
rect 41003 24633 41012 24667
rect 40960 24624 41012 24633
rect 41788 24599 41840 24608
rect 41788 24565 41797 24599
rect 41797 24565 41831 24599
rect 41831 24565 41840 24599
rect 41788 24556 41840 24565
rect 42064 24556 42116 24608
rect 46296 24667 46348 24676
rect 43260 24599 43312 24608
rect 43260 24565 43269 24599
rect 43269 24565 43303 24599
rect 43303 24565 43312 24599
rect 43260 24556 43312 24565
rect 43536 24599 43588 24608
rect 43536 24565 43545 24599
rect 43545 24565 43579 24599
rect 43579 24565 43588 24599
rect 43536 24556 43588 24565
rect 46296 24633 46305 24667
rect 46305 24633 46339 24667
rect 46339 24633 46348 24667
rect 46296 24624 46348 24633
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 18144 24352 18196 24404
rect 18236 24352 18288 24404
rect 18972 24352 19024 24404
rect 19064 24352 19116 24404
rect 16304 24284 16356 24336
rect 16764 24327 16816 24336
rect 16764 24293 16773 24327
rect 16773 24293 16807 24327
rect 16807 24293 16816 24327
rect 16764 24284 16816 24293
rect 17868 24216 17920 24268
rect 22468 24352 22520 24404
rect 22652 24352 22704 24404
rect 25320 24352 25372 24404
rect 27160 24352 27212 24404
rect 28540 24395 28592 24404
rect 28540 24361 28549 24395
rect 28549 24361 28583 24395
rect 28583 24361 28592 24395
rect 28540 24352 28592 24361
rect 28816 24352 28868 24404
rect 30564 24395 30616 24404
rect 30564 24361 30573 24395
rect 30573 24361 30607 24395
rect 30607 24361 30616 24395
rect 30564 24352 30616 24361
rect 31668 24395 31720 24404
rect 31668 24361 31677 24395
rect 31677 24361 31711 24395
rect 31711 24361 31720 24395
rect 31668 24352 31720 24361
rect 33232 24395 33284 24404
rect 33232 24361 33241 24395
rect 33241 24361 33275 24395
rect 33275 24361 33284 24395
rect 33232 24352 33284 24361
rect 35532 24395 35584 24404
rect 35532 24361 35541 24395
rect 35541 24361 35575 24395
rect 35575 24361 35584 24395
rect 35532 24352 35584 24361
rect 41788 24352 41840 24404
rect 43536 24352 43588 24404
rect 19340 24327 19392 24336
rect 19340 24293 19349 24327
rect 19349 24293 19383 24327
rect 19383 24293 19392 24327
rect 19340 24284 19392 24293
rect 20076 24284 20128 24336
rect 21824 24327 21876 24336
rect 21824 24293 21833 24327
rect 21833 24293 21867 24327
rect 21867 24293 21876 24327
rect 21824 24284 21876 24293
rect 22192 24284 22244 24336
rect 23480 24327 23532 24336
rect 23480 24293 23489 24327
rect 23489 24293 23523 24327
rect 23523 24293 23532 24327
rect 23480 24284 23532 24293
rect 25412 24284 25464 24336
rect 26700 24327 26752 24336
rect 26700 24293 26709 24327
rect 26709 24293 26743 24327
rect 26743 24293 26752 24327
rect 26700 24284 26752 24293
rect 27252 24327 27304 24336
rect 27252 24293 27261 24327
rect 27261 24293 27295 24327
rect 27295 24293 27304 24327
rect 27252 24284 27304 24293
rect 29276 24284 29328 24336
rect 32220 24327 32272 24336
rect 32220 24293 32229 24327
rect 32229 24293 32263 24327
rect 32263 24293 32272 24327
rect 32220 24284 32272 24293
rect 32312 24327 32364 24336
rect 32312 24293 32321 24327
rect 32321 24293 32355 24327
rect 32355 24293 32364 24327
rect 32312 24284 32364 24293
rect 33508 24284 33560 24336
rect 34520 24284 34572 24336
rect 35900 24284 35952 24336
rect 36452 24284 36504 24336
rect 39488 24284 39540 24336
rect 40316 24284 40368 24336
rect 42064 24284 42116 24336
rect 44364 24284 44416 24336
rect 45284 24352 45336 24404
rect 45468 24395 45520 24404
rect 45468 24361 45477 24395
rect 45477 24361 45511 24395
rect 45511 24361 45520 24395
rect 45468 24352 45520 24361
rect 45836 24284 45888 24336
rect 46296 24284 46348 24336
rect 27712 24216 27764 24268
rect 30196 24216 30248 24268
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 17040 24148 17092 24200
rect 19248 24191 19300 24200
rect 19248 24157 19257 24191
rect 19257 24157 19291 24191
rect 19291 24157 19300 24191
rect 19248 24148 19300 24157
rect 19984 24148 20036 24200
rect 20168 24148 20220 24200
rect 22744 24148 22796 24200
rect 23388 24191 23440 24200
rect 23388 24157 23397 24191
rect 23397 24157 23431 24191
rect 23431 24157 23440 24191
rect 23388 24148 23440 24157
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 16028 24080 16080 24132
rect 22928 24080 22980 24132
rect 23940 24123 23992 24132
rect 23940 24089 23949 24123
rect 23949 24089 23983 24123
rect 23983 24089 23992 24123
rect 23940 24080 23992 24089
rect 25872 24148 25924 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 31300 24216 31352 24268
rect 26332 24080 26384 24132
rect 18144 24012 18196 24064
rect 19708 24012 19760 24064
rect 29092 24055 29144 24064
rect 29092 24021 29101 24055
rect 29101 24021 29135 24055
rect 29135 24021 29144 24055
rect 29092 24012 29144 24021
rect 34060 24012 34112 24064
rect 37004 24216 37056 24268
rect 37924 24259 37976 24268
rect 37924 24225 37933 24259
rect 37933 24225 37967 24259
rect 37967 24225 37976 24259
rect 37924 24216 37976 24225
rect 38384 24216 38436 24268
rect 39396 24216 39448 24268
rect 36176 24191 36228 24200
rect 36176 24157 36185 24191
rect 36185 24157 36219 24191
rect 36219 24157 36228 24191
rect 36176 24148 36228 24157
rect 36636 24148 36688 24200
rect 39488 24191 39540 24200
rect 39488 24157 39497 24191
rect 39497 24157 39531 24191
rect 39531 24157 39540 24191
rect 39488 24148 39540 24157
rect 41236 24191 41288 24200
rect 41236 24157 41245 24191
rect 41245 24157 41279 24191
rect 41279 24157 41288 24191
rect 41236 24148 41288 24157
rect 44272 24191 44324 24200
rect 44272 24157 44281 24191
rect 44281 24157 44315 24191
rect 44315 24157 44324 24191
rect 44272 24148 44324 24157
rect 46112 24191 46164 24200
rect 46112 24157 46121 24191
rect 46121 24157 46155 24191
rect 46155 24157 46164 24191
rect 46112 24148 46164 24157
rect 46480 24191 46532 24200
rect 46480 24157 46489 24191
rect 46489 24157 46523 24191
rect 46523 24157 46532 24191
rect 46480 24148 46532 24157
rect 35256 24123 35308 24132
rect 35256 24089 35265 24123
rect 35265 24089 35299 24123
rect 35299 24089 35308 24123
rect 35256 24080 35308 24089
rect 35900 24055 35952 24064
rect 35900 24021 35909 24055
rect 35909 24021 35943 24055
rect 35943 24021 35952 24055
rect 35900 24012 35952 24021
rect 37280 24080 37332 24132
rect 36912 24012 36964 24064
rect 40868 24055 40920 24064
rect 40868 24021 40877 24055
rect 40877 24021 40911 24055
rect 40911 24021 40920 24055
rect 40868 24012 40920 24021
rect 42432 24055 42484 24064
rect 42432 24021 42441 24055
rect 42441 24021 42475 24055
rect 42475 24021 42484 24055
rect 42432 24012 42484 24021
rect 42892 24012 42944 24064
rect 44824 24012 44876 24064
rect 47032 24012 47084 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 16304 23808 16356 23860
rect 17868 23851 17920 23860
rect 17868 23817 17877 23851
rect 17877 23817 17911 23851
rect 17911 23817 17920 23851
rect 17868 23808 17920 23817
rect 19340 23808 19392 23860
rect 20260 23808 20312 23860
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 22192 23808 22244 23860
rect 22652 23808 22704 23860
rect 17040 23783 17092 23792
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 19984 23740 20036 23792
rect 14464 23672 14516 23724
rect 16672 23672 16724 23724
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 19064 23672 19116 23724
rect 19708 23715 19760 23724
rect 19708 23681 19717 23715
rect 19717 23681 19751 23715
rect 19751 23681 19760 23715
rect 19708 23672 19760 23681
rect 19800 23672 19852 23724
rect 15844 23604 15896 23656
rect 15476 23536 15528 23588
rect 17500 23579 17552 23588
rect 17500 23545 17509 23579
rect 17509 23545 17543 23579
rect 17543 23545 17552 23579
rect 18236 23579 18288 23588
rect 17500 23536 17552 23545
rect 18236 23545 18245 23579
rect 18245 23545 18279 23579
rect 18279 23545 18288 23579
rect 18236 23536 18288 23545
rect 15200 23468 15252 23520
rect 19708 23536 19760 23588
rect 20168 23536 20220 23588
rect 21364 23604 21416 23656
rect 22836 23808 22888 23860
rect 23388 23808 23440 23860
rect 25412 23808 25464 23860
rect 25872 23851 25924 23860
rect 25872 23817 25881 23851
rect 25881 23817 25915 23851
rect 25915 23817 25924 23851
rect 25872 23808 25924 23817
rect 26332 23808 26384 23860
rect 26700 23808 26752 23860
rect 26884 23808 26936 23860
rect 28540 23808 28592 23860
rect 29092 23851 29144 23860
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 30104 23808 30156 23860
rect 31300 23851 31352 23860
rect 31300 23817 31309 23851
rect 31309 23817 31343 23851
rect 31343 23817 31352 23851
rect 31300 23808 31352 23817
rect 32220 23808 32272 23860
rect 36636 23808 36688 23860
rect 36912 23808 36964 23860
rect 37924 23851 37976 23860
rect 37924 23817 37933 23851
rect 37933 23817 37967 23851
rect 37967 23817 37976 23851
rect 37924 23808 37976 23817
rect 38384 23851 38436 23860
rect 38384 23817 38393 23851
rect 38393 23817 38427 23851
rect 38427 23817 38436 23851
rect 38384 23808 38436 23817
rect 41236 23808 41288 23860
rect 43260 23808 43312 23860
rect 44548 23808 44600 23860
rect 45836 23851 45888 23860
rect 45836 23817 45845 23851
rect 45845 23817 45879 23851
rect 45879 23817 45888 23851
rect 45836 23808 45888 23817
rect 22928 23740 22980 23792
rect 23480 23672 23532 23724
rect 24952 23740 25004 23792
rect 28172 23715 28224 23724
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 29828 23715 29880 23724
rect 29828 23681 29837 23715
rect 29837 23681 29871 23715
rect 29871 23681 29880 23715
rect 29828 23672 29880 23681
rect 30196 23672 30248 23724
rect 26332 23604 26384 23656
rect 27344 23604 27396 23656
rect 28264 23604 28316 23656
rect 34244 23740 34296 23792
rect 32312 23672 32364 23724
rect 35900 23740 35952 23792
rect 35992 23740 36044 23792
rect 35348 23715 35400 23724
rect 35348 23681 35357 23715
rect 35357 23681 35391 23715
rect 35391 23681 35400 23715
rect 35348 23672 35400 23681
rect 31852 23604 31904 23656
rect 33324 23604 33376 23656
rect 19432 23468 19484 23520
rect 23848 23536 23900 23588
rect 24124 23536 24176 23588
rect 27712 23536 27764 23588
rect 29368 23579 29420 23588
rect 29368 23545 29377 23579
rect 29377 23545 29411 23579
rect 29411 23545 29420 23579
rect 29368 23536 29420 23545
rect 26332 23468 26384 23520
rect 29092 23468 29144 23520
rect 33600 23536 33652 23588
rect 29644 23468 29696 23520
rect 34520 23468 34572 23520
rect 35256 23536 35308 23588
rect 40040 23740 40092 23792
rect 40868 23740 40920 23792
rect 46112 23740 46164 23792
rect 37280 23672 37332 23724
rect 38476 23672 38528 23724
rect 39948 23672 40000 23724
rect 40684 23715 40736 23724
rect 40684 23681 40693 23715
rect 40693 23681 40727 23715
rect 40727 23681 40736 23715
rect 40684 23672 40736 23681
rect 43352 23672 43404 23724
rect 43628 23715 43680 23724
rect 43628 23681 43637 23715
rect 43637 23681 43671 23715
rect 43671 23681 43680 23715
rect 43628 23672 43680 23681
rect 45376 23672 45428 23724
rect 45836 23672 45888 23724
rect 38660 23604 38712 23656
rect 39396 23647 39448 23656
rect 39396 23613 39405 23647
rect 39405 23613 39439 23647
rect 39439 23613 39448 23647
rect 39396 23604 39448 23613
rect 42432 23604 42484 23656
rect 45100 23604 45152 23656
rect 45652 23604 45704 23656
rect 36912 23579 36964 23588
rect 36912 23545 36921 23579
rect 36921 23545 36955 23579
rect 36955 23545 36964 23579
rect 36912 23536 36964 23545
rect 37004 23579 37056 23588
rect 37004 23545 37013 23579
rect 37013 23545 37047 23579
rect 37047 23545 37056 23579
rect 37004 23536 37056 23545
rect 38660 23511 38712 23520
rect 38660 23477 38669 23511
rect 38669 23477 38703 23511
rect 38703 23477 38712 23511
rect 38660 23468 38712 23477
rect 40316 23511 40368 23520
rect 40316 23477 40325 23511
rect 40325 23477 40359 23511
rect 40359 23477 40368 23511
rect 43352 23579 43404 23588
rect 43352 23545 43361 23579
rect 43361 23545 43395 23579
rect 43395 23545 43404 23579
rect 43352 23536 43404 23545
rect 40316 23468 40368 23477
rect 44364 23468 44416 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 14464 23264 14516 23316
rect 19248 23307 19300 23316
rect 15844 23239 15896 23248
rect 15844 23205 15853 23239
rect 15853 23205 15887 23239
rect 15887 23205 15896 23239
rect 15844 23196 15896 23205
rect 16120 23196 16172 23248
rect 18328 23196 18380 23248
rect 19248 23273 19257 23307
rect 19257 23273 19291 23307
rect 19291 23273 19300 23307
rect 19248 23264 19300 23273
rect 21824 23307 21876 23316
rect 21824 23273 21833 23307
rect 21833 23273 21867 23307
rect 21867 23273 21876 23307
rect 21824 23264 21876 23273
rect 23388 23307 23440 23316
rect 23388 23273 23397 23307
rect 23397 23273 23431 23307
rect 23431 23273 23440 23307
rect 23388 23264 23440 23273
rect 24952 23307 25004 23316
rect 24952 23273 24961 23307
rect 24961 23273 24995 23307
rect 24995 23273 25004 23307
rect 24952 23264 25004 23273
rect 28172 23307 28224 23316
rect 28172 23273 28181 23307
rect 28181 23273 28215 23307
rect 28215 23273 28224 23307
rect 28172 23264 28224 23273
rect 20628 23196 20680 23248
rect 23296 23196 23348 23248
rect 26424 23196 26476 23248
rect 26608 23196 26660 23248
rect 27252 23239 27304 23248
rect 27252 23205 27261 23239
rect 27261 23205 27295 23239
rect 27295 23205 27304 23239
rect 27252 23196 27304 23205
rect 27528 23196 27580 23248
rect 29552 23239 29604 23248
rect 29552 23205 29561 23239
rect 29561 23205 29595 23239
rect 29595 23205 29604 23239
rect 29552 23196 29604 23205
rect 29644 23239 29696 23248
rect 29644 23205 29653 23239
rect 29653 23205 29687 23239
rect 29687 23205 29696 23239
rect 29644 23196 29696 23205
rect 31852 23196 31904 23248
rect 32496 23196 32548 23248
rect 33508 23264 33560 23316
rect 34060 23307 34112 23316
rect 34060 23273 34069 23307
rect 34069 23273 34103 23307
rect 34103 23273 34112 23307
rect 34060 23264 34112 23273
rect 35256 23264 35308 23316
rect 36176 23307 36228 23316
rect 36176 23273 36185 23307
rect 36185 23273 36219 23307
rect 36219 23273 36228 23307
rect 36176 23264 36228 23273
rect 36912 23264 36964 23316
rect 37096 23264 37148 23316
rect 14280 23128 14332 23180
rect 19616 23171 19668 23180
rect 19616 23137 19625 23171
rect 19625 23137 19659 23171
rect 19659 23137 19668 23171
rect 19616 23128 19668 23137
rect 21364 23171 21416 23180
rect 21364 23137 21373 23171
rect 21373 23137 21407 23171
rect 21407 23137 21416 23171
rect 21364 23128 21416 23137
rect 24860 23128 24912 23180
rect 25044 23128 25096 23180
rect 26056 23128 26108 23180
rect 33876 23128 33928 23180
rect 38844 23196 38896 23248
rect 39488 23264 39540 23316
rect 40684 23307 40736 23316
rect 40684 23273 40693 23307
rect 40693 23273 40727 23307
rect 40727 23273 40736 23307
rect 40684 23264 40736 23273
rect 44272 23307 44324 23316
rect 41236 23196 41288 23248
rect 44272 23273 44281 23307
rect 44281 23273 44315 23307
rect 44315 23273 44324 23307
rect 44272 23264 44324 23273
rect 45468 23264 45520 23316
rect 46112 23307 46164 23316
rect 46112 23273 46121 23307
rect 46121 23273 46155 23307
rect 46155 23273 46164 23307
rect 46112 23264 46164 23273
rect 34152 23128 34204 23180
rect 35992 23128 36044 23180
rect 36636 23128 36688 23180
rect 37740 23128 37792 23180
rect 39304 23171 39356 23180
rect 39304 23137 39313 23171
rect 39313 23137 39347 23171
rect 39347 23137 39356 23171
rect 39304 23128 39356 23137
rect 39396 23128 39448 23180
rect 40868 23171 40920 23180
rect 16120 23060 16172 23112
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18236 23060 18288 23112
rect 22468 23103 22520 23112
rect 22468 23069 22477 23103
rect 22477 23069 22511 23103
rect 22511 23069 22520 23103
rect 22468 23060 22520 23069
rect 22744 23103 22796 23112
rect 22744 23069 22753 23103
rect 22753 23069 22787 23103
rect 22787 23069 22796 23103
rect 22744 23060 22796 23069
rect 24400 23060 24452 23112
rect 24492 23060 24544 23112
rect 27344 23060 27396 23112
rect 28540 23060 28592 23112
rect 30012 23103 30064 23112
rect 30012 23069 30021 23103
rect 30021 23069 30055 23103
rect 30055 23069 30064 23103
rect 30012 23060 30064 23069
rect 32220 23103 32272 23112
rect 32220 23069 32229 23103
rect 32229 23069 32263 23103
rect 32263 23069 32272 23103
rect 32220 23060 32272 23069
rect 33324 23060 33376 23112
rect 37924 23060 37976 23112
rect 38936 23103 38988 23112
rect 38936 23069 38945 23103
rect 38945 23069 38979 23103
rect 38979 23069 38988 23103
rect 40868 23137 40877 23171
rect 40877 23137 40911 23171
rect 40911 23137 40920 23171
rect 40868 23128 40920 23137
rect 40960 23128 41012 23180
rect 43628 23128 43680 23180
rect 43996 23128 44048 23180
rect 44640 23171 44692 23180
rect 44640 23137 44658 23171
rect 44658 23137 44692 23171
rect 44640 23128 44692 23137
rect 45008 23128 45060 23180
rect 38936 23060 38988 23069
rect 21916 22992 21968 23044
rect 15660 22924 15712 22976
rect 16672 22967 16724 22976
rect 16672 22933 16681 22967
rect 16681 22933 16715 22967
rect 16715 22933 16724 22967
rect 16672 22924 16724 22933
rect 20168 22967 20220 22976
rect 20168 22933 20177 22967
rect 20177 22933 20211 22967
rect 20211 22933 20220 22967
rect 20168 22924 20220 22933
rect 24768 22992 24820 23044
rect 25412 22992 25464 23044
rect 38200 22992 38252 23044
rect 40224 22992 40276 23044
rect 43168 22992 43220 23044
rect 43904 22992 43956 23044
rect 23848 22967 23900 22976
rect 23848 22933 23857 22967
rect 23857 22933 23891 22967
rect 23891 22933 23900 22967
rect 23848 22924 23900 22933
rect 25504 22924 25556 22976
rect 27712 22967 27764 22976
rect 27712 22933 27721 22967
rect 27721 22933 27755 22967
rect 27755 22933 27764 22967
rect 27712 22924 27764 22933
rect 28264 22924 28316 22976
rect 29184 22924 29236 22976
rect 29368 22967 29420 22976
rect 29368 22933 29377 22967
rect 29377 22933 29411 22967
rect 29411 22933 29420 22967
rect 29368 22924 29420 22933
rect 35256 22924 35308 22976
rect 37188 22924 37240 22976
rect 42616 22924 42668 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 15844 22720 15896 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 22192 22720 22244 22772
rect 23296 22720 23348 22772
rect 25044 22720 25096 22772
rect 26424 22763 26476 22772
rect 26424 22729 26433 22763
rect 26433 22729 26467 22763
rect 26467 22729 26476 22763
rect 26424 22720 26476 22729
rect 29368 22720 29420 22772
rect 31852 22763 31904 22772
rect 31852 22729 31861 22763
rect 31861 22729 31895 22763
rect 31895 22729 31904 22763
rect 31852 22720 31904 22729
rect 32220 22763 32272 22772
rect 32220 22729 32229 22763
rect 32229 22729 32263 22763
rect 32263 22729 32272 22763
rect 32220 22720 32272 22729
rect 33876 22763 33928 22772
rect 33876 22729 33885 22763
rect 33885 22729 33919 22763
rect 33919 22729 33928 22763
rect 33876 22720 33928 22729
rect 36636 22763 36688 22772
rect 20628 22695 20680 22704
rect 20628 22661 20637 22695
rect 20637 22661 20671 22695
rect 20671 22661 20680 22695
rect 20628 22652 20680 22661
rect 21364 22652 21416 22704
rect 23756 22652 23808 22704
rect 24400 22652 24452 22704
rect 16120 22584 16172 22636
rect 19156 22584 19208 22636
rect 22376 22627 22428 22636
rect 22376 22593 22385 22627
rect 22385 22593 22419 22627
rect 22419 22593 22428 22627
rect 22376 22584 22428 22593
rect 22928 22584 22980 22636
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25780 22652 25832 22704
rect 30380 22652 30432 22704
rect 26332 22584 26384 22636
rect 26976 22627 27028 22636
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 27160 22584 27212 22636
rect 29184 22584 29236 22636
rect 32496 22627 32548 22636
rect 14648 22516 14700 22568
rect 32496 22593 32505 22627
rect 32505 22593 32539 22627
rect 32539 22593 32548 22627
rect 32496 22584 32548 22593
rect 32680 22584 32732 22636
rect 35256 22652 35308 22704
rect 35348 22652 35400 22704
rect 36636 22729 36645 22763
rect 36645 22729 36679 22763
rect 36679 22729 36688 22763
rect 36636 22720 36688 22729
rect 38200 22720 38252 22772
rect 38936 22763 38988 22772
rect 38936 22729 38945 22763
rect 38945 22729 38979 22763
rect 38979 22729 38988 22763
rect 38936 22720 38988 22729
rect 37740 22652 37792 22704
rect 37188 22627 37240 22636
rect 37188 22593 37197 22627
rect 37197 22593 37231 22627
rect 37231 22593 37240 22627
rect 37188 22584 37240 22593
rect 37280 22584 37332 22636
rect 15660 22448 15712 22500
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 15936 22491 15988 22500
rect 15936 22457 15945 22491
rect 15945 22457 15979 22491
rect 15979 22457 15988 22491
rect 15936 22448 15988 22457
rect 17960 22448 18012 22500
rect 18328 22448 18380 22500
rect 19616 22448 19668 22500
rect 20076 22491 20128 22500
rect 20076 22457 20085 22491
rect 20085 22457 20119 22491
rect 20119 22457 20128 22491
rect 20076 22448 20128 22457
rect 20168 22491 20220 22500
rect 20168 22457 20177 22491
rect 20177 22457 20211 22491
rect 20211 22457 20220 22491
rect 22100 22491 22152 22500
rect 20168 22448 20220 22457
rect 22100 22457 22109 22491
rect 22109 22457 22143 22491
rect 22143 22457 22152 22491
rect 22100 22448 22152 22457
rect 22192 22491 22244 22500
rect 22192 22457 22201 22491
rect 22201 22457 22235 22491
rect 22235 22457 22244 22491
rect 22192 22448 22244 22457
rect 23480 22491 23532 22500
rect 23480 22457 23489 22491
rect 23489 22457 23523 22491
rect 23523 22457 23532 22491
rect 23480 22448 23532 22457
rect 24308 22448 24360 22500
rect 24492 22491 24544 22500
rect 24492 22457 24501 22491
rect 24501 22457 24535 22491
rect 24535 22457 24544 22491
rect 24492 22448 24544 22457
rect 25412 22491 25464 22500
rect 25412 22457 25421 22491
rect 25421 22457 25455 22491
rect 25455 22457 25464 22491
rect 25412 22448 25464 22457
rect 25596 22448 25648 22500
rect 20352 22380 20404 22432
rect 29644 22448 29696 22500
rect 30748 22448 30800 22500
rect 40040 22720 40092 22772
rect 43996 22763 44048 22772
rect 43996 22729 44005 22763
rect 44005 22729 44039 22763
rect 44039 22729 44048 22763
rect 43996 22720 44048 22729
rect 42708 22652 42760 22704
rect 43168 22652 43220 22704
rect 43076 22627 43128 22636
rect 43076 22593 43085 22627
rect 43085 22593 43119 22627
rect 43119 22593 43128 22627
rect 43076 22584 43128 22593
rect 40224 22516 40276 22568
rect 44456 22516 44508 22568
rect 45836 22516 45888 22568
rect 34796 22448 34848 22500
rect 35808 22448 35860 22500
rect 37832 22448 37884 22500
rect 28540 22423 28592 22432
rect 28540 22389 28549 22423
rect 28549 22389 28583 22423
rect 28583 22389 28592 22423
rect 28540 22380 28592 22389
rect 33048 22380 33100 22432
rect 34152 22423 34204 22432
rect 34152 22389 34161 22423
rect 34161 22389 34195 22423
rect 34195 22389 34204 22423
rect 34152 22380 34204 22389
rect 35992 22423 36044 22432
rect 35992 22389 36001 22423
rect 36001 22389 36035 22423
rect 36035 22389 36044 22423
rect 35992 22380 36044 22389
rect 37556 22380 37608 22432
rect 39672 22448 39724 22500
rect 40868 22491 40920 22500
rect 40868 22457 40877 22491
rect 40877 22457 40911 22491
rect 40911 22457 40920 22491
rect 40868 22448 40920 22457
rect 43168 22491 43220 22500
rect 43168 22457 43177 22491
rect 43177 22457 43211 22491
rect 43211 22457 43220 22491
rect 43168 22448 43220 22457
rect 45192 22448 45244 22500
rect 39304 22423 39356 22432
rect 39304 22389 39313 22423
rect 39313 22389 39347 22423
rect 39347 22389 39356 22423
rect 39304 22380 39356 22389
rect 40776 22380 40828 22432
rect 41604 22380 41656 22432
rect 43444 22380 43496 22432
rect 45008 22423 45060 22432
rect 45008 22389 45017 22423
rect 45017 22389 45051 22423
rect 45051 22389 45060 22423
rect 45008 22380 45060 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 15844 22219 15896 22228
rect 15844 22185 15853 22219
rect 15853 22185 15887 22219
rect 15887 22185 15896 22219
rect 15844 22176 15896 22185
rect 16120 22219 16172 22228
rect 16120 22185 16129 22219
rect 16129 22185 16163 22219
rect 16163 22185 16172 22219
rect 16120 22176 16172 22185
rect 18144 22176 18196 22228
rect 20168 22176 20220 22228
rect 22100 22219 22152 22228
rect 22100 22185 22109 22219
rect 22109 22185 22143 22219
rect 22143 22185 22152 22219
rect 22100 22176 22152 22185
rect 22468 22219 22520 22228
rect 22468 22185 22477 22219
rect 22477 22185 22511 22219
rect 22511 22185 22520 22219
rect 22468 22176 22520 22185
rect 23296 22176 23348 22228
rect 23940 22176 23992 22228
rect 25504 22176 25556 22228
rect 26976 22219 27028 22228
rect 26976 22185 26985 22219
rect 26985 22185 27019 22219
rect 27019 22185 27028 22219
rect 26976 22176 27028 22185
rect 27344 22219 27396 22228
rect 27344 22185 27353 22219
rect 27353 22185 27387 22219
rect 27387 22185 27396 22219
rect 27344 22176 27396 22185
rect 32496 22219 32548 22228
rect 32496 22185 32505 22219
rect 32505 22185 32539 22219
rect 32539 22185 32548 22219
rect 32496 22176 32548 22185
rect 33048 22219 33100 22228
rect 33048 22185 33057 22219
rect 33057 22185 33091 22219
rect 33091 22185 33100 22219
rect 33048 22176 33100 22185
rect 34796 22219 34848 22228
rect 34796 22185 34805 22219
rect 34805 22185 34839 22219
rect 34839 22185 34848 22219
rect 34796 22176 34848 22185
rect 35256 22176 35308 22228
rect 37188 22219 37240 22228
rect 37188 22185 37197 22219
rect 37197 22185 37231 22219
rect 37231 22185 37240 22219
rect 37188 22176 37240 22185
rect 37648 22176 37700 22228
rect 40960 22219 41012 22228
rect 16672 22108 16724 22160
rect 19432 22151 19484 22160
rect 19432 22117 19441 22151
rect 19441 22117 19475 22151
rect 19475 22117 19484 22151
rect 19432 22108 19484 22117
rect 19984 22151 20036 22160
rect 19984 22117 19993 22151
rect 19993 22117 20027 22151
rect 20027 22117 20036 22151
rect 19984 22108 20036 22117
rect 23020 22108 23072 22160
rect 24308 22151 24360 22160
rect 24308 22117 24317 22151
rect 24317 22117 24351 22151
rect 24351 22117 24360 22151
rect 24308 22108 24360 22117
rect 25412 22108 25464 22160
rect 28632 22108 28684 22160
rect 30564 22151 30616 22160
rect 30564 22117 30573 22151
rect 30573 22117 30607 22151
rect 30607 22117 30616 22151
rect 30564 22108 30616 22117
rect 34520 22108 34572 22160
rect 35808 22151 35860 22160
rect 35808 22117 35817 22151
rect 35817 22117 35851 22151
rect 35851 22117 35860 22151
rect 35808 22108 35860 22117
rect 36360 22151 36412 22160
rect 36360 22117 36369 22151
rect 36369 22117 36403 22151
rect 36403 22117 36412 22151
rect 36360 22108 36412 22117
rect 37832 22108 37884 22160
rect 40960 22185 40969 22219
rect 40969 22185 41003 22219
rect 41003 22185 41012 22219
rect 40960 22176 41012 22185
rect 43076 22219 43128 22228
rect 43076 22185 43085 22219
rect 43085 22185 43119 22219
rect 43119 22185 43128 22219
rect 43076 22176 43128 22185
rect 43352 22176 43404 22228
rect 45652 22176 45704 22228
rect 41420 22151 41472 22160
rect 41420 22117 41429 22151
rect 41429 22117 41463 22151
rect 41463 22117 41472 22151
rect 41420 22108 41472 22117
rect 43444 22151 43496 22160
rect 43444 22117 43453 22151
rect 43453 22117 43487 22151
rect 43487 22117 43496 22151
rect 43444 22108 43496 22117
rect 43536 22151 43588 22160
rect 43536 22117 43545 22151
rect 43545 22117 43579 22151
rect 43579 22117 43588 22151
rect 45376 22151 45428 22160
rect 43536 22108 43588 22117
rect 45376 22117 45385 22151
rect 45385 22117 45419 22151
rect 45419 22117 45428 22151
rect 45376 22108 45428 22117
rect 15200 22040 15252 22092
rect 17224 22040 17276 22092
rect 18144 22040 18196 22092
rect 20352 22040 20404 22092
rect 22008 22040 22060 22092
rect 26608 22083 26660 22092
rect 26608 22049 26626 22083
rect 26626 22049 26660 22083
rect 26608 22040 26660 22049
rect 27252 22040 27304 22092
rect 27436 22040 27488 22092
rect 29552 22040 29604 22092
rect 32680 22040 32732 22092
rect 39212 22040 39264 22092
rect 39856 22040 39908 22092
rect 46480 22040 46532 22092
rect 46756 22083 46808 22092
rect 46756 22049 46765 22083
rect 46765 22049 46799 22083
rect 46799 22049 46808 22083
rect 46756 22040 46808 22049
rect 19340 22015 19392 22024
rect 19340 21981 19349 22015
rect 19349 21981 19383 22015
rect 19383 21981 19392 22015
rect 19340 21972 19392 21981
rect 22744 21972 22796 22024
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 24216 22015 24268 22024
rect 24216 21981 24225 22015
rect 24225 21981 24259 22015
rect 24259 21981 24268 22015
rect 24216 21972 24268 21981
rect 24400 21972 24452 22024
rect 25596 21972 25648 22024
rect 28356 21972 28408 22024
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 32128 22015 32180 22024
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 33876 22015 33928 22024
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 35716 22015 35768 22024
rect 35716 21981 35725 22015
rect 35725 21981 35759 22015
rect 35759 21981 35768 22015
rect 35716 21972 35768 21981
rect 20076 21904 20128 21956
rect 21640 21836 21692 21888
rect 27988 21904 28040 21956
rect 25320 21836 25372 21888
rect 30012 21836 30064 21888
rect 31668 21836 31720 21888
rect 36728 21879 36780 21888
rect 36728 21845 36737 21879
rect 36737 21845 36771 21879
rect 36771 21845 36780 21879
rect 36728 21836 36780 21845
rect 37464 21879 37516 21888
rect 37464 21845 37473 21879
rect 37473 21845 37507 21879
rect 37507 21845 37516 21879
rect 41052 21972 41104 22024
rect 41512 21972 41564 22024
rect 45284 22015 45336 22024
rect 45284 21981 45293 22015
rect 45293 21981 45327 22015
rect 45327 21981 45336 22015
rect 45284 21972 45336 21981
rect 42984 21904 43036 21956
rect 45468 21972 45520 22024
rect 44548 21879 44600 21888
rect 37464 21836 37516 21845
rect 44548 21845 44557 21879
rect 44557 21845 44591 21879
rect 44591 21845 44600 21879
rect 44548 21836 44600 21845
rect 45744 21836 45796 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 17960 21632 18012 21684
rect 19340 21632 19392 21684
rect 19064 21564 19116 21616
rect 16488 21539 16540 21548
rect 16488 21505 16497 21539
rect 16497 21505 16531 21539
rect 16531 21505 16540 21539
rect 16488 21496 16540 21505
rect 19432 21496 19484 21548
rect 20260 21632 20312 21684
rect 22468 21632 22520 21684
rect 23020 21675 23072 21684
rect 23020 21641 23029 21675
rect 23029 21641 23063 21675
rect 23063 21641 23072 21675
rect 23020 21632 23072 21641
rect 24308 21632 24360 21684
rect 25596 21632 25648 21684
rect 26608 21675 26660 21684
rect 26608 21641 26617 21675
rect 26617 21641 26651 21675
rect 26651 21641 26660 21675
rect 26608 21632 26660 21641
rect 27436 21675 27488 21684
rect 27436 21641 27445 21675
rect 27445 21641 27479 21675
rect 27479 21641 27488 21675
rect 27436 21632 27488 21641
rect 28632 21675 28684 21684
rect 28632 21641 28641 21675
rect 28641 21641 28675 21675
rect 28675 21641 28684 21675
rect 28632 21632 28684 21641
rect 30564 21675 30616 21684
rect 20536 21428 20588 21480
rect 21548 21428 21600 21480
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 25504 21496 25556 21548
rect 27620 21471 27672 21480
rect 22744 21360 22796 21412
rect 23572 21360 23624 21412
rect 23940 21403 23992 21412
rect 23940 21369 23949 21403
rect 23949 21369 23983 21403
rect 23983 21369 23992 21403
rect 23940 21360 23992 21369
rect 25596 21360 25648 21412
rect 13820 21292 13872 21344
rect 15200 21292 15252 21344
rect 17224 21292 17276 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18144 21292 18196 21344
rect 20536 21292 20588 21344
rect 21640 21292 21692 21344
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 23664 21292 23716 21344
rect 23756 21292 23808 21344
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 27712 21360 27764 21412
rect 28356 21403 28408 21412
rect 28356 21369 28365 21403
rect 28365 21369 28399 21403
rect 28399 21369 28408 21403
rect 28356 21360 28408 21369
rect 30564 21641 30573 21675
rect 30573 21641 30607 21675
rect 30607 21641 30616 21675
rect 30564 21632 30616 21641
rect 30748 21632 30800 21684
rect 32496 21632 32548 21684
rect 34520 21632 34572 21684
rect 35716 21675 35768 21684
rect 35716 21641 35725 21675
rect 35725 21641 35759 21675
rect 35759 21641 35768 21675
rect 35716 21632 35768 21641
rect 35808 21632 35860 21684
rect 37832 21632 37884 21684
rect 38108 21632 38160 21684
rect 39856 21675 39908 21684
rect 30472 21564 30524 21616
rect 31208 21564 31260 21616
rect 32772 21564 32824 21616
rect 31668 21539 31720 21548
rect 31668 21505 31677 21539
rect 31677 21505 31711 21539
rect 31711 21505 31720 21539
rect 31668 21496 31720 21505
rect 29276 21471 29328 21480
rect 29276 21437 29285 21471
rect 29285 21437 29319 21471
rect 29319 21437 29328 21471
rect 29276 21428 29328 21437
rect 33876 21496 33928 21548
rect 30748 21360 30800 21412
rect 31760 21403 31812 21412
rect 31760 21369 31769 21403
rect 31769 21369 31803 21403
rect 31803 21369 31812 21403
rect 32312 21403 32364 21412
rect 31760 21360 31812 21369
rect 32312 21369 32321 21403
rect 32321 21369 32355 21403
rect 32355 21369 32364 21403
rect 32312 21360 32364 21369
rect 32680 21360 32732 21412
rect 33324 21428 33376 21480
rect 34152 21428 34204 21480
rect 37556 21496 37608 21548
rect 36728 21428 36780 21480
rect 39856 21641 39865 21675
rect 39865 21641 39899 21675
rect 39899 21641 39908 21675
rect 39856 21632 39908 21641
rect 41420 21675 41472 21684
rect 41420 21641 41429 21675
rect 41429 21641 41463 21675
rect 41463 21641 41472 21675
rect 41420 21632 41472 21641
rect 42708 21632 42760 21684
rect 43444 21632 43496 21684
rect 45284 21632 45336 21684
rect 42892 21564 42944 21616
rect 40776 21496 40828 21548
rect 42340 21539 42392 21548
rect 42340 21505 42349 21539
rect 42349 21505 42383 21539
rect 42383 21505 42392 21539
rect 42340 21496 42392 21505
rect 42984 21539 43036 21548
rect 42984 21505 42993 21539
rect 42993 21505 43027 21539
rect 43027 21505 43036 21539
rect 42984 21496 43036 21505
rect 45652 21564 45704 21616
rect 46756 21564 46808 21616
rect 43536 21496 43588 21548
rect 44548 21539 44600 21548
rect 44548 21505 44557 21539
rect 44557 21505 44591 21539
rect 44591 21505 44600 21539
rect 44548 21496 44600 21505
rect 40500 21471 40552 21480
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 34520 21292 34572 21344
rect 38016 21360 38068 21412
rect 40500 21437 40509 21471
rect 40509 21437 40543 21471
rect 40543 21437 40552 21471
rect 40500 21428 40552 21437
rect 37556 21335 37608 21344
rect 37556 21301 37565 21335
rect 37565 21301 37599 21335
rect 37599 21301 37608 21335
rect 37556 21292 37608 21301
rect 38384 21292 38436 21344
rect 39764 21360 39816 21412
rect 44640 21403 44692 21412
rect 40316 21335 40368 21344
rect 40316 21301 40325 21335
rect 40325 21301 40359 21335
rect 40359 21301 40368 21335
rect 40316 21292 40368 21301
rect 41420 21292 41472 21344
rect 44640 21369 44649 21403
rect 44649 21369 44683 21403
rect 44683 21369 44692 21403
rect 44640 21360 44692 21369
rect 45192 21403 45244 21412
rect 45192 21369 45201 21403
rect 45201 21369 45235 21403
rect 45235 21369 45244 21403
rect 45192 21360 45244 21369
rect 46940 21428 46992 21480
rect 47584 21471 47636 21480
rect 47584 21437 47593 21471
rect 47593 21437 47627 21471
rect 47627 21437 47636 21471
rect 47584 21428 47636 21437
rect 45376 21292 45428 21344
rect 46664 21335 46716 21344
rect 46664 21301 46673 21335
rect 46673 21301 46707 21335
rect 46707 21301 46716 21335
rect 46664 21292 46716 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 15292 21088 15344 21140
rect 17224 21088 17276 21140
rect 19248 21088 19300 21140
rect 22744 21131 22796 21140
rect 18972 21020 19024 21072
rect 18880 20952 18932 21004
rect 22744 21097 22753 21131
rect 22753 21097 22787 21131
rect 22787 21097 22796 21131
rect 22744 21088 22796 21097
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 24216 21131 24268 21140
rect 24216 21097 24225 21131
rect 24225 21097 24259 21131
rect 24259 21097 24268 21131
rect 24216 21088 24268 21097
rect 27620 21131 27672 21140
rect 27620 21097 27629 21131
rect 27629 21097 27663 21131
rect 27663 21097 27672 21131
rect 27620 21088 27672 21097
rect 28356 21088 28408 21140
rect 32128 21088 32180 21140
rect 32588 21088 32640 21140
rect 29276 21063 29328 21072
rect 29276 21029 29285 21063
rect 29285 21029 29319 21063
rect 29319 21029 29328 21063
rect 29276 21020 29328 21029
rect 30196 21020 30248 21072
rect 32312 21020 32364 21072
rect 22652 20952 22704 21004
rect 25872 20952 25924 21004
rect 27068 20952 27120 21004
rect 28080 20995 28132 21004
rect 28080 20961 28089 20995
rect 28089 20961 28123 20995
rect 28123 20961 28132 20995
rect 28080 20952 28132 20961
rect 28172 20952 28224 21004
rect 17500 20884 17552 20936
rect 18052 20927 18104 20936
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 18696 20927 18748 20936
rect 18696 20893 18705 20927
rect 18705 20893 18739 20927
rect 18739 20893 18748 20927
rect 18696 20884 18748 20893
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 16948 20816 17000 20868
rect 27712 20816 27764 20868
rect 32680 20995 32732 21004
rect 32680 20961 32689 20995
rect 32689 20961 32723 20995
rect 32723 20961 32732 20995
rect 32680 20952 32732 20961
rect 37832 21088 37884 21140
rect 40500 21131 40552 21140
rect 40500 21097 40509 21131
rect 40509 21097 40543 21131
rect 40543 21097 40552 21131
rect 40500 21088 40552 21097
rect 41052 21131 41104 21140
rect 41052 21097 41061 21131
rect 41061 21097 41095 21131
rect 41095 21097 41104 21131
rect 41052 21088 41104 21097
rect 42340 21131 42392 21140
rect 42340 21097 42349 21131
rect 42349 21097 42383 21131
rect 42383 21097 42392 21131
rect 42340 21088 42392 21097
rect 44640 21088 44692 21140
rect 35900 21020 35952 21072
rect 37556 21020 37608 21072
rect 41420 21063 41472 21072
rect 41420 21029 41429 21063
rect 41429 21029 41463 21063
rect 41463 21029 41472 21063
rect 41420 21020 41472 21029
rect 43996 21020 44048 21072
rect 45376 21020 45428 21072
rect 45560 21020 45612 21072
rect 45744 21063 45796 21072
rect 45744 21029 45753 21063
rect 45753 21029 45787 21063
rect 45787 21029 45796 21063
rect 45744 21020 45796 21029
rect 45836 21063 45888 21072
rect 45836 21029 45845 21063
rect 45845 21029 45879 21063
rect 45879 21029 45888 21063
rect 45836 21020 45888 21029
rect 34152 20995 34204 21004
rect 34152 20961 34161 20995
rect 34161 20961 34195 20995
rect 34195 20961 34204 20995
rect 34152 20952 34204 20961
rect 35256 20952 35308 21004
rect 39028 20952 39080 21004
rect 39764 20995 39816 21004
rect 39764 20961 39773 20995
rect 39773 20961 39807 20995
rect 39807 20961 39816 20995
rect 39764 20952 39816 20961
rect 29828 20884 29880 20936
rect 34796 20927 34848 20936
rect 34796 20893 34805 20927
rect 34805 20893 34839 20927
rect 34839 20893 34848 20927
rect 34796 20884 34848 20893
rect 36360 20884 36412 20936
rect 37280 20884 37332 20936
rect 38108 20884 38160 20936
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 41328 20927 41380 20936
rect 30932 20816 30984 20868
rect 41328 20893 41337 20927
rect 41337 20893 41371 20927
rect 41371 20893 41380 20927
rect 41328 20884 41380 20893
rect 44364 20884 44416 20936
rect 45560 20884 45612 20936
rect 41512 20816 41564 20868
rect 18788 20748 18840 20800
rect 26516 20748 26568 20800
rect 31024 20791 31076 20800
rect 31024 20757 31033 20791
rect 31033 20757 31067 20791
rect 31067 20757 31076 20791
rect 31024 20748 31076 20757
rect 33324 20791 33376 20800
rect 33324 20757 33333 20791
rect 33333 20757 33367 20791
rect 33367 20757 33376 20791
rect 33324 20748 33376 20757
rect 38936 20791 38988 20800
rect 38936 20757 38945 20791
rect 38945 20757 38979 20791
rect 38979 20757 38988 20791
rect 38936 20748 38988 20757
rect 44732 20748 44784 20800
rect 46848 20748 46900 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 17132 20544 17184 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 17776 20587 17828 20596
rect 17776 20553 17785 20587
rect 17785 20553 17819 20587
rect 17819 20553 17828 20587
rect 17776 20544 17828 20553
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 21272 20544 21324 20596
rect 22652 20587 22704 20596
rect 16948 20476 17000 20528
rect 18696 20476 18748 20528
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 25872 20587 25924 20596
rect 25872 20553 25881 20587
rect 25881 20553 25915 20587
rect 25915 20553 25924 20587
rect 25872 20544 25924 20553
rect 28172 20544 28224 20596
rect 30196 20544 30248 20596
rect 30748 20544 30800 20596
rect 31760 20544 31812 20596
rect 32588 20544 32640 20596
rect 32680 20587 32732 20596
rect 32680 20553 32689 20587
rect 32689 20553 32723 20587
rect 32723 20553 32732 20587
rect 32956 20587 33008 20596
rect 32680 20544 32732 20553
rect 32956 20553 32965 20587
rect 32965 20553 32999 20587
rect 32999 20553 33008 20587
rect 32956 20544 33008 20553
rect 34520 20544 34572 20596
rect 37556 20544 37608 20596
rect 38108 20587 38160 20596
rect 38108 20553 38117 20587
rect 38117 20553 38151 20587
rect 38151 20553 38160 20587
rect 38108 20544 38160 20553
rect 38844 20544 38896 20596
rect 39028 20544 39080 20596
rect 42892 20587 42944 20596
rect 42892 20553 42901 20587
rect 42901 20553 42935 20587
rect 42935 20553 42944 20587
rect 42892 20544 42944 20553
rect 44364 20587 44416 20596
rect 44364 20553 44373 20587
rect 44373 20553 44407 20587
rect 44407 20553 44416 20587
rect 44364 20544 44416 20553
rect 45744 20544 45796 20596
rect 45836 20587 45888 20596
rect 45836 20553 45845 20587
rect 45845 20553 45879 20587
rect 45879 20553 45888 20587
rect 45836 20544 45888 20553
rect 28080 20476 28132 20528
rect 33048 20476 33100 20528
rect 33324 20476 33376 20528
rect 43996 20519 44048 20528
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 17776 20272 17828 20324
rect 18236 20204 18288 20256
rect 20076 20340 20128 20392
rect 20904 20272 20956 20324
rect 26884 20408 26936 20460
rect 25136 20383 25188 20392
rect 25136 20349 25154 20383
rect 25154 20349 25188 20383
rect 25136 20340 25188 20349
rect 26516 20383 26568 20392
rect 26516 20349 26525 20383
rect 26525 20349 26559 20383
rect 26559 20349 26568 20383
rect 26516 20340 26568 20349
rect 27712 20383 27764 20392
rect 27712 20349 27721 20383
rect 27721 20349 27755 20383
rect 27755 20349 27764 20383
rect 27712 20340 27764 20349
rect 30104 20408 30156 20460
rect 31024 20451 31076 20460
rect 31024 20417 31033 20451
rect 31033 20417 31067 20451
rect 31067 20417 31076 20451
rect 31024 20408 31076 20417
rect 33140 20408 33192 20460
rect 34796 20408 34848 20460
rect 35256 20408 35308 20460
rect 21824 20272 21876 20324
rect 21548 20204 21600 20256
rect 23480 20272 23532 20324
rect 26056 20315 26108 20324
rect 26056 20281 26065 20315
rect 26065 20281 26099 20315
rect 26099 20281 26108 20315
rect 26056 20272 26108 20281
rect 27252 20272 27304 20324
rect 29000 20272 29052 20324
rect 33232 20383 33284 20392
rect 33232 20349 33241 20383
rect 33241 20349 33275 20383
rect 33275 20349 33284 20383
rect 33232 20340 33284 20349
rect 33416 20340 33468 20392
rect 36636 20383 36688 20392
rect 36636 20349 36645 20383
rect 36645 20349 36679 20383
rect 36679 20349 36688 20383
rect 36636 20340 36688 20349
rect 36820 20340 36872 20392
rect 38844 20383 38896 20392
rect 38844 20349 38853 20383
rect 38853 20349 38887 20383
rect 38887 20349 38896 20383
rect 38844 20340 38896 20349
rect 38936 20340 38988 20392
rect 40500 20383 40552 20392
rect 40500 20349 40509 20383
rect 40509 20349 40543 20383
rect 40543 20349 40552 20383
rect 40500 20340 40552 20349
rect 30196 20272 30248 20324
rect 30748 20272 30800 20324
rect 34520 20272 34572 20324
rect 22376 20204 22428 20256
rect 25044 20204 25096 20256
rect 30104 20247 30156 20256
rect 30104 20213 30113 20247
rect 30113 20213 30147 20247
rect 30147 20213 30156 20247
rect 30104 20204 30156 20213
rect 34152 20247 34204 20256
rect 34152 20213 34161 20247
rect 34161 20213 34195 20247
rect 34195 20213 34204 20247
rect 34152 20204 34204 20213
rect 35808 20247 35860 20256
rect 35808 20213 35817 20247
rect 35817 20213 35851 20247
rect 35851 20213 35860 20247
rect 35808 20204 35860 20213
rect 36728 20247 36780 20256
rect 36728 20213 36737 20247
rect 36737 20213 36771 20247
rect 36771 20213 36780 20247
rect 36728 20204 36780 20213
rect 38016 20204 38068 20256
rect 40316 20272 40368 20324
rect 43996 20485 44005 20519
rect 44005 20485 44039 20519
rect 44039 20485 44048 20519
rect 43996 20476 44048 20485
rect 45376 20476 45428 20528
rect 47032 20476 47084 20528
rect 43168 20408 43220 20460
rect 41328 20272 41380 20324
rect 43076 20315 43128 20324
rect 43076 20281 43085 20315
rect 43085 20281 43119 20315
rect 43119 20281 43128 20315
rect 43076 20272 43128 20281
rect 46204 20315 46256 20324
rect 41420 20247 41472 20256
rect 41420 20213 41429 20247
rect 41429 20213 41463 20247
rect 41463 20213 41472 20247
rect 41420 20204 41472 20213
rect 41880 20204 41932 20256
rect 42892 20204 42944 20256
rect 46204 20281 46213 20315
rect 46213 20281 46247 20315
rect 46247 20281 46256 20315
rect 46204 20272 46256 20281
rect 46848 20315 46900 20324
rect 45744 20204 45796 20256
rect 46848 20281 46857 20315
rect 46857 20281 46891 20315
rect 46891 20281 46900 20315
rect 46848 20272 46900 20281
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 18052 20043 18104 20052
rect 18052 20009 18061 20043
rect 18061 20009 18095 20043
rect 18095 20009 18104 20043
rect 18052 20000 18104 20009
rect 16856 19864 16908 19916
rect 17500 19864 17552 19916
rect 18236 19864 18288 19916
rect 18512 19864 18564 19916
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 21824 20043 21876 20052
rect 21824 20009 21833 20043
rect 21833 20009 21867 20043
rect 21867 20009 21876 20043
rect 21824 20000 21876 20009
rect 26516 20000 26568 20052
rect 27712 20043 27764 20052
rect 27712 20009 27721 20043
rect 27721 20009 27755 20043
rect 27755 20009 27764 20043
rect 27712 20000 27764 20009
rect 29828 20043 29880 20052
rect 29828 20009 29837 20043
rect 29837 20009 29871 20043
rect 29871 20009 29880 20043
rect 29828 20000 29880 20009
rect 32404 20000 32456 20052
rect 33784 20000 33836 20052
rect 34520 20000 34572 20052
rect 35808 20000 35860 20052
rect 36360 20000 36412 20052
rect 37464 20000 37516 20052
rect 38936 20000 38988 20052
rect 40500 20043 40552 20052
rect 40500 20009 40509 20043
rect 40509 20009 40543 20043
rect 40543 20009 40552 20043
rect 40500 20000 40552 20009
rect 43076 20043 43128 20052
rect 43076 20009 43085 20043
rect 43085 20009 43119 20043
rect 43119 20009 43128 20043
rect 43076 20000 43128 20009
rect 45744 20043 45796 20052
rect 45744 20009 45753 20043
rect 45753 20009 45787 20043
rect 45787 20009 45796 20043
rect 45744 20000 45796 20009
rect 46204 20000 46256 20052
rect 23296 19975 23348 19984
rect 23296 19941 23305 19975
rect 23305 19941 23339 19975
rect 23339 19941 23348 19975
rect 23296 19932 23348 19941
rect 27252 19932 27304 19984
rect 29000 19975 29052 19984
rect 29000 19941 29009 19975
rect 29009 19941 29043 19975
rect 29043 19941 29052 19975
rect 29000 19932 29052 19941
rect 32680 19932 32732 19984
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 22376 19864 22428 19916
rect 24952 19907 25004 19916
rect 24952 19873 24961 19907
rect 24961 19873 24995 19907
rect 24995 19873 25004 19907
rect 24952 19864 25004 19873
rect 29276 19864 29328 19916
rect 30840 19864 30892 19916
rect 30932 19907 30984 19916
rect 30932 19873 30941 19907
rect 30941 19873 30975 19907
rect 30975 19873 30984 19907
rect 30932 19864 30984 19873
rect 31944 19864 31996 19916
rect 33876 19932 33928 19984
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 26884 19839 26936 19848
rect 25688 19728 25740 19780
rect 26884 19805 26893 19839
rect 26893 19805 26927 19839
rect 26927 19805 26936 19839
rect 26884 19796 26936 19805
rect 31024 19839 31076 19848
rect 31024 19805 31033 19839
rect 31033 19805 31067 19839
rect 31067 19805 31076 19839
rect 31024 19796 31076 19805
rect 32956 19796 33008 19848
rect 35624 19907 35676 19916
rect 35624 19873 35633 19907
rect 35633 19873 35667 19907
rect 35667 19873 35676 19907
rect 35624 19864 35676 19873
rect 36176 19864 36228 19916
rect 39304 19907 39356 19916
rect 27620 19728 27672 19780
rect 27712 19728 27764 19780
rect 31116 19728 31168 19780
rect 39304 19873 39313 19907
rect 39313 19873 39347 19907
rect 39347 19873 39356 19907
rect 39304 19864 39356 19873
rect 41604 19932 41656 19984
rect 41880 19975 41932 19984
rect 41880 19941 41889 19975
rect 41889 19941 41923 19975
rect 41923 19941 41932 19975
rect 41880 19932 41932 19941
rect 40040 19839 40092 19848
rect 40040 19805 40049 19839
rect 40049 19805 40083 19839
rect 40083 19805 40092 19839
rect 40040 19796 40092 19805
rect 43720 19932 43772 19984
rect 44824 19864 44876 19916
rect 45836 19907 45888 19916
rect 45836 19873 45845 19907
rect 45845 19873 45879 19907
rect 45879 19873 45888 19907
rect 45836 19864 45888 19873
rect 43444 19839 43496 19848
rect 43444 19805 43453 19839
rect 43453 19805 43487 19839
rect 43487 19805 43496 19839
rect 43444 19796 43496 19805
rect 43628 19796 43680 19848
rect 38384 19728 38436 19780
rect 45284 19728 45336 19780
rect 20076 19703 20128 19712
rect 20076 19669 20085 19703
rect 20085 19669 20119 19703
rect 20119 19669 20128 19703
rect 20076 19660 20128 19669
rect 25412 19660 25464 19712
rect 34612 19703 34664 19712
rect 34612 19669 34621 19703
rect 34621 19669 34655 19703
rect 34655 19669 34664 19703
rect 34612 19660 34664 19669
rect 35256 19703 35308 19712
rect 35256 19669 35265 19703
rect 35265 19669 35299 19703
rect 35299 19669 35308 19703
rect 35256 19660 35308 19669
rect 41420 19703 41472 19712
rect 41420 19669 41429 19703
rect 41429 19669 41463 19703
rect 41463 19669 41472 19703
rect 41420 19660 41472 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 20904 19456 20956 19508
rect 23388 19499 23440 19508
rect 23388 19465 23397 19499
rect 23397 19465 23431 19499
rect 23431 19465 23440 19499
rect 23388 19456 23440 19465
rect 24952 19499 25004 19508
rect 24952 19465 24961 19499
rect 24961 19465 24995 19499
rect 24995 19465 25004 19499
rect 24952 19456 25004 19465
rect 25688 19499 25740 19508
rect 25688 19465 25697 19499
rect 25697 19465 25731 19499
rect 25731 19465 25740 19499
rect 25688 19456 25740 19465
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 27252 19499 27304 19508
rect 27252 19465 27261 19499
rect 27261 19465 27295 19499
rect 27295 19465 27304 19499
rect 27252 19456 27304 19465
rect 30840 19456 30892 19508
rect 30932 19499 30984 19508
rect 30932 19465 30941 19499
rect 30941 19465 30975 19499
rect 30975 19465 30984 19499
rect 30932 19456 30984 19465
rect 31116 19456 31168 19508
rect 33508 19456 33560 19508
rect 35624 19456 35676 19508
rect 38384 19499 38436 19508
rect 38384 19465 38393 19499
rect 38393 19465 38427 19499
rect 38427 19465 38436 19499
rect 38384 19456 38436 19465
rect 38936 19499 38988 19508
rect 38936 19465 38945 19499
rect 38945 19465 38979 19499
rect 38979 19465 38988 19499
rect 38936 19456 38988 19465
rect 41328 19456 41380 19508
rect 41880 19456 41932 19508
rect 44824 19456 44876 19508
rect 45836 19456 45888 19508
rect 18052 19388 18104 19440
rect 25412 19388 25464 19440
rect 26884 19388 26936 19440
rect 36452 19388 36504 19440
rect 36636 19388 36688 19440
rect 39304 19388 39356 19440
rect 20260 19363 20312 19372
rect 16488 19252 16540 19304
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 20720 19320 20772 19372
rect 18512 19295 18564 19304
rect 17132 19227 17184 19236
rect 17132 19193 17141 19227
rect 17141 19193 17175 19227
rect 17175 19193 17184 19227
rect 17132 19184 17184 19193
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 19248 19252 19300 19304
rect 22652 19320 22704 19372
rect 23756 19320 23808 19372
rect 34704 19320 34756 19372
rect 35256 19320 35308 19372
rect 37648 19320 37700 19372
rect 37924 19320 37976 19372
rect 23112 19252 23164 19304
rect 23664 19295 23716 19304
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 20260 19184 20312 19236
rect 20628 19184 20680 19236
rect 21272 19184 21324 19236
rect 23296 19184 23348 19236
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 26240 19227 26292 19236
rect 26240 19193 26249 19227
rect 26249 19193 26283 19227
rect 26283 19193 26292 19227
rect 26240 19184 26292 19193
rect 27804 19227 27856 19236
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 21364 19159 21416 19168
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 21364 19116 21416 19125
rect 22744 19159 22796 19168
rect 22744 19125 22753 19159
rect 22753 19125 22787 19159
rect 22787 19125 22796 19159
rect 22744 19116 22796 19125
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 23940 19116 23992 19168
rect 26056 19116 26108 19168
rect 27804 19193 27813 19227
rect 27813 19193 27847 19227
rect 27847 19193 27856 19227
rect 27804 19184 27856 19193
rect 30104 19252 30156 19304
rect 30748 19252 30800 19304
rect 32404 19252 32456 19304
rect 34520 19252 34572 19304
rect 36176 19252 36228 19304
rect 37464 19184 37516 19236
rect 37556 19227 37608 19236
rect 37556 19193 37565 19227
rect 37565 19193 37599 19227
rect 37599 19193 37608 19227
rect 37556 19184 37608 19193
rect 38200 19184 38252 19236
rect 41420 19227 41472 19236
rect 41420 19193 41429 19227
rect 41429 19193 41463 19227
rect 41463 19193 41472 19227
rect 41420 19184 41472 19193
rect 43260 19320 43312 19372
rect 43628 19363 43680 19372
rect 43628 19329 43637 19363
rect 43637 19329 43671 19363
rect 43671 19329 43680 19363
rect 43628 19320 43680 19329
rect 42984 19227 43036 19236
rect 31484 19159 31536 19168
rect 31484 19125 31493 19159
rect 31493 19125 31527 19159
rect 31527 19125 31536 19159
rect 31484 19116 31536 19125
rect 31944 19159 31996 19168
rect 31944 19125 31953 19159
rect 31953 19125 31987 19159
rect 31987 19125 31996 19159
rect 31944 19116 31996 19125
rect 32404 19116 32456 19168
rect 33140 19116 33192 19168
rect 33416 19116 33468 19168
rect 33600 19159 33652 19168
rect 33600 19125 33609 19159
rect 33609 19125 33643 19159
rect 33643 19125 33652 19159
rect 33600 19116 33652 19125
rect 33876 19159 33928 19168
rect 33876 19125 33885 19159
rect 33885 19125 33919 19159
rect 33919 19125 33928 19159
rect 33876 19116 33928 19125
rect 34520 19159 34572 19168
rect 34520 19125 34529 19159
rect 34529 19125 34563 19159
rect 34563 19125 34572 19159
rect 34520 19116 34572 19125
rect 35624 19116 35676 19168
rect 41328 19116 41380 19168
rect 42984 19193 42993 19227
rect 42993 19193 43027 19227
rect 43027 19193 43036 19227
rect 42984 19184 43036 19193
rect 42616 19116 42668 19168
rect 43444 19184 43496 19236
rect 45192 19184 45244 19236
rect 46756 19184 46808 19236
rect 43720 19116 43772 19168
rect 45008 19159 45060 19168
rect 45008 19125 45017 19159
rect 45017 19125 45051 19159
rect 45051 19125 45060 19159
rect 45008 19116 45060 19125
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 16856 18955 16908 18964
rect 16856 18921 16865 18955
rect 16865 18921 16899 18955
rect 16899 18921 16908 18955
rect 16856 18912 16908 18921
rect 17408 18912 17460 18964
rect 17776 18955 17828 18964
rect 17776 18921 17785 18955
rect 17785 18921 17819 18955
rect 17819 18921 17828 18955
rect 17776 18912 17828 18921
rect 18512 18912 18564 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 29000 18955 29052 18964
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 21364 18844 21416 18896
rect 21548 18844 21600 18896
rect 26700 18887 26752 18896
rect 26700 18853 26709 18887
rect 26709 18853 26743 18887
rect 26743 18853 26752 18887
rect 26700 18844 26752 18853
rect 27804 18844 27856 18896
rect 32036 18912 32088 18964
rect 32404 18912 32456 18964
rect 34612 18912 34664 18964
rect 34796 18912 34848 18964
rect 35348 18955 35400 18964
rect 35348 18921 35357 18955
rect 35357 18921 35391 18955
rect 35391 18921 35400 18955
rect 35348 18912 35400 18921
rect 37556 18912 37608 18964
rect 41604 18912 41656 18964
rect 43168 18912 43220 18964
rect 29828 18844 29880 18896
rect 30564 18887 30616 18896
rect 30564 18853 30573 18887
rect 30573 18853 30607 18887
rect 30607 18853 30616 18887
rect 30564 18844 30616 18853
rect 34704 18887 34756 18896
rect 17132 18776 17184 18828
rect 19432 18776 19484 18828
rect 22744 18776 22796 18828
rect 23112 18819 23164 18828
rect 23112 18785 23121 18819
rect 23121 18785 23155 18819
rect 23155 18785 23164 18819
rect 23112 18776 23164 18785
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 28356 18776 28408 18828
rect 29276 18776 29328 18828
rect 30748 18819 30800 18828
rect 30748 18785 30757 18819
rect 30757 18785 30791 18819
rect 30791 18785 30800 18819
rect 30748 18776 30800 18785
rect 31852 18776 31904 18828
rect 34704 18853 34713 18887
rect 34713 18853 34747 18887
rect 34747 18853 34756 18887
rect 34704 18844 34756 18853
rect 35624 18844 35676 18896
rect 37648 18844 37700 18896
rect 38016 18887 38068 18896
rect 38016 18853 38025 18887
rect 38025 18853 38059 18887
rect 38059 18853 38068 18887
rect 38016 18844 38068 18853
rect 40960 18844 41012 18896
rect 43628 18844 43680 18896
rect 45100 18844 45152 18896
rect 45560 18887 45612 18896
rect 45560 18853 45569 18887
rect 45569 18853 45603 18887
rect 45603 18853 45612 18887
rect 45560 18844 45612 18853
rect 46480 18887 46532 18896
rect 46480 18853 46489 18887
rect 46489 18853 46523 18887
rect 46523 18853 46532 18887
rect 46480 18844 46532 18853
rect 46572 18887 46624 18896
rect 46572 18853 46581 18887
rect 46581 18853 46615 18887
rect 46615 18853 46624 18887
rect 46572 18844 46624 18853
rect 32772 18776 32824 18828
rect 33508 18776 33560 18828
rect 34336 18776 34388 18828
rect 21548 18708 21600 18760
rect 26608 18751 26660 18760
rect 26608 18717 26617 18751
rect 26617 18717 26651 18751
rect 26651 18717 26660 18751
rect 26608 18708 26660 18717
rect 27620 18708 27672 18760
rect 30840 18708 30892 18760
rect 22744 18640 22796 18692
rect 31484 18640 31536 18692
rect 34060 18640 34112 18692
rect 38200 18776 38252 18828
rect 39948 18776 40000 18828
rect 40040 18776 40092 18828
rect 41696 18776 41748 18828
rect 42800 18776 42852 18828
rect 35348 18708 35400 18760
rect 37740 18751 37792 18760
rect 37740 18717 37749 18751
rect 37749 18717 37783 18751
rect 37783 18717 37792 18751
rect 37740 18708 37792 18717
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 20720 18572 20772 18624
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 26240 18572 26292 18581
rect 27896 18572 27948 18624
rect 29552 18572 29604 18624
rect 32312 18572 32364 18624
rect 43720 18708 43772 18760
rect 44916 18751 44968 18760
rect 44916 18717 44925 18751
rect 44925 18717 44959 18751
rect 44959 18717 44968 18751
rect 44916 18708 44968 18717
rect 46756 18751 46808 18760
rect 46756 18717 46765 18751
rect 46765 18717 46799 18751
rect 46799 18717 46808 18751
rect 46756 18708 46808 18717
rect 36820 18572 36872 18624
rect 39764 18572 39816 18624
rect 40500 18615 40552 18624
rect 40500 18581 40509 18615
rect 40509 18581 40543 18615
rect 40543 18581 40552 18615
rect 40500 18572 40552 18581
rect 43628 18615 43680 18624
rect 43628 18581 43637 18615
rect 43637 18581 43671 18615
rect 43671 18581 43680 18615
rect 43628 18572 43680 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 17132 18411 17184 18420
rect 17132 18377 17141 18411
rect 17141 18377 17175 18411
rect 17175 18377 17184 18411
rect 17132 18368 17184 18377
rect 17776 18368 17828 18420
rect 21364 18368 21416 18420
rect 21548 18411 21600 18420
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 22744 18411 22796 18420
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 24952 18368 25004 18420
rect 25136 18411 25188 18420
rect 25136 18377 25145 18411
rect 25145 18377 25179 18411
rect 25179 18377 25188 18411
rect 25136 18368 25188 18377
rect 25596 18411 25648 18420
rect 25596 18377 25605 18411
rect 25605 18377 25639 18411
rect 25639 18377 25648 18411
rect 25596 18368 25648 18377
rect 26700 18411 26752 18420
rect 26700 18377 26709 18411
rect 26709 18377 26743 18411
rect 26743 18377 26752 18411
rect 26700 18368 26752 18377
rect 29276 18368 29328 18420
rect 30748 18368 30800 18420
rect 31852 18411 31904 18420
rect 31852 18377 31861 18411
rect 31861 18377 31895 18411
rect 31895 18377 31904 18411
rect 31852 18368 31904 18377
rect 36452 18368 36504 18420
rect 18696 18343 18748 18352
rect 18696 18309 18705 18343
rect 18705 18309 18739 18343
rect 18739 18309 18748 18343
rect 18696 18300 18748 18309
rect 18512 18232 18564 18284
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 25044 18300 25096 18352
rect 29184 18300 29236 18352
rect 34796 18300 34848 18352
rect 27620 18275 27672 18284
rect 19984 18164 20036 18216
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 29828 18275 29880 18284
rect 29828 18241 29837 18275
rect 29837 18241 29871 18275
rect 29871 18241 29880 18275
rect 29828 18232 29880 18241
rect 31852 18232 31904 18284
rect 32864 18232 32916 18284
rect 33232 18232 33284 18284
rect 18328 18096 18380 18148
rect 20076 18096 20128 18148
rect 22560 18164 22612 18216
rect 25136 18164 25188 18216
rect 29552 18164 29604 18216
rect 30840 18164 30892 18216
rect 32404 18164 32456 18216
rect 32772 18207 32824 18216
rect 32772 18173 32781 18207
rect 32781 18173 32815 18207
rect 32815 18173 32824 18207
rect 32772 18164 32824 18173
rect 25780 18139 25832 18148
rect 25780 18105 25789 18139
rect 25789 18105 25823 18139
rect 25823 18105 25832 18139
rect 25780 18096 25832 18105
rect 19432 18028 19484 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 21916 18071 21968 18080
rect 21916 18037 21925 18071
rect 21925 18037 21959 18071
rect 21959 18037 21968 18071
rect 21916 18028 21968 18037
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 23940 18028 23992 18080
rect 24216 18071 24268 18080
rect 24216 18037 24225 18071
rect 24225 18037 24259 18071
rect 24259 18037 24268 18071
rect 24216 18028 24268 18037
rect 25596 18028 25648 18080
rect 26240 18096 26292 18148
rect 26792 18096 26844 18148
rect 27344 18139 27396 18148
rect 27344 18105 27353 18139
rect 27353 18105 27387 18139
rect 27387 18105 27396 18139
rect 27344 18096 27396 18105
rect 31116 18139 31168 18148
rect 28356 18071 28408 18080
rect 28356 18037 28365 18071
rect 28365 18037 28399 18071
rect 28399 18037 28408 18071
rect 28356 18028 28408 18037
rect 29368 18028 29420 18080
rect 31116 18105 31125 18139
rect 31125 18105 31159 18139
rect 31159 18105 31168 18139
rect 31116 18096 31168 18105
rect 31208 18096 31260 18148
rect 33324 18139 33376 18148
rect 33324 18105 33333 18139
rect 33333 18105 33367 18139
rect 33367 18105 33376 18139
rect 33324 18096 33376 18105
rect 34796 18164 34848 18216
rect 37740 18368 37792 18420
rect 38936 18368 38988 18420
rect 41328 18368 41380 18420
rect 41696 18411 41748 18420
rect 41696 18377 41705 18411
rect 41705 18377 41739 18411
rect 41739 18377 41748 18411
rect 41696 18368 41748 18377
rect 42800 18368 42852 18420
rect 45008 18368 45060 18420
rect 38016 18300 38068 18352
rect 37556 18232 37608 18284
rect 39212 18232 39264 18284
rect 35808 18207 35860 18216
rect 35808 18173 35817 18207
rect 35817 18173 35851 18207
rect 35851 18173 35860 18207
rect 35808 18164 35860 18173
rect 36452 18207 36504 18216
rect 36452 18173 36461 18207
rect 36461 18173 36495 18207
rect 36495 18173 36504 18207
rect 36452 18164 36504 18173
rect 36820 18207 36872 18216
rect 36820 18173 36829 18207
rect 36829 18173 36863 18207
rect 36863 18173 36872 18207
rect 36820 18164 36872 18173
rect 36912 18164 36964 18216
rect 38936 18164 38988 18216
rect 39396 18164 39448 18216
rect 39672 18164 39724 18216
rect 40500 18207 40552 18216
rect 40500 18173 40509 18207
rect 40509 18173 40543 18207
rect 40543 18173 40552 18207
rect 40500 18164 40552 18173
rect 44916 18300 44968 18352
rect 43352 18232 43404 18284
rect 43812 18232 43864 18284
rect 46848 18275 46900 18284
rect 46848 18241 46857 18275
rect 46857 18241 46891 18275
rect 46891 18241 46900 18275
rect 46848 18232 46900 18241
rect 43444 18164 43496 18216
rect 45928 18164 45980 18216
rect 37648 18096 37700 18148
rect 38016 18096 38068 18148
rect 40684 18096 40736 18148
rect 40960 18096 41012 18148
rect 43628 18096 43680 18148
rect 31484 18071 31536 18080
rect 31484 18037 31493 18071
rect 31493 18037 31527 18071
rect 31527 18037 31536 18071
rect 31484 18028 31536 18037
rect 33600 18071 33652 18080
rect 33600 18037 33609 18071
rect 33609 18037 33643 18071
rect 33643 18037 33652 18071
rect 33600 18028 33652 18037
rect 34244 18071 34296 18080
rect 34244 18037 34253 18071
rect 34253 18037 34287 18071
rect 34287 18037 34296 18071
rect 34244 18028 34296 18037
rect 34336 18028 34388 18080
rect 35256 18028 35308 18080
rect 38292 18028 38344 18080
rect 45100 18028 45152 18080
rect 46204 18028 46256 18080
rect 46572 18028 46624 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 20996 17867 21048 17876
rect 20996 17833 21005 17867
rect 21005 17833 21039 17867
rect 21039 17833 21048 17867
rect 20996 17824 21048 17833
rect 26608 17824 26660 17876
rect 27344 17824 27396 17876
rect 28356 17824 28408 17876
rect 33324 17867 33376 17876
rect 33324 17833 33333 17867
rect 33333 17833 33367 17867
rect 33367 17833 33376 17867
rect 33324 17824 33376 17833
rect 34060 17867 34112 17876
rect 34060 17833 34069 17867
rect 34069 17833 34103 17867
rect 34103 17833 34112 17867
rect 34060 17824 34112 17833
rect 35624 17867 35676 17876
rect 35624 17833 35633 17867
rect 35633 17833 35667 17867
rect 35667 17833 35676 17867
rect 35624 17824 35676 17833
rect 36452 17824 36504 17876
rect 39948 17867 40000 17876
rect 39948 17833 39957 17867
rect 39957 17833 39991 17867
rect 39991 17833 40000 17867
rect 39948 17824 40000 17833
rect 40040 17824 40092 17876
rect 43444 17824 43496 17876
rect 43536 17824 43588 17876
rect 46204 17867 46256 17876
rect 17776 17756 17828 17808
rect 26700 17799 26752 17808
rect 16856 17688 16908 17740
rect 18144 17688 18196 17740
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 26700 17765 26709 17799
rect 26709 17765 26743 17799
rect 26743 17765 26752 17799
rect 26700 17756 26752 17765
rect 26792 17756 26844 17808
rect 29184 17799 29236 17808
rect 29184 17765 29193 17799
rect 29193 17765 29227 17799
rect 29227 17765 29236 17799
rect 29184 17756 29236 17765
rect 30564 17799 30616 17808
rect 30564 17765 30573 17799
rect 30573 17765 30607 17799
rect 30607 17765 30616 17799
rect 30564 17756 30616 17765
rect 31484 17756 31536 17808
rect 32772 17756 32824 17808
rect 46204 17833 46213 17867
rect 46213 17833 46247 17867
rect 46247 17833 46256 17867
rect 46204 17824 46256 17833
rect 46480 17867 46532 17876
rect 46480 17833 46489 17867
rect 46489 17833 46523 17867
rect 46523 17833 46532 17867
rect 46480 17824 46532 17833
rect 38660 17756 38712 17808
rect 39672 17799 39724 17808
rect 19892 17663 19944 17672
rect 19892 17629 19901 17663
rect 19901 17629 19935 17663
rect 19935 17629 19944 17663
rect 19892 17620 19944 17629
rect 20352 17620 20404 17672
rect 21180 17688 21232 17740
rect 21916 17688 21968 17740
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 24216 17688 24268 17740
rect 25044 17688 25096 17740
rect 25504 17688 25556 17740
rect 28264 17688 28316 17740
rect 29276 17688 29328 17740
rect 30656 17731 30708 17740
rect 30656 17697 30665 17731
rect 30665 17697 30699 17731
rect 30699 17697 30708 17731
rect 30656 17688 30708 17697
rect 30840 17731 30892 17740
rect 30840 17697 30849 17731
rect 30849 17697 30883 17731
rect 30883 17697 30892 17731
rect 30840 17688 30892 17697
rect 32220 17688 32272 17740
rect 34520 17731 34572 17740
rect 34520 17697 34529 17731
rect 34529 17697 34563 17731
rect 34563 17697 34572 17731
rect 34520 17688 34572 17697
rect 35348 17688 35400 17740
rect 37648 17688 37700 17740
rect 39672 17765 39681 17799
rect 39681 17765 39715 17799
rect 39715 17765 39724 17799
rect 39672 17756 39724 17765
rect 40960 17756 41012 17808
rect 44916 17799 44968 17808
rect 44916 17765 44925 17799
rect 44925 17765 44959 17799
rect 44959 17765 44968 17799
rect 44916 17756 44968 17765
rect 45100 17756 45152 17808
rect 45468 17799 45520 17808
rect 45468 17765 45477 17799
rect 45477 17765 45511 17799
rect 45511 17765 45520 17799
rect 45468 17756 45520 17765
rect 39396 17731 39448 17740
rect 39396 17697 39405 17731
rect 39405 17697 39439 17731
rect 39439 17697 39448 17731
rect 39396 17688 39448 17697
rect 43260 17731 43312 17740
rect 43260 17697 43269 17731
rect 43269 17697 43303 17731
rect 43303 17697 43312 17731
rect 43260 17688 43312 17697
rect 22744 17620 22796 17672
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 22284 17552 22336 17604
rect 34244 17620 34296 17672
rect 35532 17620 35584 17672
rect 40592 17663 40644 17672
rect 40592 17629 40601 17663
rect 40601 17629 40635 17663
rect 40635 17629 40644 17663
rect 40592 17620 40644 17629
rect 44824 17663 44876 17672
rect 44824 17629 44833 17663
rect 44833 17629 44867 17663
rect 44867 17629 44876 17663
rect 44824 17620 44876 17629
rect 31576 17595 31628 17604
rect 31576 17561 31585 17595
rect 31585 17561 31619 17595
rect 31619 17561 31628 17595
rect 31576 17552 31628 17561
rect 32496 17552 32548 17604
rect 18236 17484 18288 17536
rect 18512 17527 18564 17536
rect 18512 17493 18521 17527
rect 18521 17493 18555 17527
rect 18555 17493 18564 17527
rect 18512 17484 18564 17493
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 24584 17527 24636 17536
rect 24584 17493 24593 17527
rect 24593 17493 24627 17527
rect 24627 17493 24636 17527
rect 24584 17484 24636 17493
rect 25688 17484 25740 17536
rect 25780 17484 25832 17536
rect 29460 17484 29512 17536
rect 30104 17527 30156 17536
rect 30104 17493 30113 17527
rect 30113 17493 30147 17527
rect 30147 17493 30156 17527
rect 30104 17484 30156 17493
rect 30932 17527 30984 17536
rect 30932 17493 30941 17527
rect 30941 17493 30975 17527
rect 30975 17493 30984 17527
rect 30932 17484 30984 17493
rect 32404 17484 32456 17536
rect 36544 17527 36596 17536
rect 36544 17493 36553 17527
rect 36553 17493 36587 17527
rect 36587 17493 36596 17527
rect 36544 17484 36596 17493
rect 37924 17527 37976 17536
rect 37924 17493 37933 17527
rect 37933 17493 37967 17527
rect 37967 17493 37976 17527
rect 37924 17484 37976 17493
rect 43260 17484 43312 17536
rect 43628 17484 43680 17536
rect 43812 17527 43864 17536
rect 43812 17493 43821 17527
rect 43821 17493 43855 17527
rect 43855 17493 43864 17527
rect 43812 17484 43864 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 16856 17280 16908 17289
rect 18512 17280 18564 17332
rect 18604 17280 18656 17332
rect 20352 17323 20404 17332
rect 20352 17289 20361 17323
rect 20361 17289 20395 17323
rect 20395 17289 20404 17323
rect 20352 17280 20404 17289
rect 20628 17323 20680 17332
rect 20628 17289 20637 17323
rect 20637 17289 20671 17323
rect 20671 17289 20680 17323
rect 20628 17280 20680 17289
rect 22744 17323 22796 17332
rect 22744 17289 22753 17323
rect 22753 17289 22787 17323
rect 22787 17289 22796 17323
rect 22744 17280 22796 17289
rect 23388 17323 23440 17332
rect 23388 17289 23397 17323
rect 23397 17289 23431 17323
rect 23431 17289 23440 17323
rect 23388 17280 23440 17289
rect 23940 17323 23992 17332
rect 23940 17289 23949 17323
rect 23949 17289 23983 17323
rect 23983 17289 23992 17323
rect 23940 17280 23992 17289
rect 25044 17323 25096 17332
rect 25044 17289 25053 17323
rect 25053 17289 25087 17323
rect 25087 17289 25096 17323
rect 25044 17280 25096 17289
rect 26700 17280 26752 17332
rect 29276 17280 29328 17332
rect 30656 17323 30708 17332
rect 30656 17289 30665 17323
rect 30665 17289 30699 17323
rect 30699 17289 30708 17323
rect 30656 17280 30708 17289
rect 31300 17280 31352 17332
rect 32220 17280 32272 17332
rect 34520 17323 34572 17332
rect 34520 17289 34529 17323
rect 34529 17289 34563 17323
rect 34563 17289 34572 17323
rect 34520 17280 34572 17289
rect 17776 17212 17828 17264
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 18880 17144 18932 17196
rect 20996 17144 21048 17196
rect 20352 17076 20404 17128
rect 18236 17051 18288 17060
rect 18236 17017 18245 17051
rect 18245 17017 18279 17051
rect 18279 17017 18288 17051
rect 18236 17008 18288 17017
rect 19524 17008 19576 17060
rect 20076 17008 20128 17060
rect 20628 17008 20680 17060
rect 23940 17076 23992 17128
rect 25964 17212 26016 17264
rect 27712 17212 27764 17264
rect 29736 17212 29788 17264
rect 31668 17212 31720 17264
rect 26608 17144 26660 17196
rect 29184 17144 29236 17196
rect 30104 17144 30156 17196
rect 34152 17212 34204 17264
rect 36912 17280 36964 17332
rect 37648 17280 37700 17332
rect 38292 17323 38344 17332
rect 38292 17289 38301 17323
rect 38301 17289 38335 17323
rect 38335 17289 38344 17323
rect 38292 17280 38344 17289
rect 38660 17323 38712 17332
rect 38660 17289 38669 17323
rect 38669 17289 38703 17323
rect 38703 17289 38712 17323
rect 38660 17280 38712 17289
rect 39396 17280 39448 17332
rect 42616 17323 42668 17332
rect 42616 17289 42625 17323
rect 42625 17289 42659 17323
rect 42659 17289 42668 17323
rect 42616 17280 42668 17289
rect 43260 17323 43312 17332
rect 43260 17289 43269 17323
rect 43269 17289 43303 17323
rect 43303 17289 43312 17323
rect 43260 17280 43312 17289
rect 44824 17280 44876 17332
rect 35440 17212 35492 17264
rect 36360 17255 36412 17264
rect 36360 17221 36369 17255
rect 36369 17221 36403 17255
rect 36403 17221 36412 17255
rect 36360 17212 36412 17221
rect 36544 17255 36596 17264
rect 36544 17221 36553 17255
rect 36553 17221 36587 17255
rect 36587 17221 36596 17255
rect 36544 17212 36596 17221
rect 34612 17144 34664 17196
rect 40592 17212 40644 17264
rect 43168 17212 43220 17264
rect 31576 17076 31628 17128
rect 24952 17008 25004 17060
rect 26148 17008 26200 17060
rect 18420 16940 18472 16992
rect 19340 16940 19392 16992
rect 21548 16940 21600 16992
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 25504 16983 25556 16992
rect 25504 16949 25513 16983
rect 25513 16949 25547 16983
rect 25547 16949 25556 16983
rect 25504 16940 25556 16949
rect 25872 16940 25924 16992
rect 25964 16940 26016 16992
rect 26792 16983 26844 16992
rect 26792 16949 26801 16983
rect 26801 16949 26835 16983
rect 26835 16949 26844 16983
rect 26792 16940 26844 16949
rect 27252 17008 27304 17060
rect 30840 17008 30892 17060
rect 32036 17076 32088 17128
rect 32404 17076 32456 17128
rect 34336 17076 34388 17128
rect 40684 17144 40736 17196
rect 41696 17187 41748 17196
rect 41696 17153 41705 17187
rect 41705 17153 41739 17187
rect 41739 17153 41748 17187
rect 41696 17144 41748 17153
rect 44916 17144 44968 17196
rect 35532 17076 35584 17128
rect 36360 17076 36412 17128
rect 38292 17076 38344 17128
rect 39396 17119 39448 17128
rect 39396 17085 39405 17119
rect 39405 17085 39439 17119
rect 39439 17085 39448 17119
rect 39396 17076 39448 17085
rect 45192 17076 45244 17128
rect 27712 16940 27764 16992
rect 29000 16983 29052 16992
rect 29000 16949 29009 16983
rect 29009 16949 29043 16983
rect 29043 16949 29052 16983
rect 29000 16940 29052 16949
rect 32496 16940 32548 16992
rect 32772 16940 32824 16992
rect 33416 16983 33468 16992
rect 33416 16949 33425 16983
rect 33425 16949 33459 16983
rect 33459 16949 33468 16983
rect 33416 16940 33468 16949
rect 34796 16940 34848 16992
rect 35348 16983 35400 16992
rect 35348 16949 35357 16983
rect 35357 16949 35391 16983
rect 35391 16949 35400 16983
rect 35348 16940 35400 16949
rect 36360 16940 36412 16992
rect 40224 16983 40276 16992
rect 40224 16949 40233 16983
rect 40233 16949 40267 16983
rect 40267 16949 40276 16983
rect 40224 16940 40276 16949
rect 40316 16940 40368 16992
rect 40960 16983 41012 16992
rect 40960 16949 40969 16983
rect 40969 16949 41003 16983
rect 41003 16949 41012 16983
rect 43536 17051 43588 17060
rect 43536 17017 43545 17051
rect 43545 17017 43579 17051
rect 43579 17017 43588 17051
rect 43536 17008 43588 17017
rect 40960 16940 41012 16949
rect 43260 16940 43312 16992
rect 44640 17008 44692 17060
rect 46388 16940 46440 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 18144 16736 18196 16788
rect 16948 16600 17000 16652
rect 17500 16600 17552 16652
rect 18604 16668 18656 16720
rect 18512 16600 18564 16652
rect 19340 16736 19392 16788
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 23388 16736 23440 16788
rect 26608 16736 26660 16788
rect 27712 16779 27764 16788
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 19708 16600 19760 16652
rect 21548 16711 21600 16720
rect 21548 16677 21557 16711
rect 21557 16677 21591 16711
rect 21591 16677 21600 16711
rect 21548 16668 21600 16677
rect 26792 16668 26844 16720
rect 26884 16711 26936 16720
rect 26884 16677 26893 16711
rect 26893 16677 26927 16711
rect 26927 16677 26936 16711
rect 27712 16745 27721 16779
rect 27721 16745 27755 16779
rect 27755 16745 27764 16779
rect 27712 16736 27764 16745
rect 34336 16779 34388 16788
rect 34336 16745 34345 16779
rect 34345 16745 34379 16779
rect 34379 16745 34388 16779
rect 34336 16736 34388 16745
rect 35348 16736 35400 16788
rect 36912 16736 36964 16788
rect 37924 16736 37976 16788
rect 39396 16736 39448 16788
rect 40592 16736 40644 16788
rect 41696 16779 41748 16788
rect 41696 16745 41705 16779
rect 41705 16745 41739 16779
rect 41739 16745 41748 16779
rect 41696 16736 41748 16745
rect 43536 16736 43588 16788
rect 44824 16736 44876 16788
rect 26884 16668 26936 16677
rect 29092 16668 29144 16720
rect 36544 16668 36596 16720
rect 38016 16668 38068 16720
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 24584 16643 24636 16652
rect 24584 16609 24593 16643
rect 24593 16609 24627 16643
rect 24627 16609 24636 16643
rect 24584 16600 24636 16609
rect 31116 16600 31168 16652
rect 32220 16600 32272 16652
rect 33508 16600 33560 16652
rect 34152 16643 34204 16652
rect 34152 16609 34161 16643
rect 34161 16609 34195 16643
rect 34195 16609 34204 16643
rect 34152 16600 34204 16609
rect 35808 16643 35860 16652
rect 35808 16609 35817 16643
rect 35817 16609 35851 16643
rect 35851 16609 35860 16643
rect 35808 16600 35860 16609
rect 39580 16643 39632 16652
rect 39580 16609 39589 16643
rect 39589 16609 39623 16643
rect 39623 16609 39632 16643
rect 39580 16600 39632 16609
rect 43812 16668 43864 16720
rect 47308 16668 47360 16720
rect 41144 16643 41196 16652
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 27068 16532 27120 16584
rect 28356 16532 28408 16584
rect 31668 16532 31720 16584
rect 33416 16532 33468 16584
rect 33692 16532 33744 16584
rect 37832 16575 37884 16584
rect 37832 16541 37841 16575
rect 37841 16541 37875 16575
rect 37875 16541 37884 16575
rect 37832 16532 37884 16541
rect 20352 16507 20404 16516
rect 20352 16473 20361 16507
rect 20361 16473 20395 16507
rect 20395 16473 20404 16507
rect 20352 16464 20404 16473
rect 27896 16464 27948 16516
rect 41144 16609 41188 16643
rect 41188 16609 41196 16643
rect 41144 16600 41196 16609
rect 42432 16600 42484 16652
rect 43444 16643 43496 16652
rect 43444 16609 43462 16643
rect 43462 16609 43496 16643
rect 43444 16600 43496 16609
rect 43904 16600 43956 16652
rect 44640 16643 44692 16652
rect 44640 16609 44649 16643
rect 44649 16609 44683 16643
rect 44683 16609 44692 16643
rect 44640 16600 44692 16609
rect 45560 16600 45612 16652
rect 47216 16643 47268 16652
rect 47216 16609 47225 16643
rect 47225 16609 47259 16643
rect 47259 16609 47268 16643
rect 47216 16600 47268 16609
rect 42340 16532 42392 16584
rect 40592 16464 40644 16516
rect 44272 16464 44324 16516
rect 45560 16464 45612 16516
rect 25228 16439 25280 16448
rect 25228 16405 25237 16439
rect 25237 16405 25271 16439
rect 25271 16405 25280 16439
rect 25228 16396 25280 16405
rect 28264 16439 28316 16448
rect 28264 16405 28273 16439
rect 28273 16405 28307 16439
rect 28307 16405 28316 16439
rect 28264 16396 28316 16405
rect 30380 16396 30432 16448
rect 31208 16439 31260 16448
rect 31208 16405 31217 16439
rect 31217 16405 31251 16439
rect 31251 16405 31260 16439
rect 31208 16396 31260 16405
rect 31576 16439 31628 16448
rect 31576 16405 31585 16439
rect 31585 16405 31619 16439
rect 31619 16405 31628 16439
rect 31576 16396 31628 16405
rect 32036 16396 32088 16448
rect 34520 16396 34572 16448
rect 35532 16396 35584 16448
rect 42156 16396 42208 16448
rect 43720 16396 43772 16448
rect 46296 16396 46348 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 19248 16235 19300 16244
rect 19248 16201 19257 16235
rect 19257 16201 19291 16235
rect 19291 16201 19300 16235
rect 19248 16192 19300 16201
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 20628 16192 20680 16244
rect 21548 16192 21600 16244
rect 24584 16192 24636 16244
rect 25964 16192 26016 16244
rect 26148 16235 26200 16244
rect 26148 16201 26157 16235
rect 26157 16201 26191 16235
rect 26191 16201 26200 16235
rect 26148 16192 26200 16201
rect 26884 16192 26936 16244
rect 30380 16235 30432 16244
rect 30380 16201 30389 16235
rect 30389 16201 30423 16235
rect 30423 16201 30432 16235
rect 30380 16192 30432 16201
rect 31116 16192 31168 16244
rect 31668 16235 31720 16244
rect 31668 16201 31677 16235
rect 31677 16201 31711 16235
rect 31711 16201 31720 16235
rect 31668 16192 31720 16201
rect 34152 16192 34204 16244
rect 35808 16192 35860 16244
rect 21088 16124 21140 16176
rect 22468 16124 22520 16176
rect 22928 16167 22980 16176
rect 22928 16133 22937 16167
rect 22937 16133 22971 16167
rect 22971 16133 22980 16167
rect 22928 16124 22980 16133
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 19984 16056 20036 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 21456 16056 21508 16108
rect 25228 16056 25280 16108
rect 25688 16056 25740 16108
rect 34244 16124 34296 16176
rect 35256 16124 35308 16176
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 29736 16099 29788 16108
rect 29736 16065 29745 16099
rect 29745 16065 29779 16099
rect 29779 16065 29788 16099
rect 29736 16056 29788 16065
rect 30104 16056 30156 16108
rect 33324 16056 33376 16108
rect 33876 16056 33928 16108
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 22468 16031 22520 16040
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 23296 15988 23348 16040
rect 20628 15920 20680 15972
rect 26148 15920 26200 15972
rect 30380 15988 30432 16040
rect 32128 16031 32180 16040
rect 32128 15997 32137 16031
rect 32137 15997 32171 16031
rect 32171 15997 32180 16031
rect 32128 15988 32180 15997
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 34704 15988 34756 16040
rect 35348 15988 35400 16040
rect 36360 16192 36412 16244
rect 40224 16192 40276 16244
rect 42432 16192 42484 16244
rect 43444 16235 43496 16244
rect 39396 16124 39448 16176
rect 39580 16167 39632 16176
rect 39580 16133 39589 16167
rect 39589 16133 39623 16167
rect 39623 16133 39632 16167
rect 39580 16124 39632 16133
rect 43444 16201 43453 16235
rect 43453 16201 43487 16235
rect 43487 16201 43496 16235
rect 43444 16192 43496 16201
rect 44640 16235 44692 16244
rect 44640 16201 44649 16235
rect 44649 16201 44683 16235
rect 44683 16201 44692 16235
rect 44640 16192 44692 16201
rect 45560 16235 45612 16244
rect 45560 16201 45569 16235
rect 45569 16201 45603 16235
rect 45603 16201 45612 16235
rect 45560 16192 45612 16201
rect 47216 16167 47268 16176
rect 47216 16133 47225 16167
rect 47225 16133 47259 16167
rect 47259 16133 47268 16167
rect 47216 16124 47268 16133
rect 40592 16099 40644 16108
rect 40592 16065 40601 16099
rect 40601 16065 40635 16099
rect 40635 16065 40644 16099
rect 40592 16056 40644 16065
rect 40776 16056 40828 16108
rect 36912 16031 36964 16040
rect 33508 15920 33560 15972
rect 16948 15852 17000 15904
rect 21364 15895 21416 15904
rect 21364 15861 21373 15895
rect 21373 15861 21407 15895
rect 21407 15861 21416 15895
rect 21364 15852 21416 15861
rect 22652 15895 22704 15904
rect 22652 15861 22661 15895
rect 22661 15861 22695 15895
rect 22695 15861 22704 15895
rect 22652 15852 22704 15861
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 28632 15895 28684 15904
rect 28632 15861 28641 15895
rect 28641 15861 28675 15895
rect 28675 15861 28684 15895
rect 28632 15852 28684 15861
rect 29092 15895 29144 15904
rect 29092 15861 29101 15895
rect 29101 15861 29135 15895
rect 29135 15861 29144 15895
rect 29092 15852 29144 15861
rect 30380 15852 30432 15904
rect 32036 15895 32088 15904
rect 32036 15861 32045 15895
rect 32045 15861 32079 15895
rect 32079 15861 32088 15895
rect 32036 15852 32088 15861
rect 32220 15852 32272 15904
rect 33784 15852 33836 15904
rect 36912 15997 36921 16031
rect 36921 15997 36955 16031
rect 36955 15997 36964 16031
rect 36912 15988 36964 15997
rect 37924 16031 37976 16040
rect 37924 15997 37933 16031
rect 37933 15997 37967 16031
rect 37967 15997 37976 16031
rect 37924 15988 37976 15997
rect 42156 16031 42208 16040
rect 42156 15997 42165 16031
rect 42165 15997 42199 16031
rect 42199 15997 42208 16031
rect 42156 15988 42208 15997
rect 44272 16031 44324 16040
rect 44272 15997 44281 16031
rect 44281 15997 44315 16031
rect 44315 15997 44324 16031
rect 44272 15988 44324 15997
rect 46388 16031 46440 16040
rect 46388 15997 46397 16031
rect 46397 15997 46431 16031
rect 46431 15997 46440 16031
rect 46388 15988 46440 15997
rect 37832 15920 37884 15972
rect 40224 15920 40276 15972
rect 43536 15920 43588 15972
rect 46112 15963 46164 15972
rect 46112 15929 46121 15963
rect 46121 15929 46155 15963
rect 46155 15929 46164 15963
rect 46112 15920 46164 15929
rect 34704 15895 34756 15904
rect 34704 15861 34713 15895
rect 34713 15861 34747 15895
rect 34747 15861 34756 15895
rect 34704 15852 34756 15861
rect 38016 15852 38068 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 18512 15512 18564 15564
rect 20720 15580 20772 15632
rect 21364 15580 21416 15632
rect 21732 15623 21784 15632
rect 21732 15589 21741 15623
rect 21741 15589 21775 15623
rect 21775 15589 21784 15623
rect 21732 15580 21784 15589
rect 22652 15512 22704 15564
rect 26424 15648 26476 15700
rect 25228 15580 25280 15632
rect 25872 15580 25924 15632
rect 28356 15648 28408 15700
rect 29460 15648 29512 15700
rect 31668 15648 31720 15700
rect 32220 15648 32272 15700
rect 28632 15580 28684 15632
rect 24216 15555 24268 15564
rect 24216 15521 24225 15555
rect 24225 15521 24259 15555
rect 24259 15521 24268 15555
rect 24216 15512 24268 15521
rect 24860 15512 24912 15564
rect 29368 15555 29420 15564
rect 18972 15444 19024 15496
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 27068 15487 27120 15496
rect 23388 15444 23440 15453
rect 27068 15453 27077 15487
rect 27077 15453 27111 15487
rect 27111 15453 27120 15487
rect 27068 15444 27120 15453
rect 28724 15444 28776 15496
rect 29368 15521 29377 15555
rect 29377 15521 29411 15555
rect 29411 15521 29420 15555
rect 29368 15512 29420 15521
rect 32036 15580 32088 15632
rect 31576 15555 31628 15564
rect 31576 15521 31585 15555
rect 31585 15521 31619 15555
rect 31619 15521 31628 15555
rect 32404 15648 32456 15700
rect 34336 15648 34388 15700
rect 34428 15648 34480 15700
rect 35440 15648 35492 15700
rect 36912 15691 36964 15700
rect 36912 15657 36921 15691
rect 36921 15657 36955 15691
rect 36955 15657 36964 15691
rect 36912 15648 36964 15657
rect 37832 15648 37884 15700
rect 37924 15648 37976 15700
rect 41144 15691 41196 15700
rect 41144 15657 41153 15691
rect 41153 15657 41187 15691
rect 41187 15657 41196 15691
rect 41144 15648 41196 15657
rect 44272 15648 44324 15700
rect 33508 15580 33560 15632
rect 35532 15580 35584 15632
rect 32772 15555 32824 15564
rect 31576 15512 31628 15521
rect 32772 15521 32781 15555
rect 32781 15521 32815 15555
rect 32815 15521 32824 15555
rect 32772 15512 32824 15521
rect 33968 15512 34020 15564
rect 34336 15512 34388 15564
rect 35440 15512 35492 15564
rect 36452 15555 36504 15564
rect 36452 15521 36461 15555
rect 36461 15521 36495 15555
rect 36495 15521 36504 15555
rect 36452 15512 36504 15521
rect 37740 15555 37792 15564
rect 37740 15521 37749 15555
rect 37749 15521 37783 15555
rect 37783 15521 37792 15555
rect 37740 15512 37792 15521
rect 39948 15580 40000 15632
rect 42892 15580 42944 15632
rect 43536 15623 43588 15632
rect 43536 15589 43545 15623
rect 43545 15589 43579 15623
rect 43579 15589 43588 15623
rect 43536 15580 43588 15589
rect 46112 15580 46164 15632
rect 38292 15512 38344 15564
rect 42340 15512 42392 15564
rect 47308 15555 47360 15564
rect 47308 15521 47317 15555
rect 47317 15521 47351 15555
rect 47351 15521 47360 15555
rect 47308 15512 47360 15521
rect 29184 15444 29236 15496
rect 33784 15444 33836 15496
rect 34244 15444 34296 15496
rect 36544 15444 36596 15496
rect 39580 15444 39632 15496
rect 40316 15444 40368 15496
rect 40868 15444 40920 15496
rect 43444 15487 43496 15496
rect 43444 15453 43453 15487
rect 43453 15453 43487 15487
rect 43487 15453 43496 15487
rect 43444 15444 43496 15453
rect 45836 15487 45888 15496
rect 45836 15453 45845 15487
rect 45845 15453 45879 15487
rect 45879 15453 45888 15487
rect 45836 15444 45888 15453
rect 46480 15487 46532 15496
rect 46480 15453 46489 15487
rect 46489 15453 46523 15487
rect 46523 15453 46532 15487
rect 46480 15444 46532 15453
rect 21824 15376 21876 15428
rect 33140 15376 33192 15428
rect 34520 15376 34572 15428
rect 38476 15376 38528 15428
rect 43996 15419 44048 15428
rect 43996 15385 44005 15419
rect 44005 15385 44039 15419
rect 44039 15385 44048 15419
rect 43996 15376 44048 15385
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 33232 15351 33284 15360
rect 33232 15317 33241 15351
rect 33241 15317 33275 15351
rect 33275 15317 33284 15351
rect 33232 15308 33284 15317
rect 34336 15351 34388 15360
rect 34336 15317 34345 15351
rect 34345 15317 34379 15351
rect 34379 15317 34388 15351
rect 34336 15308 34388 15317
rect 35256 15308 35308 15360
rect 36820 15308 36872 15360
rect 42248 15308 42300 15360
rect 46204 15308 46256 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 18144 15104 18196 15156
rect 18512 15104 18564 15156
rect 21088 15104 21140 15156
rect 22652 15104 22704 15156
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 25872 15147 25924 15156
rect 25872 15113 25881 15147
rect 25881 15113 25915 15147
rect 25915 15113 25924 15147
rect 25872 15104 25924 15113
rect 26148 15147 26200 15156
rect 26148 15113 26157 15147
rect 26157 15113 26191 15147
rect 26191 15113 26200 15147
rect 26148 15104 26200 15113
rect 28264 15104 28316 15156
rect 32036 15104 32088 15156
rect 33784 15104 33836 15156
rect 34244 15104 34296 15156
rect 34428 15104 34480 15156
rect 35532 15104 35584 15156
rect 36544 15104 36596 15156
rect 38292 15147 38344 15156
rect 38292 15113 38301 15147
rect 38301 15113 38335 15147
rect 38335 15113 38344 15147
rect 38292 15104 38344 15113
rect 39580 15147 39632 15156
rect 39580 15113 39589 15147
rect 39589 15113 39623 15147
rect 39623 15113 39632 15147
rect 39580 15104 39632 15113
rect 40224 15147 40276 15156
rect 40224 15113 40233 15147
rect 40233 15113 40267 15147
rect 40267 15113 40276 15147
rect 40224 15104 40276 15113
rect 42340 15104 42392 15156
rect 42892 15147 42944 15156
rect 42892 15113 42901 15147
rect 42901 15113 42935 15147
rect 42935 15113 42944 15147
rect 42892 15104 42944 15113
rect 46112 15104 46164 15156
rect 47308 15147 47360 15156
rect 47308 15113 47317 15147
rect 47317 15113 47351 15147
rect 47351 15113 47360 15147
rect 47308 15104 47360 15113
rect 19156 15036 19208 15088
rect 19064 14900 19116 14952
rect 23480 15036 23532 15088
rect 24216 15036 24268 15088
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 22008 14968 22060 15020
rect 23756 15011 23808 15020
rect 17592 14807 17644 14816
rect 17592 14773 17601 14807
rect 17601 14773 17635 14807
rect 17635 14773 17644 14807
rect 17592 14764 17644 14773
rect 21916 14943 21968 14952
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 23756 14977 23765 15011
rect 23765 14977 23799 15011
rect 23799 14977 23808 15011
rect 25504 15036 25556 15088
rect 28724 15079 28776 15088
rect 28724 15045 28733 15079
rect 28733 15045 28767 15079
rect 28767 15045 28776 15079
rect 28724 15036 28776 15045
rect 29092 15079 29144 15088
rect 29092 15045 29101 15079
rect 29101 15045 29135 15079
rect 29135 15045 29144 15079
rect 29092 15036 29144 15045
rect 29460 15036 29512 15088
rect 33508 15079 33560 15088
rect 33508 15045 33517 15079
rect 33517 15045 33551 15079
rect 33551 15045 33560 15079
rect 33508 15036 33560 15045
rect 34520 15036 34572 15088
rect 34980 15036 35032 15088
rect 38108 15036 38160 15088
rect 23756 14968 23808 14977
rect 24768 14900 24820 14952
rect 25228 14943 25280 14952
rect 25228 14909 25272 14943
rect 25272 14909 25280 14943
rect 25228 14900 25280 14909
rect 20628 14832 20680 14884
rect 23388 14832 23440 14884
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 24400 14875 24452 14884
rect 24400 14841 24409 14875
rect 24409 14841 24443 14875
rect 24443 14841 24452 14875
rect 24400 14832 24452 14841
rect 24584 14832 24636 14884
rect 24860 14832 24912 14884
rect 29368 14968 29420 15020
rect 26516 14900 26568 14952
rect 28264 14900 28316 14952
rect 29276 14943 29328 14952
rect 29276 14909 29285 14943
rect 29285 14909 29319 14943
rect 29319 14909 29328 14943
rect 29276 14900 29328 14909
rect 31484 14900 31536 14952
rect 33232 14968 33284 15020
rect 35256 15011 35308 15020
rect 35256 14977 35265 15011
rect 35265 14977 35299 15011
rect 35299 14977 35308 15011
rect 35256 14968 35308 14977
rect 32772 14943 32824 14952
rect 32772 14909 32781 14943
rect 32781 14909 32815 14943
rect 32815 14909 32824 14943
rect 32772 14900 32824 14909
rect 26148 14832 26200 14884
rect 29460 14832 29512 14884
rect 34428 14900 34480 14952
rect 34612 14900 34664 14952
rect 35440 14900 35492 14952
rect 36912 14943 36964 14952
rect 36912 14909 36921 14943
rect 36921 14909 36955 14943
rect 36955 14909 36964 14943
rect 36912 14900 36964 14909
rect 37280 14900 37332 14952
rect 38292 14900 38344 14952
rect 38476 14943 38528 14952
rect 38476 14909 38485 14943
rect 38485 14909 38519 14943
rect 38519 14909 38528 14943
rect 40040 15036 40092 15088
rect 43536 15036 43588 15088
rect 43996 15079 44048 15088
rect 43996 15045 44005 15079
rect 44005 15045 44039 15079
rect 44039 15045 44048 15079
rect 43996 15036 44048 15045
rect 40592 15011 40644 15020
rect 40592 14977 40601 15011
rect 40601 14977 40635 15011
rect 40635 14977 40644 15011
rect 40592 14968 40644 14977
rect 40868 15011 40920 15020
rect 40868 14977 40877 15011
rect 40877 14977 40911 15011
rect 40911 14977 40920 15011
rect 40868 14968 40920 14977
rect 38476 14900 38528 14909
rect 41972 14900 42024 14952
rect 46204 15011 46256 15020
rect 46204 14977 46213 15011
rect 46213 14977 46247 15011
rect 46247 14977 46256 15011
rect 46204 14968 46256 14977
rect 46480 15011 46532 15020
rect 46480 14977 46489 15011
rect 46489 14977 46523 15011
rect 46523 14977 46532 15011
rect 46480 14968 46532 14977
rect 33968 14875 34020 14884
rect 33968 14841 33977 14875
rect 33977 14841 34011 14875
rect 34011 14841 34020 14875
rect 33968 14832 34020 14841
rect 35164 14832 35216 14884
rect 35624 14875 35676 14884
rect 35624 14841 35633 14875
rect 35633 14841 35667 14875
rect 35667 14841 35676 14875
rect 35624 14832 35676 14841
rect 37832 14832 37884 14884
rect 40224 14832 40276 14884
rect 41696 14832 41748 14884
rect 28540 14764 28592 14816
rect 30288 14764 30340 14816
rect 32404 14807 32456 14816
rect 32404 14773 32413 14807
rect 32413 14773 32447 14807
rect 32447 14773 32456 14807
rect 32404 14764 32456 14773
rect 36820 14764 36872 14816
rect 37740 14764 37792 14816
rect 39948 14807 40000 14816
rect 39948 14773 39957 14807
rect 39957 14773 39991 14807
rect 39991 14773 40000 14807
rect 42248 14832 42300 14884
rect 43536 14875 43588 14884
rect 43536 14841 43545 14875
rect 43545 14841 43579 14875
rect 43579 14841 43588 14875
rect 43536 14832 43588 14841
rect 46296 14875 46348 14884
rect 46296 14841 46305 14875
rect 46305 14841 46339 14875
rect 46339 14841 46348 14875
rect 46296 14832 46348 14841
rect 39948 14764 40000 14773
rect 41880 14764 41932 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 21180 14560 21232 14612
rect 23572 14560 23624 14612
rect 25228 14560 25280 14612
rect 30564 14603 30616 14612
rect 30564 14569 30573 14603
rect 30573 14569 30607 14603
rect 30607 14569 30616 14603
rect 30564 14560 30616 14569
rect 33784 14603 33836 14612
rect 33784 14569 33793 14603
rect 33793 14569 33827 14603
rect 33827 14569 33836 14603
rect 33784 14560 33836 14569
rect 33968 14560 34020 14612
rect 35532 14603 35584 14612
rect 35532 14569 35541 14603
rect 35541 14569 35575 14603
rect 35575 14569 35584 14603
rect 35532 14560 35584 14569
rect 36452 14603 36504 14612
rect 36452 14569 36461 14603
rect 36461 14569 36495 14603
rect 36495 14569 36504 14603
rect 36452 14560 36504 14569
rect 40592 14603 40644 14612
rect 18696 14492 18748 14544
rect 19892 14492 19944 14544
rect 20812 14492 20864 14544
rect 21732 14492 21784 14544
rect 23296 14492 23348 14544
rect 24952 14535 25004 14544
rect 24952 14501 24961 14535
rect 24961 14501 24995 14535
rect 24995 14501 25004 14535
rect 24952 14492 25004 14501
rect 26700 14492 26752 14544
rect 26792 14492 26844 14544
rect 29276 14492 29328 14544
rect 32864 14535 32916 14544
rect 32864 14501 32873 14535
rect 32873 14501 32907 14535
rect 32907 14501 32916 14535
rect 32864 14492 32916 14501
rect 19248 14424 19300 14476
rect 28724 14467 28776 14476
rect 28724 14433 28733 14467
rect 28733 14433 28767 14467
rect 28767 14433 28776 14467
rect 28724 14424 28776 14433
rect 29368 14424 29420 14476
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 24400 14356 24452 14408
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 26424 14356 26476 14408
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27344 14399 27396 14408
rect 27344 14365 27353 14399
rect 27353 14365 27387 14399
rect 27387 14365 27396 14399
rect 27344 14356 27396 14365
rect 30104 14356 30156 14408
rect 31760 14424 31812 14476
rect 33508 14492 33560 14544
rect 35256 14492 35308 14544
rect 38016 14492 38068 14544
rect 39948 14492 40000 14544
rect 40592 14569 40601 14603
rect 40601 14569 40635 14603
rect 40635 14569 40644 14603
rect 40592 14560 40644 14569
rect 41972 14492 42024 14544
rect 33140 14356 33192 14408
rect 33416 14399 33468 14408
rect 33416 14365 33425 14399
rect 33425 14365 33459 14399
rect 33459 14365 33468 14399
rect 33416 14356 33468 14365
rect 34612 14356 34664 14408
rect 35624 14424 35676 14476
rect 36268 14424 36320 14476
rect 40776 14424 40828 14476
rect 41604 14424 41656 14476
rect 42064 14424 42116 14476
rect 35164 14356 35216 14408
rect 37832 14399 37884 14408
rect 37832 14365 37841 14399
rect 37841 14365 37875 14399
rect 37875 14365 37884 14399
rect 37832 14356 37884 14365
rect 39672 14399 39724 14408
rect 39672 14365 39681 14399
rect 39681 14365 39715 14399
rect 39715 14365 39724 14399
rect 39672 14356 39724 14365
rect 43444 14560 43496 14612
rect 43536 14560 43588 14612
rect 46296 14560 46348 14612
rect 43996 14492 44048 14544
rect 45192 14535 45244 14544
rect 45192 14501 45201 14535
rect 45201 14501 45235 14535
rect 45235 14501 45244 14535
rect 45192 14492 45244 14501
rect 45560 14492 45612 14544
rect 45836 14535 45888 14544
rect 45836 14501 45845 14535
rect 45845 14501 45879 14535
rect 45879 14501 45888 14535
rect 45836 14492 45888 14501
rect 43720 14467 43772 14476
rect 43720 14433 43729 14467
rect 43729 14433 43763 14467
rect 43763 14433 43772 14467
rect 43720 14424 43772 14433
rect 46020 14424 46072 14476
rect 46848 14424 46900 14476
rect 19432 14288 19484 14340
rect 34336 14288 34388 14340
rect 28264 14263 28316 14272
rect 28264 14229 28273 14263
rect 28273 14229 28307 14263
rect 28307 14229 28316 14263
rect 28264 14220 28316 14229
rect 35808 14220 35860 14272
rect 36360 14220 36412 14272
rect 36912 14263 36964 14272
rect 36912 14229 36921 14263
rect 36921 14229 36955 14263
rect 36955 14229 36964 14263
rect 36912 14220 36964 14229
rect 41420 14220 41472 14272
rect 41604 14263 41656 14272
rect 41604 14229 41613 14263
rect 41613 14229 41647 14263
rect 41647 14229 41656 14263
rect 41604 14220 41656 14229
rect 42432 14220 42484 14272
rect 46940 14220 46992 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 17592 14016 17644 14068
rect 20812 14016 20864 14068
rect 23204 14059 23256 14068
rect 23204 14025 23213 14059
rect 23213 14025 23247 14059
rect 23247 14025 23256 14059
rect 23204 14016 23256 14025
rect 23296 14016 23348 14068
rect 24860 14016 24912 14068
rect 26792 14016 26844 14068
rect 30104 14059 30156 14068
rect 20628 13948 20680 14000
rect 24308 13991 24360 14000
rect 19064 13880 19116 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 24308 13957 24317 13991
rect 24317 13957 24351 13991
rect 24351 13957 24360 13991
rect 24308 13948 24360 13957
rect 24952 13948 25004 14000
rect 29276 13948 29328 14000
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 31484 14059 31536 14068
rect 31484 14025 31493 14059
rect 31493 14025 31527 14059
rect 31527 14025 31536 14059
rect 31484 14016 31536 14025
rect 31760 14059 31812 14068
rect 31760 14025 31769 14059
rect 31769 14025 31803 14059
rect 31803 14025 31812 14059
rect 31760 14016 31812 14025
rect 32864 14016 32916 14068
rect 34612 14059 34664 14068
rect 34612 14025 34621 14059
rect 34621 14025 34655 14059
rect 34655 14025 34664 14059
rect 34612 14016 34664 14025
rect 34704 14016 34756 14068
rect 36268 14059 36320 14068
rect 36268 14025 36277 14059
rect 36277 14025 36311 14059
rect 36311 14025 36320 14059
rect 36268 14016 36320 14025
rect 37832 14016 37884 14068
rect 39672 14016 39724 14068
rect 43720 14016 43772 14068
rect 45192 14016 45244 14068
rect 46848 14059 46900 14068
rect 46848 14025 46857 14059
rect 46857 14025 46891 14059
rect 46891 14025 46900 14059
rect 46848 14016 46900 14025
rect 35440 13948 35492 14000
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 19340 13812 19392 13864
rect 25780 13880 25832 13932
rect 27068 13880 27120 13932
rect 27344 13923 27396 13932
rect 27344 13889 27353 13923
rect 27353 13889 27387 13923
rect 27387 13889 27396 13923
rect 27344 13880 27396 13889
rect 30564 13923 30616 13932
rect 30564 13889 30573 13923
rect 30573 13889 30607 13923
rect 30607 13889 30616 13923
rect 30564 13880 30616 13889
rect 35256 13923 35308 13932
rect 29368 13812 29420 13864
rect 16212 13744 16264 13796
rect 17960 13744 18012 13796
rect 18788 13744 18840 13796
rect 22192 13787 22244 13796
rect 22192 13753 22195 13787
rect 22195 13753 22229 13787
rect 22229 13753 22244 13787
rect 24492 13787 24544 13796
rect 22192 13744 22244 13753
rect 24492 13753 24501 13787
rect 24501 13753 24535 13787
rect 24535 13753 24544 13787
rect 24492 13744 24544 13753
rect 17040 13676 17092 13728
rect 20904 13676 20956 13728
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 24308 13676 24360 13728
rect 27068 13744 27120 13796
rect 28724 13787 28776 13796
rect 28724 13753 28733 13787
rect 28733 13753 28767 13787
rect 28767 13753 28776 13787
rect 31944 13812 31996 13864
rect 32404 13812 32456 13864
rect 32772 13812 32824 13864
rect 33416 13812 33468 13864
rect 28724 13744 28776 13753
rect 27804 13719 27856 13728
rect 27804 13685 27813 13719
rect 27813 13685 27847 13719
rect 27847 13685 27856 13719
rect 27804 13676 27856 13685
rect 28540 13676 28592 13728
rect 29460 13676 29512 13728
rect 34520 13744 34572 13796
rect 35256 13889 35265 13923
rect 35265 13889 35299 13923
rect 35299 13889 35308 13923
rect 35256 13880 35308 13889
rect 37188 13880 37240 13932
rect 38016 13880 38068 13932
rect 39948 13880 40000 13932
rect 37004 13855 37056 13864
rect 37004 13821 37013 13855
rect 37013 13821 37047 13855
rect 37047 13821 37056 13855
rect 37004 13812 37056 13821
rect 42892 13948 42944 14000
rect 43812 13948 43864 14000
rect 41420 13880 41472 13932
rect 46848 13812 46900 13864
rect 42340 13787 42392 13796
rect 32404 13676 32456 13728
rect 33876 13719 33928 13728
rect 33876 13685 33885 13719
rect 33885 13685 33919 13719
rect 33919 13685 33928 13719
rect 33876 13676 33928 13685
rect 37188 13676 37240 13728
rect 38936 13719 38988 13728
rect 38936 13685 38945 13719
rect 38945 13685 38979 13719
rect 38979 13685 38988 13719
rect 38936 13676 38988 13685
rect 41696 13676 41748 13728
rect 42340 13753 42349 13787
rect 42349 13753 42383 13787
rect 42383 13753 42392 13787
rect 42340 13744 42392 13753
rect 41972 13676 42024 13728
rect 42064 13676 42116 13728
rect 43812 13787 43864 13796
rect 43812 13753 43821 13787
rect 43821 13753 43855 13787
rect 43855 13753 43864 13787
rect 44364 13787 44416 13796
rect 43812 13744 43864 13753
rect 44364 13753 44373 13787
rect 44373 13753 44407 13787
rect 44407 13753 44416 13787
rect 44364 13744 44416 13753
rect 45468 13676 45520 13728
rect 46572 13719 46624 13728
rect 46572 13685 46581 13719
rect 46581 13685 46615 13719
rect 46615 13685 46624 13719
rect 46572 13676 46624 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 20996 13472 21048 13524
rect 24492 13515 24544 13524
rect 24492 13481 24501 13515
rect 24501 13481 24535 13515
rect 24535 13481 24544 13515
rect 24492 13472 24544 13481
rect 17132 13404 17184 13456
rect 22192 13404 22244 13456
rect 22836 13404 22888 13456
rect 25136 13472 25188 13524
rect 25780 13404 25832 13456
rect 29368 13472 29420 13524
rect 30564 13472 30616 13524
rect 33416 13472 33468 13524
rect 34520 13515 34572 13524
rect 34520 13481 34529 13515
rect 34529 13481 34563 13515
rect 34563 13481 34572 13515
rect 34520 13472 34572 13481
rect 35256 13472 35308 13524
rect 41512 13472 41564 13524
rect 26792 13404 26844 13456
rect 28540 13404 28592 13456
rect 30104 13404 30156 13456
rect 30380 13447 30432 13456
rect 30380 13413 30389 13447
rect 30389 13413 30423 13447
rect 30423 13413 30432 13447
rect 30380 13404 30432 13413
rect 32864 13404 32916 13456
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 20904 13336 20956 13388
rect 24768 13336 24820 13388
rect 28264 13336 28316 13388
rect 32772 13379 32824 13388
rect 32772 13345 32781 13379
rect 32781 13345 32815 13379
rect 32815 13345 32824 13379
rect 32772 13336 32824 13345
rect 34704 13336 34756 13388
rect 34796 13379 34848 13388
rect 34796 13345 34805 13379
rect 34805 13345 34839 13379
rect 34839 13345 34848 13379
rect 35992 13379 36044 13388
rect 34796 13336 34848 13345
rect 35992 13345 36001 13379
rect 36001 13345 36035 13379
rect 36035 13345 36044 13379
rect 35992 13336 36044 13345
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 16948 13268 17000 13320
rect 20996 13268 21048 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 26608 13311 26660 13320
rect 26608 13277 26617 13311
rect 26617 13277 26651 13311
rect 26651 13277 26660 13311
rect 26608 13268 26660 13277
rect 26700 13268 26752 13320
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 30288 13311 30340 13320
rect 30288 13277 30297 13311
rect 30297 13277 30331 13311
rect 30331 13277 30340 13311
rect 30288 13268 30340 13277
rect 30656 13268 30708 13320
rect 32588 13268 32640 13320
rect 36176 13268 36228 13320
rect 37004 13447 37056 13456
rect 37004 13413 37013 13447
rect 37013 13413 37047 13447
rect 37047 13413 37056 13447
rect 37004 13404 37056 13413
rect 37280 13336 37332 13388
rect 37924 13379 37976 13388
rect 37924 13345 37933 13379
rect 37933 13345 37967 13379
rect 37967 13345 37976 13379
rect 37924 13336 37976 13345
rect 39120 13404 39172 13456
rect 40960 13404 41012 13456
rect 43444 13404 43496 13456
rect 45376 13447 45428 13456
rect 45376 13413 45385 13447
rect 45385 13413 45419 13447
rect 45419 13413 45428 13447
rect 45376 13404 45428 13413
rect 45468 13404 45520 13456
rect 39856 13336 39908 13388
rect 42616 13336 42668 13388
rect 46940 13336 46992 13388
rect 47124 13379 47176 13388
rect 47124 13345 47133 13379
rect 47133 13345 47167 13379
rect 47167 13345 47176 13379
rect 47124 13336 47176 13345
rect 38660 13311 38712 13320
rect 38660 13277 38669 13311
rect 38669 13277 38703 13311
rect 38703 13277 38712 13311
rect 38660 13268 38712 13277
rect 40316 13268 40368 13320
rect 43720 13311 43772 13320
rect 43720 13277 43729 13311
rect 43729 13277 43763 13311
rect 43763 13277 43772 13311
rect 43720 13268 43772 13277
rect 44364 13311 44416 13320
rect 44364 13277 44373 13311
rect 44373 13277 44407 13311
rect 44407 13277 44416 13311
rect 45284 13311 45336 13320
rect 44364 13268 44416 13277
rect 45284 13277 45293 13311
rect 45293 13277 45327 13311
rect 45327 13277 45336 13311
rect 45284 13268 45336 13277
rect 27804 13200 27856 13252
rect 30748 13200 30800 13252
rect 45836 13243 45888 13252
rect 45836 13209 45845 13243
rect 45845 13209 45879 13243
rect 45879 13209 45888 13243
rect 45836 13200 45888 13209
rect 17132 13132 17184 13184
rect 18788 13132 18840 13184
rect 22008 13132 22060 13184
rect 27068 13132 27120 13184
rect 28080 13132 28132 13184
rect 29276 13132 29328 13184
rect 33508 13175 33560 13184
rect 33508 13141 33517 13175
rect 33517 13141 33551 13175
rect 33551 13141 33560 13175
rect 33508 13132 33560 13141
rect 39672 13175 39724 13184
rect 39672 13141 39681 13175
rect 39681 13141 39715 13175
rect 39715 13141 39724 13175
rect 39672 13132 39724 13141
rect 40960 13132 41012 13184
rect 42156 13175 42208 13184
rect 42156 13141 42165 13175
rect 42165 13141 42199 13175
rect 42199 13141 42208 13175
rect 42156 13132 42208 13141
rect 43536 13132 43588 13184
rect 46296 13175 46348 13184
rect 46296 13141 46305 13175
rect 46305 13141 46339 13175
rect 46339 13141 46348 13175
rect 46296 13132 46348 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 16120 12928 16172 12980
rect 17868 12928 17920 12980
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 22836 12971 22888 12980
rect 22836 12937 22845 12971
rect 22845 12937 22879 12971
rect 22879 12937 22888 12971
rect 22836 12928 22888 12937
rect 24584 12971 24636 12980
rect 24584 12937 24593 12971
rect 24593 12937 24627 12971
rect 24627 12937 24636 12971
rect 24584 12928 24636 12937
rect 25136 12971 25188 12980
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 26792 12928 26844 12980
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 27068 12860 27120 12912
rect 30012 12860 30064 12912
rect 22192 12792 22244 12844
rect 23296 12792 23348 12844
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 17132 12656 17184 12708
rect 19248 12656 19300 12708
rect 19340 12656 19392 12708
rect 22008 12656 22060 12708
rect 22744 12724 22796 12776
rect 24584 12724 24636 12776
rect 25688 12724 25740 12776
rect 26332 12792 26384 12844
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 28632 12792 28684 12844
rect 29368 12835 29420 12844
rect 29368 12801 29377 12835
rect 29377 12801 29411 12835
rect 29411 12801 29420 12835
rect 29368 12792 29420 12801
rect 27896 12767 27948 12776
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 17960 12588 18012 12640
rect 18512 12588 18564 12640
rect 26056 12656 26108 12708
rect 27896 12733 27905 12767
rect 27905 12733 27939 12767
rect 27939 12733 27948 12767
rect 27896 12724 27948 12733
rect 28080 12767 28132 12776
rect 28080 12733 28089 12767
rect 28089 12733 28123 12767
rect 28123 12733 28132 12767
rect 28080 12724 28132 12733
rect 37280 12971 37332 12980
rect 37280 12937 37289 12971
rect 37289 12937 37323 12971
rect 37323 12937 37332 12971
rect 37280 12928 37332 12937
rect 41604 12928 41656 12980
rect 43444 12928 43496 12980
rect 47124 12971 47176 12980
rect 47124 12937 47133 12971
rect 47133 12937 47167 12971
rect 47167 12937 47176 12971
rect 47124 12928 47176 12937
rect 32404 12860 32456 12912
rect 21088 12588 21140 12640
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 28540 12588 28592 12640
rect 28908 12588 28960 12640
rect 29092 12656 29144 12708
rect 30012 12699 30064 12708
rect 30012 12665 30021 12699
rect 30021 12665 30055 12699
rect 30055 12665 30064 12699
rect 30012 12656 30064 12665
rect 32864 12860 32916 12912
rect 35992 12860 36044 12912
rect 39856 12903 39908 12912
rect 39856 12869 39865 12903
rect 39865 12869 39899 12903
rect 39899 12869 39908 12903
rect 39856 12860 39908 12869
rect 40868 12860 40920 12912
rect 32956 12656 33008 12708
rect 33324 12767 33376 12776
rect 33324 12733 33333 12767
rect 33333 12733 33367 12767
rect 33367 12733 33376 12767
rect 33324 12724 33376 12733
rect 33508 12767 33560 12776
rect 33508 12733 33517 12767
rect 33517 12733 33551 12767
rect 33551 12733 33560 12767
rect 35348 12792 35400 12844
rect 33508 12724 33560 12733
rect 38108 12792 38160 12844
rect 38660 12835 38712 12844
rect 38660 12801 38669 12835
rect 38669 12801 38703 12835
rect 38703 12801 38712 12835
rect 38660 12792 38712 12801
rect 34796 12656 34848 12708
rect 36176 12724 36228 12776
rect 37280 12724 37332 12776
rect 38844 12724 38896 12776
rect 42156 12835 42208 12844
rect 42156 12801 42165 12835
rect 42165 12801 42199 12835
rect 42199 12801 42208 12835
rect 42156 12792 42208 12801
rect 42248 12792 42300 12844
rect 42524 12792 42576 12844
rect 43720 12792 43772 12844
rect 46020 12792 46072 12844
rect 46204 12792 46256 12844
rect 40960 12767 41012 12776
rect 40960 12733 40969 12767
rect 40969 12733 41003 12767
rect 41003 12733 41012 12767
rect 40960 12724 41012 12733
rect 36544 12656 36596 12708
rect 30104 12588 30156 12640
rect 30380 12588 30432 12640
rect 31300 12631 31352 12640
rect 31300 12597 31309 12631
rect 31309 12597 31343 12631
rect 31343 12597 31352 12631
rect 31300 12588 31352 12597
rect 32588 12588 32640 12640
rect 37556 12656 37608 12708
rect 37924 12699 37976 12708
rect 37924 12665 37933 12699
rect 37933 12665 37967 12699
rect 37967 12665 37976 12699
rect 37924 12656 37976 12665
rect 37648 12631 37700 12640
rect 37648 12597 37657 12631
rect 37657 12597 37691 12631
rect 37691 12597 37700 12631
rect 37648 12588 37700 12597
rect 38016 12588 38068 12640
rect 40316 12588 40368 12640
rect 41972 12631 42024 12640
rect 41972 12597 41981 12631
rect 41981 12597 42015 12631
rect 42015 12597 42024 12631
rect 41972 12588 42024 12597
rect 42524 12588 42576 12640
rect 43536 12656 43588 12708
rect 44456 12656 44508 12708
rect 46204 12699 46256 12708
rect 46204 12665 46213 12699
rect 46213 12665 46247 12699
rect 46247 12665 46256 12699
rect 46204 12656 46256 12665
rect 45376 12588 45428 12640
rect 46848 12656 46900 12708
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 17868 12384 17920 12436
rect 19340 12427 19392 12436
rect 19340 12393 19349 12427
rect 19349 12393 19383 12427
rect 19383 12393 19392 12427
rect 19340 12384 19392 12393
rect 22192 12427 22244 12436
rect 22192 12393 22201 12427
rect 22201 12393 22235 12427
rect 22235 12393 22244 12427
rect 22192 12384 22244 12393
rect 24768 12427 24820 12436
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 26056 12427 26108 12436
rect 26056 12393 26065 12427
rect 26065 12393 26099 12427
rect 26099 12393 26108 12427
rect 26056 12384 26108 12393
rect 26608 12384 26660 12436
rect 28356 12427 28408 12436
rect 28356 12393 28365 12427
rect 28365 12393 28399 12427
rect 28399 12393 28408 12427
rect 28356 12384 28408 12393
rect 29368 12427 29420 12436
rect 29368 12393 29377 12427
rect 29377 12393 29411 12427
rect 29411 12393 29420 12427
rect 29368 12384 29420 12393
rect 33324 12427 33376 12436
rect 33324 12393 33333 12427
rect 33333 12393 33367 12427
rect 33367 12393 33376 12427
rect 33324 12384 33376 12393
rect 34704 12427 34756 12436
rect 34704 12393 34713 12427
rect 34713 12393 34747 12427
rect 34747 12393 34756 12427
rect 34704 12384 34756 12393
rect 35348 12384 35400 12436
rect 36084 12384 36136 12436
rect 37280 12384 37332 12436
rect 40316 12427 40368 12436
rect 40316 12393 40325 12427
rect 40325 12393 40359 12427
rect 40359 12393 40368 12427
rect 40316 12384 40368 12393
rect 42064 12384 42116 12436
rect 42156 12384 42208 12436
rect 42616 12427 42668 12436
rect 42616 12393 42625 12427
rect 42625 12393 42659 12427
rect 42659 12393 42668 12427
rect 42616 12384 42668 12393
rect 43536 12384 43588 12436
rect 45284 12384 45336 12436
rect 21088 12359 21140 12368
rect 21088 12325 21097 12359
rect 21097 12325 21131 12359
rect 21131 12325 21140 12359
rect 21088 12316 21140 12325
rect 23204 12316 23256 12368
rect 26792 12316 26844 12368
rect 27804 12359 27856 12368
rect 27804 12325 27813 12359
rect 27813 12325 27847 12359
rect 27847 12325 27856 12359
rect 27804 12316 27856 12325
rect 28908 12316 28960 12368
rect 30748 12316 30800 12368
rect 32496 12359 32548 12368
rect 32496 12325 32505 12359
rect 32505 12325 32539 12359
rect 32539 12325 32548 12359
rect 32496 12316 32548 12325
rect 33692 12316 33744 12368
rect 38016 12316 38068 12368
rect 40868 12316 40920 12368
rect 45468 12359 45520 12368
rect 45468 12325 45477 12359
rect 45477 12325 45511 12359
rect 45511 12325 45520 12359
rect 45468 12316 45520 12325
rect 46020 12359 46072 12368
rect 46020 12325 46029 12359
rect 46029 12325 46063 12359
rect 46063 12325 46072 12359
rect 46020 12316 46072 12325
rect 46848 12359 46900 12368
rect 46848 12325 46857 12359
rect 46857 12325 46891 12359
rect 46891 12325 46900 12359
rect 46848 12316 46900 12325
rect 17408 12248 17460 12300
rect 18972 12291 19024 12300
rect 18972 12257 18981 12291
rect 18981 12257 19015 12291
rect 19015 12257 19024 12291
rect 18972 12248 19024 12257
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 24860 12248 24912 12300
rect 26240 12248 26292 12300
rect 28448 12248 28500 12300
rect 32588 12248 32640 12300
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 28172 12180 28224 12232
rect 29092 12180 29144 12232
rect 30380 12180 30432 12232
rect 24492 12112 24544 12164
rect 33876 12180 33928 12232
rect 34796 12248 34848 12300
rect 36084 12248 36136 12300
rect 36544 12248 36596 12300
rect 42156 12291 42208 12300
rect 42156 12257 42200 12291
rect 42200 12257 42208 12291
rect 42156 12248 42208 12257
rect 43260 12248 43312 12300
rect 46572 12248 46624 12300
rect 34428 12223 34480 12232
rect 34428 12189 34437 12223
rect 34437 12189 34471 12223
rect 34471 12189 34480 12223
rect 34428 12180 34480 12189
rect 37924 12180 37976 12232
rect 40592 12180 40644 12232
rect 43628 12180 43680 12232
rect 44732 12180 44784 12232
rect 45376 12223 45428 12232
rect 45376 12189 45385 12223
rect 45385 12189 45419 12223
rect 45419 12189 45428 12223
rect 45376 12180 45428 12189
rect 36452 12112 36504 12164
rect 36636 12112 36688 12164
rect 38844 12112 38896 12164
rect 19892 12087 19944 12096
rect 19892 12053 19901 12087
rect 19901 12053 19935 12087
rect 19935 12053 19944 12087
rect 19892 12044 19944 12053
rect 24676 12044 24728 12096
rect 24952 12044 25004 12096
rect 25320 12044 25372 12096
rect 35532 12087 35584 12096
rect 35532 12053 35541 12087
rect 35541 12053 35575 12087
rect 35575 12053 35584 12087
rect 35532 12044 35584 12053
rect 37648 12044 37700 12096
rect 39120 12087 39172 12096
rect 39120 12053 39129 12087
rect 39129 12053 39163 12087
rect 39163 12053 39172 12087
rect 39120 12044 39172 12053
rect 41788 12044 41840 12096
rect 43628 12044 43680 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 18972 11840 19024 11892
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 23204 11840 23256 11892
rect 23388 11883 23440 11892
rect 23388 11849 23397 11883
rect 23397 11849 23431 11883
rect 23431 11849 23440 11883
rect 23388 11840 23440 11849
rect 26240 11883 26292 11892
rect 26240 11849 26249 11883
rect 26249 11849 26283 11883
rect 26283 11849 26292 11883
rect 26240 11840 26292 11849
rect 26792 11840 26844 11892
rect 28172 11883 28224 11892
rect 28172 11849 28181 11883
rect 28181 11849 28215 11883
rect 28215 11849 28224 11883
rect 28172 11840 28224 11849
rect 29092 11883 29144 11892
rect 29092 11849 29101 11883
rect 29101 11849 29135 11883
rect 29135 11849 29144 11883
rect 29092 11840 29144 11849
rect 33692 11840 33744 11892
rect 36084 11883 36136 11892
rect 36084 11849 36093 11883
rect 36093 11849 36127 11883
rect 36127 11849 36136 11883
rect 36084 11840 36136 11849
rect 36544 11840 36596 11892
rect 40868 11840 40920 11892
rect 42248 11840 42300 11892
rect 43260 11883 43312 11892
rect 43260 11849 43269 11883
rect 43269 11849 43303 11883
rect 43303 11849 43312 11883
rect 43260 11840 43312 11849
rect 43444 11840 43496 11892
rect 45468 11840 45520 11892
rect 46572 11840 46624 11892
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 20628 11772 20680 11824
rect 23848 11704 23900 11756
rect 24492 11704 24544 11756
rect 24676 11704 24728 11756
rect 30012 11704 30064 11756
rect 37648 11704 37700 11756
rect 42432 11772 42484 11824
rect 20444 11679 20496 11688
rect 20444 11645 20462 11679
rect 20462 11645 20496 11679
rect 20444 11636 20496 11645
rect 21272 11636 21324 11688
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 22008 11636 22060 11688
rect 27620 11636 27672 11688
rect 28908 11636 28960 11688
rect 32588 11679 32640 11688
rect 32588 11645 32597 11679
rect 32597 11645 32631 11679
rect 32631 11645 32640 11679
rect 32588 11636 32640 11645
rect 33048 11636 33100 11688
rect 35532 11679 35584 11688
rect 23388 11568 23440 11620
rect 17408 11500 17460 11552
rect 19432 11500 19484 11552
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 21732 11500 21784 11509
rect 25320 11611 25372 11620
rect 25320 11577 25329 11611
rect 25329 11577 25363 11611
rect 25363 11577 25372 11611
rect 25320 11568 25372 11577
rect 24492 11500 24544 11552
rect 26700 11500 26752 11552
rect 26792 11500 26844 11552
rect 26976 11611 27028 11620
rect 26976 11577 26985 11611
rect 26985 11577 27019 11611
rect 27019 11577 27028 11611
rect 26976 11568 27028 11577
rect 29828 11568 29880 11620
rect 28448 11500 28500 11552
rect 30104 11611 30156 11620
rect 30104 11577 30113 11611
rect 30113 11577 30147 11611
rect 30147 11577 30156 11611
rect 31576 11611 31628 11620
rect 30104 11568 30156 11577
rect 31576 11577 31585 11611
rect 31585 11577 31619 11611
rect 31619 11577 31628 11611
rect 31576 11568 31628 11577
rect 32680 11568 32732 11620
rect 33324 11568 33376 11620
rect 33508 11611 33560 11620
rect 33508 11577 33517 11611
rect 33517 11577 33551 11611
rect 33551 11577 33560 11611
rect 33508 11568 33560 11577
rect 30840 11500 30892 11552
rect 35532 11645 35541 11679
rect 35541 11645 35575 11679
rect 35575 11645 35584 11679
rect 35532 11636 35584 11645
rect 36728 11636 36780 11688
rect 35716 11611 35768 11620
rect 35716 11577 35725 11611
rect 35725 11577 35759 11611
rect 35759 11577 35768 11611
rect 35716 11568 35768 11577
rect 35900 11500 35952 11552
rect 37924 11611 37976 11620
rect 37924 11577 37933 11611
rect 37933 11577 37967 11611
rect 37967 11577 37976 11611
rect 37924 11568 37976 11577
rect 37832 11500 37884 11552
rect 38016 11500 38068 11552
rect 38568 11500 38620 11552
rect 38936 11636 38988 11688
rect 39120 11636 39172 11688
rect 42340 11704 42392 11756
rect 40500 11679 40552 11688
rect 40500 11645 40509 11679
rect 40509 11645 40543 11679
rect 40543 11645 40552 11679
rect 40500 11636 40552 11645
rect 40960 11679 41012 11688
rect 40960 11645 40969 11679
rect 40969 11645 41003 11679
rect 41003 11645 41012 11679
rect 40960 11636 41012 11645
rect 39580 11611 39632 11620
rect 39580 11577 39589 11611
rect 39589 11577 39623 11611
rect 39623 11577 39632 11611
rect 39580 11568 39632 11577
rect 42248 11568 42300 11620
rect 43628 11568 43680 11620
rect 44456 11611 44508 11620
rect 40592 11543 40644 11552
rect 40592 11509 40601 11543
rect 40601 11509 40635 11543
rect 40635 11509 40644 11543
rect 40592 11500 40644 11509
rect 42064 11500 42116 11552
rect 43260 11500 43312 11552
rect 43444 11500 43496 11552
rect 44456 11577 44465 11611
rect 44465 11577 44499 11611
rect 44499 11577 44508 11611
rect 44456 11568 44508 11577
rect 44548 11568 44600 11620
rect 45376 11568 45428 11620
rect 43996 11500 44048 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 18604 11339 18656 11348
rect 18604 11305 18613 11339
rect 18613 11305 18647 11339
rect 18647 11305 18656 11339
rect 18604 11296 18656 11305
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 21088 11296 21140 11348
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 28724 11339 28776 11348
rect 28724 11305 28733 11339
rect 28733 11305 28767 11339
rect 28767 11305 28776 11339
rect 28724 11296 28776 11305
rect 29828 11296 29880 11348
rect 30104 11296 30156 11348
rect 31576 11339 31628 11348
rect 31576 11305 31585 11339
rect 31585 11305 31619 11339
rect 31619 11305 31628 11339
rect 31576 11296 31628 11305
rect 32496 11339 32548 11348
rect 32496 11305 32505 11339
rect 32505 11305 32539 11339
rect 32539 11305 32548 11339
rect 32496 11296 32548 11305
rect 19156 11228 19208 11280
rect 19892 11228 19944 11280
rect 17868 11160 17920 11212
rect 20076 11160 20128 11212
rect 20628 11228 20680 11280
rect 21272 11228 21324 11280
rect 26700 11228 26752 11280
rect 27620 11228 27672 11280
rect 27804 11271 27856 11280
rect 27804 11237 27813 11271
rect 27813 11237 27847 11271
rect 27847 11237 27856 11271
rect 27804 11228 27856 11237
rect 33600 11296 33652 11348
rect 33876 11339 33928 11348
rect 33876 11305 33885 11339
rect 33885 11305 33919 11339
rect 33919 11305 33928 11339
rect 33876 11296 33928 11305
rect 36728 11339 36780 11348
rect 36728 11305 36737 11339
rect 36737 11305 36771 11339
rect 36771 11305 36780 11339
rect 36728 11296 36780 11305
rect 37648 11296 37700 11348
rect 37924 11339 37976 11348
rect 37924 11305 37933 11339
rect 37933 11305 37967 11339
rect 37967 11305 37976 11339
rect 37924 11296 37976 11305
rect 40592 11296 40644 11348
rect 42156 11339 42208 11348
rect 42156 11305 42165 11339
rect 42165 11305 42199 11339
rect 42199 11305 42208 11339
rect 42156 11296 42208 11305
rect 38752 11271 38804 11280
rect 20996 11160 21048 11212
rect 23388 11203 23440 11212
rect 23388 11169 23432 11203
rect 23432 11169 23440 11203
rect 28632 11203 28684 11212
rect 23388 11160 23440 11169
rect 28632 11169 28641 11203
rect 28641 11169 28675 11203
rect 28675 11169 28684 11203
rect 28632 11160 28684 11169
rect 29276 11160 29328 11212
rect 30472 11203 30524 11212
rect 30472 11169 30481 11203
rect 30481 11169 30515 11203
rect 30515 11169 30524 11203
rect 30472 11160 30524 11169
rect 18972 11092 19024 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 27436 11092 27488 11144
rect 30012 11092 30064 11144
rect 33876 11160 33928 11212
rect 34612 11160 34664 11212
rect 35532 11203 35584 11212
rect 35532 11169 35541 11203
rect 35541 11169 35575 11203
rect 35575 11169 35584 11203
rect 35532 11160 35584 11169
rect 38752 11237 38761 11271
rect 38761 11237 38795 11271
rect 38795 11237 38804 11271
rect 38752 11228 38804 11237
rect 40868 11228 40920 11280
rect 43996 11271 44048 11280
rect 43996 11237 44005 11271
rect 44005 11237 44039 11271
rect 44039 11237 44048 11271
rect 43996 11228 44048 11237
rect 37280 11160 37332 11212
rect 45192 11160 45244 11212
rect 30932 11135 30984 11144
rect 30932 11101 30941 11135
rect 30941 11101 30975 11135
rect 30975 11101 30984 11135
rect 30932 11092 30984 11101
rect 37832 11092 37884 11144
rect 39488 11092 39540 11144
rect 39948 11092 40000 11144
rect 43904 11135 43956 11144
rect 43904 11101 43913 11135
rect 43913 11101 43947 11135
rect 43947 11101 43956 11135
rect 43904 11092 43956 11101
rect 44548 11135 44600 11144
rect 44548 11101 44557 11135
rect 44557 11101 44591 11135
rect 44591 11101 44600 11135
rect 44548 11092 44600 11101
rect 39304 11024 39356 11076
rect 19524 10956 19576 11008
rect 23848 10999 23900 11008
rect 23848 10965 23857 10999
rect 23857 10965 23891 10999
rect 23891 10965 23900 10999
rect 23848 10956 23900 10965
rect 25504 10999 25556 11008
rect 25504 10965 25513 10999
rect 25513 10965 25547 10999
rect 25547 10965 25556 10999
rect 25504 10956 25556 10965
rect 26792 10999 26844 11008
rect 26792 10965 26801 10999
rect 26801 10965 26835 10999
rect 26835 10965 26844 10999
rect 26792 10956 26844 10965
rect 27528 10956 27580 11008
rect 37740 10956 37792 11008
rect 40500 10999 40552 11008
rect 40500 10965 40509 10999
rect 40509 10965 40543 10999
rect 40543 10965 40552 10999
rect 40500 10956 40552 10965
rect 41604 10999 41656 11008
rect 41604 10965 41613 10999
rect 41613 10965 41647 10999
rect 41647 10965 41656 10999
rect 41604 10956 41656 10965
rect 46020 10956 46072 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 16120 10752 16172 10804
rect 18972 10752 19024 10804
rect 19156 10795 19208 10804
rect 19156 10761 19165 10795
rect 19165 10761 19199 10795
rect 19199 10761 19208 10795
rect 19156 10752 19208 10761
rect 17776 10684 17828 10736
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 23388 10795 23440 10804
rect 20076 10727 20128 10736
rect 20076 10693 20085 10727
rect 20085 10693 20119 10727
rect 20119 10693 20128 10727
rect 20076 10684 20128 10693
rect 16304 10480 16356 10532
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 19984 10616 20036 10668
rect 23388 10761 23397 10795
rect 23397 10761 23431 10795
rect 23431 10761 23440 10795
rect 23388 10752 23440 10761
rect 25320 10752 25372 10804
rect 26700 10752 26752 10804
rect 29000 10752 29052 10804
rect 29276 10752 29328 10804
rect 31300 10795 31352 10804
rect 31300 10761 31309 10795
rect 31309 10761 31343 10795
rect 31343 10761 31352 10795
rect 31300 10752 31352 10761
rect 33600 10752 33652 10804
rect 33876 10752 33928 10804
rect 37280 10795 37332 10804
rect 37280 10761 37289 10795
rect 37289 10761 37323 10795
rect 37323 10761 37332 10795
rect 37280 10752 37332 10761
rect 39856 10752 39908 10804
rect 40868 10752 40920 10804
rect 41604 10752 41656 10804
rect 30472 10684 30524 10736
rect 21732 10659 21784 10668
rect 21732 10625 21741 10659
rect 21741 10625 21775 10659
rect 21775 10625 21784 10659
rect 21732 10616 21784 10625
rect 24768 10616 24820 10668
rect 30932 10616 30984 10668
rect 32312 10616 32364 10668
rect 34612 10659 34664 10668
rect 34612 10625 34621 10659
rect 34621 10625 34655 10659
rect 34655 10625 34664 10659
rect 42064 10684 42116 10736
rect 34612 10616 34664 10625
rect 35716 10616 35768 10668
rect 36084 10659 36136 10668
rect 36084 10625 36093 10659
rect 36093 10625 36127 10659
rect 36127 10625 36136 10659
rect 36084 10616 36136 10625
rect 37832 10659 37884 10668
rect 37832 10625 37841 10659
rect 37841 10625 37875 10659
rect 37875 10625 37884 10659
rect 37832 10616 37884 10625
rect 39580 10616 39632 10668
rect 41144 10616 41196 10668
rect 21640 10548 21692 10600
rect 27528 10548 27580 10600
rect 30380 10591 30432 10600
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 17868 10412 17920 10464
rect 18788 10412 18840 10464
rect 19432 10412 19484 10464
rect 23572 10480 23624 10532
rect 24952 10480 25004 10532
rect 27068 10480 27120 10532
rect 28540 10480 28592 10532
rect 22652 10455 22704 10464
rect 22652 10421 22661 10455
rect 22661 10421 22695 10455
rect 22695 10421 22704 10455
rect 22652 10412 22704 10421
rect 24584 10412 24636 10464
rect 28356 10455 28408 10464
rect 28356 10421 28365 10455
rect 28365 10421 28399 10455
rect 28399 10421 28408 10455
rect 28356 10412 28408 10421
rect 28632 10455 28684 10464
rect 28632 10421 28641 10455
rect 28641 10421 28675 10455
rect 28675 10421 28684 10455
rect 28632 10412 28684 10421
rect 30380 10557 30389 10591
rect 30389 10557 30423 10591
rect 30423 10557 30432 10591
rect 30380 10548 30432 10557
rect 30472 10548 30524 10600
rect 33416 10548 33468 10600
rect 33508 10548 33560 10600
rect 38752 10548 38804 10600
rect 42248 10548 42300 10600
rect 43720 10752 43772 10804
rect 43904 10752 43956 10804
rect 45192 10752 45244 10804
rect 47492 10752 47544 10804
rect 43996 10684 44048 10736
rect 44548 10727 44600 10736
rect 44548 10693 44557 10727
rect 44557 10693 44591 10727
rect 44591 10693 44600 10727
rect 44548 10684 44600 10693
rect 44088 10616 44140 10668
rect 46756 10591 46808 10600
rect 46756 10557 46765 10591
rect 46765 10557 46799 10591
rect 46799 10557 46808 10591
rect 46756 10548 46808 10557
rect 35716 10480 35768 10532
rect 38016 10480 38068 10532
rect 40868 10480 40920 10532
rect 43812 10480 43864 10532
rect 44088 10523 44140 10532
rect 44088 10489 44097 10523
rect 44097 10489 44131 10523
rect 44131 10489 44140 10523
rect 46112 10523 46164 10532
rect 44088 10480 44140 10489
rect 46112 10489 46121 10523
rect 46121 10489 46155 10523
rect 46155 10489 46164 10523
rect 46112 10480 46164 10489
rect 30104 10412 30156 10464
rect 32128 10412 32180 10464
rect 35532 10412 35584 10464
rect 37004 10455 37056 10464
rect 37004 10421 37013 10455
rect 37013 10421 37047 10455
rect 37047 10421 37056 10455
rect 37004 10412 37056 10421
rect 38752 10455 38804 10464
rect 38752 10421 38761 10455
rect 38761 10421 38795 10455
rect 38795 10421 38804 10455
rect 38752 10412 38804 10421
rect 39488 10455 39540 10464
rect 39488 10421 39497 10455
rect 39497 10421 39531 10455
rect 39531 10421 39540 10455
rect 39488 10412 39540 10421
rect 39948 10455 40000 10464
rect 39948 10421 39957 10455
rect 39957 10421 39991 10455
rect 39991 10421 40000 10455
rect 39948 10412 40000 10421
rect 42524 10412 42576 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 17500 10208 17552 10260
rect 19984 10208 20036 10260
rect 21640 10251 21692 10260
rect 21640 10217 21649 10251
rect 21649 10217 21683 10251
rect 21683 10217 21692 10251
rect 21640 10208 21692 10217
rect 21732 10208 21784 10260
rect 23848 10208 23900 10260
rect 24584 10208 24636 10260
rect 24768 10208 24820 10260
rect 26792 10208 26844 10260
rect 28448 10251 28500 10260
rect 28448 10217 28457 10251
rect 28457 10217 28491 10251
rect 28491 10217 28500 10251
rect 28448 10208 28500 10217
rect 30012 10251 30064 10260
rect 30012 10217 30021 10251
rect 30021 10217 30055 10251
rect 30055 10217 30064 10251
rect 30012 10208 30064 10217
rect 30380 10208 30432 10260
rect 32312 10251 32364 10260
rect 32312 10217 32321 10251
rect 32321 10217 32355 10251
rect 32355 10217 32364 10251
rect 32312 10208 32364 10217
rect 36084 10251 36136 10260
rect 36084 10217 36093 10251
rect 36093 10217 36127 10251
rect 36127 10217 36136 10251
rect 36084 10208 36136 10217
rect 37832 10208 37884 10260
rect 39948 10208 40000 10260
rect 41144 10251 41196 10260
rect 41144 10217 41153 10251
rect 41153 10217 41187 10251
rect 41187 10217 41196 10251
rect 41144 10208 41196 10217
rect 43812 10208 43864 10260
rect 46756 10208 46808 10260
rect 18236 10140 18288 10192
rect 16120 10072 16172 10124
rect 19156 10072 19208 10124
rect 21456 10072 21508 10124
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 22008 10004 22060 10056
rect 22652 10072 22704 10124
rect 24860 10140 24912 10192
rect 27068 10140 27120 10192
rect 33692 10140 33744 10192
rect 39028 10140 39080 10192
rect 41788 10183 41840 10192
rect 41788 10149 41797 10183
rect 41797 10149 41831 10183
rect 41831 10149 41840 10183
rect 41788 10140 41840 10149
rect 42248 10140 42300 10192
rect 43076 10140 43128 10192
rect 43904 10140 43956 10192
rect 44088 10140 44140 10192
rect 24216 10072 24268 10124
rect 25504 10072 25556 10124
rect 26240 10072 26292 10124
rect 28172 10072 28224 10124
rect 28724 10072 28776 10124
rect 30380 10115 30432 10124
rect 30380 10081 30389 10115
rect 30389 10081 30423 10115
rect 30423 10081 30432 10115
rect 30380 10072 30432 10081
rect 33048 10115 33100 10124
rect 30012 10004 30064 10056
rect 30656 10004 30708 10056
rect 33048 10081 33057 10115
rect 33057 10081 33091 10115
rect 33091 10081 33100 10115
rect 33048 10072 33100 10081
rect 35532 10072 35584 10124
rect 36452 10115 36504 10124
rect 36452 10081 36461 10115
rect 36461 10081 36495 10115
rect 36495 10081 36504 10115
rect 36452 10072 36504 10081
rect 39672 10072 39724 10124
rect 40132 10115 40184 10124
rect 40132 10081 40141 10115
rect 40141 10081 40175 10115
rect 40175 10081 40184 10115
rect 40132 10072 40184 10081
rect 40960 10072 41012 10124
rect 46020 10115 46072 10124
rect 46020 10081 46029 10115
rect 46029 10081 46063 10115
rect 46063 10081 46072 10115
rect 46020 10072 46072 10081
rect 47492 10115 47544 10124
rect 47492 10081 47501 10115
rect 47501 10081 47535 10115
rect 47535 10081 47544 10115
rect 47492 10072 47544 10081
rect 35624 10047 35676 10056
rect 35624 10013 35633 10047
rect 35633 10013 35667 10047
rect 35667 10013 35676 10047
rect 35624 10004 35676 10013
rect 38660 10047 38712 10056
rect 38660 10013 38669 10047
rect 38669 10013 38703 10047
rect 38703 10013 38712 10047
rect 38660 10004 38712 10013
rect 43904 10047 43956 10056
rect 43904 10013 43913 10047
rect 43913 10013 43947 10047
rect 43947 10013 43956 10047
rect 43904 10004 43956 10013
rect 45928 10047 45980 10056
rect 45928 10013 45937 10047
rect 45937 10013 45971 10047
rect 45971 10013 45980 10047
rect 45928 10004 45980 10013
rect 35256 9936 35308 9988
rect 35808 9936 35860 9988
rect 44456 9979 44508 9988
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 27436 9868 27488 9920
rect 29276 9911 29328 9920
rect 29276 9877 29285 9911
rect 29285 9877 29319 9911
rect 29319 9877 29328 9911
rect 29276 9868 29328 9877
rect 30104 9868 30156 9920
rect 35900 9868 35952 9920
rect 44456 9945 44465 9979
rect 44465 9945 44499 9979
rect 44499 9945 44508 9979
rect 44456 9936 44508 9945
rect 39304 9868 39356 9920
rect 43812 9868 43864 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 16120 9664 16172 9716
rect 17868 9664 17920 9716
rect 22008 9707 22060 9716
rect 22008 9673 22017 9707
rect 22017 9673 22051 9707
rect 22051 9673 22060 9707
rect 22008 9664 22060 9673
rect 22652 9664 22704 9716
rect 25688 9707 25740 9716
rect 25688 9673 25697 9707
rect 25697 9673 25731 9707
rect 25731 9673 25740 9707
rect 25688 9664 25740 9673
rect 29184 9664 29236 9716
rect 30380 9707 30432 9716
rect 30380 9673 30389 9707
rect 30389 9673 30423 9707
rect 30423 9673 30432 9707
rect 30380 9664 30432 9673
rect 30656 9707 30708 9716
rect 30656 9673 30665 9707
rect 30665 9673 30699 9707
rect 30699 9673 30708 9707
rect 30656 9664 30708 9673
rect 32404 9707 32456 9716
rect 32404 9673 32413 9707
rect 32413 9673 32447 9707
rect 32447 9673 32456 9707
rect 32404 9664 32456 9673
rect 32680 9707 32732 9716
rect 32680 9673 32689 9707
rect 32689 9673 32723 9707
rect 32723 9673 32732 9707
rect 32680 9664 32732 9673
rect 33048 9664 33100 9716
rect 33692 9707 33744 9716
rect 33692 9673 33701 9707
rect 33701 9673 33735 9707
rect 33735 9673 33744 9707
rect 33692 9664 33744 9673
rect 35532 9664 35584 9716
rect 36452 9664 36504 9716
rect 38660 9664 38712 9716
rect 39028 9707 39080 9716
rect 39028 9673 39037 9707
rect 39037 9673 39071 9707
rect 39071 9673 39080 9707
rect 39028 9664 39080 9673
rect 39488 9664 39540 9716
rect 40960 9707 41012 9716
rect 40960 9673 40969 9707
rect 40969 9673 41003 9707
rect 41003 9673 41012 9707
rect 40960 9664 41012 9673
rect 41880 9664 41932 9716
rect 42248 9664 42300 9716
rect 44088 9664 44140 9716
rect 45928 9707 45980 9716
rect 45928 9673 45937 9707
rect 45937 9673 45971 9707
rect 45971 9673 45980 9707
rect 45928 9664 45980 9673
rect 47492 9707 47544 9716
rect 47492 9673 47501 9707
rect 47501 9673 47535 9707
rect 47535 9673 47544 9707
rect 47492 9664 47544 9673
rect 10968 9392 11020 9444
rect 16212 9460 16264 9512
rect 19156 9528 19208 9580
rect 19432 9528 19484 9580
rect 18144 9392 18196 9444
rect 20168 9503 20220 9512
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 18604 9324 18656 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 23756 9503 23808 9512
rect 23480 9460 23532 9469
rect 23756 9469 23765 9503
rect 23765 9469 23799 9503
rect 23799 9469 23808 9503
rect 23756 9460 23808 9469
rect 23848 9460 23900 9512
rect 24124 9460 24176 9512
rect 25688 9460 25740 9512
rect 26516 9435 26568 9444
rect 26516 9401 26525 9435
rect 26525 9401 26559 9435
rect 26559 9401 26568 9435
rect 26516 9392 26568 9401
rect 27988 9460 28040 9512
rect 29000 9460 29052 9512
rect 29184 9460 29236 9512
rect 29368 9460 29420 9512
rect 35256 9596 35308 9648
rect 35716 9639 35768 9648
rect 35716 9605 35725 9639
rect 35725 9605 35759 9639
rect 35759 9605 35768 9639
rect 35716 9596 35768 9605
rect 40132 9639 40184 9648
rect 40132 9605 40141 9639
rect 40141 9605 40175 9639
rect 40175 9605 40184 9639
rect 40132 9596 40184 9605
rect 43076 9639 43128 9648
rect 43076 9605 43085 9639
rect 43085 9605 43119 9639
rect 43119 9605 43128 9639
rect 43076 9596 43128 9605
rect 46020 9596 46072 9648
rect 35624 9528 35676 9580
rect 37004 9528 37056 9580
rect 30196 9460 30248 9512
rect 32404 9460 32456 9512
rect 32680 9460 32732 9512
rect 34428 9460 34480 9512
rect 42524 9571 42576 9580
rect 42524 9537 42533 9571
rect 42533 9537 42567 9571
rect 42567 9537 42576 9571
rect 42524 9528 42576 9537
rect 43260 9528 43312 9580
rect 43904 9528 43956 9580
rect 46388 9528 46440 9580
rect 38752 9460 38804 9512
rect 30012 9392 30064 9444
rect 30380 9392 30432 9444
rect 35716 9392 35768 9444
rect 19984 9324 20036 9376
rect 21456 9324 21508 9376
rect 22928 9324 22980 9376
rect 23112 9367 23164 9376
rect 23112 9333 23121 9367
rect 23121 9333 23155 9367
rect 23155 9333 23164 9367
rect 23112 9324 23164 9333
rect 23848 9367 23900 9376
rect 23848 9333 23857 9367
rect 23857 9333 23891 9367
rect 23891 9333 23900 9367
rect 23848 9324 23900 9333
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 27068 9324 27120 9376
rect 27528 9324 27580 9376
rect 29644 9324 29696 9376
rect 32588 9324 32640 9376
rect 33048 9367 33100 9376
rect 33048 9333 33057 9367
rect 33057 9333 33091 9367
rect 33091 9333 33100 9367
rect 33048 9324 33100 9333
rect 36912 9324 36964 9376
rect 37740 9367 37792 9376
rect 37740 9333 37749 9367
rect 37749 9333 37783 9367
rect 37783 9333 37792 9367
rect 37740 9324 37792 9333
rect 42156 9324 42208 9376
rect 44088 9435 44140 9444
rect 44088 9401 44097 9435
rect 44097 9401 44131 9435
rect 44131 9401 44140 9435
rect 44088 9392 44140 9401
rect 46848 9435 46900 9444
rect 45928 9324 45980 9376
rect 46848 9401 46857 9435
rect 46857 9401 46891 9435
rect 46891 9401 46900 9435
rect 46848 9392 46900 9401
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 17868 9120 17920 9172
rect 17960 9120 18012 9172
rect 20168 9120 20220 9172
rect 24216 9163 24268 9172
rect 24216 9129 24225 9163
rect 24225 9129 24259 9163
rect 24259 9129 24268 9163
rect 24216 9120 24268 9129
rect 25688 9120 25740 9172
rect 26240 9163 26292 9172
rect 26240 9129 26249 9163
rect 26249 9129 26283 9163
rect 26283 9129 26292 9163
rect 26240 9120 26292 9129
rect 27988 9120 28040 9172
rect 28172 9163 28224 9172
rect 28172 9129 28181 9163
rect 28181 9129 28215 9163
rect 28215 9129 28224 9163
rect 28172 9120 28224 9129
rect 30840 9120 30892 9172
rect 35532 9163 35584 9172
rect 35532 9129 35541 9163
rect 35541 9129 35575 9163
rect 35575 9129 35584 9163
rect 35532 9120 35584 9129
rect 35624 9120 35676 9172
rect 38016 9120 38068 9172
rect 39856 9163 39908 9172
rect 39856 9129 39865 9163
rect 39865 9129 39899 9163
rect 39899 9129 39908 9163
rect 39856 9120 39908 9129
rect 41788 9120 41840 9172
rect 42524 9120 42576 9172
rect 44088 9120 44140 9172
rect 18604 9052 18656 9104
rect 18696 9027 18748 9036
rect 18696 8993 18705 9027
rect 18705 8993 18739 9027
rect 18739 8993 18748 9027
rect 18696 8984 18748 8993
rect 18788 8984 18840 9036
rect 20076 8984 20128 9036
rect 27068 9052 27120 9104
rect 21640 8984 21692 9036
rect 22744 8984 22796 9036
rect 24032 8984 24084 9036
rect 24952 8984 25004 9036
rect 28816 8984 28868 9036
rect 29276 8984 29328 9036
rect 30840 8984 30892 9036
rect 32128 8984 32180 9036
rect 32588 9027 32640 9036
rect 32588 8993 32597 9027
rect 32597 8993 32631 9027
rect 32631 8993 32640 9027
rect 32588 8984 32640 8993
rect 32956 8984 33008 9036
rect 33416 8984 33468 9036
rect 34428 9027 34480 9036
rect 34428 8993 34437 9027
rect 34437 8993 34471 9027
rect 34471 8993 34480 9027
rect 34428 8984 34480 8993
rect 41880 9095 41932 9104
rect 41880 9061 41889 9095
rect 41889 9061 41923 9095
rect 41923 9061 41932 9095
rect 41880 9052 41932 9061
rect 43260 9052 43312 9104
rect 43536 9095 43588 9104
rect 43536 9061 43545 9095
rect 43545 9061 43579 9095
rect 43579 9061 43588 9095
rect 43536 9052 43588 9061
rect 46112 9052 46164 9104
rect 36084 9027 36136 9036
rect 36084 8993 36093 9027
rect 36093 8993 36127 9027
rect 36127 8993 36136 9027
rect 36084 8984 36136 8993
rect 36360 8984 36412 9036
rect 47216 9027 47268 9036
rect 47216 8993 47225 9027
rect 47225 8993 47259 9027
rect 47259 8993 47268 9027
rect 47216 8984 47268 8993
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 25044 8916 25096 8968
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 29552 8916 29604 8968
rect 34796 8916 34848 8968
rect 36728 8916 36780 8968
rect 38108 8916 38160 8968
rect 39488 8959 39540 8968
rect 39488 8925 39497 8959
rect 39497 8925 39531 8959
rect 39531 8925 39540 8959
rect 39488 8916 39540 8925
rect 41788 8959 41840 8968
rect 41788 8925 41797 8959
rect 41797 8925 41831 8959
rect 41831 8925 41840 8959
rect 43444 8959 43496 8968
rect 41788 8916 41840 8925
rect 43444 8925 43453 8959
rect 43453 8925 43487 8959
rect 43487 8925 43496 8959
rect 43444 8916 43496 8925
rect 43720 8959 43772 8968
rect 43720 8925 43729 8959
rect 43729 8925 43763 8959
rect 43763 8925 43772 8959
rect 43720 8916 43772 8925
rect 45744 8959 45796 8968
rect 45744 8925 45753 8959
rect 45753 8925 45787 8959
rect 45787 8925 45796 8959
rect 45744 8916 45796 8925
rect 46020 8959 46072 8968
rect 46020 8925 46029 8959
rect 46029 8925 46063 8959
rect 46063 8925 46072 8959
rect 46020 8916 46072 8925
rect 46848 8916 46900 8968
rect 23940 8780 23992 8832
rect 27620 8780 27672 8832
rect 33692 8823 33744 8832
rect 33692 8789 33701 8823
rect 33701 8789 33735 8823
rect 33735 8789 33744 8823
rect 33692 8780 33744 8789
rect 38660 8823 38712 8832
rect 38660 8789 38669 8823
rect 38669 8789 38703 8823
rect 38703 8789 38712 8823
rect 38660 8780 38712 8789
rect 47492 8848 47544 8900
rect 45928 8780 45980 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 21640 8619 21692 8628
rect 21640 8585 21649 8619
rect 21649 8585 21683 8619
rect 21683 8585 21692 8619
rect 21640 8576 21692 8585
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 23112 8576 23164 8628
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 26516 8576 26568 8628
rect 27436 8576 27488 8628
rect 28816 8576 28868 8628
rect 30840 8619 30892 8628
rect 30840 8585 30849 8619
rect 30849 8585 30883 8619
rect 30883 8585 30892 8619
rect 30840 8576 30892 8585
rect 32588 8619 32640 8628
rect 32588 8585 32597 8619
rect 32597 8585 32631 8619
rect 32631 8585 32640 8619
rect 32588 8576 32640 8585
rect 33048 8619 33100 8628
rect 33048 8585 33057 8619
rect 33057 8585 33091 8619
rect 33091 8585 33100 8619
rect 33048 8576 33100 8585
rect 34428 8619 34480 8628
rect 34428 8585 34437 8619
rect 34437 8585 34471 8619
rect 34471 8585 34480 8619
rect 34428 8576 34480 8585
rect 38108 8619 38160 8628
rect 38108 8585 38117 8619
rect 38117 8585 38151 8619
rect 38151 8585 38160 8619
rect 38108 8576 38160 8585
rect 41788 8576 41840 8628
rect 41880 8576 41932 8628
rect 43536 8576 43588 8628
rect 45744 8576 45796 8628
rect 18696 8440 18748 8492
rect 24032 8508 24084 8560
rect 25688 8508 25740 8560
rect 28448 8508 28500 8560
rect 29276 8508 29328 8560
rect 23848 8440 23900 8492
rect 29552 8483 29604 8492
rect 29552 8449 29561 8483
rect 29561 8449 29595 8483
rect 29595 8449 29604 8483
rect 29552 8440 29604 8449
rect 28356 8372 28408 8424
rect 29000 8372 29052 8424
rect 31576 8508 31628 8560
rect 39764 8508 39816 8560
rect 43444 8508 43496 8560
rect 46296 8508 46348 8560
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 31484 8440 31536 8492
rect 33692 8440 33744 8492
rect 33048 8372 33100 8424
rect 34336 8372 34388 8424
rect 34888 8415 34940 8424
rect 34888 8381 34897 8415
rect 34897 8381 34931 8415
rect 34931 8381 34940 8415
rect 34888 8372 34940 8381
rect 39488 8440 39540 8492
rect 43720 8440 43772 8492
rect 46112 8440 46164 8492
rect 35532 8372 35584 8424
rect 36636 8372 36688 8424
rect 36820 8372 36872 8424
rect 19156 8347 19208 8356
rect 19156 8313 19165 8347
rect 19165 8313 19199 8347
rect 19199 8313 19208 8347
rect 19156 8304 19208 8313
rect 19432 8304 19484 8356
rect 20720 8347 20772 8356
rect 20720 8313 20729 8347
rect 20729 8313 20763 8347
rect 20763 8313 20772 8347
rect 20720 8304 20772 8313
rect 20904 8304 20956 8356
rect 23572 8304 23624 8356
rect 26056 8347 26108 8356
rect 26056 8313 26065 8347
rect 26065 8313 26099 8347
rect 26099 8313 26108 8347
rect 26056 8304 26108 8313
rect 26700 8347 26752 8356
rect 23664 8236 23716 8288
rect 26700 8313 26709 8347
rect 26709 8313 26743 8347
rect 26743 8313 26752 8347
rect 26700 8304 26752 8313
rect 27068 8279 27120 8288
rect 27068 8245 27077 8279
rect 27077 8245 27111 8279
rect 27111 8245 27120 8279
rect 30288 8304 30340 8356
rect 31576 8304 31628 8356
rect 39120 8372 39172 8424
rect 44272 8415 44324 8424
rect 38752 8304 38804 8356
rect 30472 8279 30524 8288
rect 27068 8236 27120 8245
rect 30472 8245 30481 8279
rect 30481 8245 30515 8279
rect 30515 8245 30524 8279
rect 30472 8236 30524 8245
rect 36084 8279 36136 8288
rect 36084 8245 36093 8279
rect 36093 8245 36127 8279
rect 36127 8245 36136 8279
rect 36084 8236 36136 8245
rect 36636 8236 36688 8288
rect 37004 8279 37056 8288
rect 37004 8245 37013 8279
rect 37013 8245 37047 8279
rect 37047 8245 37056 8279
rect 37004 8236 37056 8245
rect 38016 8236 38068 8288
rect 39580 8279 39632 8288
rect 39580 8245 39589 8279
rect 39589 8245 39623 8279
rect 39623 8245 39632 8279
rect 39580 8236 39632 8245
rect 39856 8279 39908 8288
rect 39856 8245 39865 8279
rect 39865 8245 39899 8279
rect 39899 8245 39908 8279
rect 39856 8236 39908 8245
rect 41512 8347 41564 8356
rect 41512 8313 41521 8347
rect 41521 8313 41555 8347
rect 41555 8313 41564 8347
rect 41512 8304 41564 8313
rect 42156 8304 42208 8356
rect 44272 8381 44281 8415
rect 44281 8381 44315 8415
rect 44315 8381 44324 8415
rect 44272 8372 44324 8381
rect 46204 8415 46256 8424
rect 46204 8381 46213 8415
rect 46213 8381 46247 8415
rect 46247 8381 46256 8415
rect 46204 8372 46256 8381
rect 43812 8304 43864 8356
rect 46112 8347 46164 8356
rect 46112 8313 46121 8347
rect 46121 8313 46155 8347
rect 46155 8313 46164 8347
rect 46112 8304 46164 8313
rect 44364 8236 44416 8288
rect 47216 8279 47268 8288
rect 47216 8245 47225 8279
rect 47225 8245 47259 8279
rect 47259 8245 47268 8279
rect 47216 8236 47268 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 23664 8075 23716 8084
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 23848 8032 23900 8084
rect 28356 8032 28408 8084
rect 32956 8032 33008 8084
rect 34888 8075 34940 8084
rect 34888 8041 34897 8075
rect 34897 8041 34931 8075
rect 34931 8041 34940 8075
rect 34888 8032 34940 8041
rect 36360 8075 36412 8084
rect 36360 8041 36369 8075
rect 36369 8041 36403 8075
rect 36403 8041 36412 8075
rect 36360 8032 36412 8041
rect 36820 8075 36872 8084
rect 36820 8041 36829 8075
rect 36829 8041 36863 8075
rect 36863 8041 36872 8075
rect 36820 8032 36872 8041
rect 38752 8075 38804 8084
rect 38752 8041 38761 8075
rect 38761 8041 38795 8075
rect 38795 8041 38804 8075
rect 38752 8032 38804 8041
rect 44272 8075 44324 8084
rect 44272 8041 44281 8075
rect 44281 8041 44315 8075
rect 44315 8041 44324 8075
rect 44272 8032 44324 8041
rect 46296 8032 46348 8084
rect 21088 8007 21140 8016
rect 21088 7973 21097 8007
rect 21097 7973 21131 8007
rect 21131 7973 21140 8007
rect 21088 7964 21140 7973
rect 22928 7964 22980 8016
rect 24952 8007 25004 8016
rect 24952 7973 24961 8007
rect 24961 7973 24995 8007
rect 24995 7973 25004 8007
rect 24952 7964 25004 7973
rect 25044 8007 25096 8016
rect 25044 7973 25053 8007
rect 25053 7973 25087 8007
rect 25087 7973 25096 8007
rect 25044 7964 25096 7973
rect 26608 7964 26660 8016
rect 26792 7964 26844 8016
rect 28172 7964 28224 8016
rect 30288 7964 30340 8016
rect 33784 7964 33836 8016
rect 35716 7964 35768 8016
rect 39856 7964 39908 8016
rect 45008 8007 45060 8016
rect 45008 7973 45017 8007
rect 45017 7973 45051 8007
rect 45051 7973 45060 8007
rect 45008 7964 45060 7973
rect 45744 7964 45796 8016
rect 46204 8007 46256 8016
rect 46204 7973 46213 8007
rect 46213 7973 46247 8007
rect 46247 7973 46256 8007
rect 46204 7964 46256 7973
rect 18880 7896 18932 7948
rect 19432 7939 19484 7948
rect 19432 7905 19476 7939
rect 19476 7905 19484 7939
rect 19432 7896 19484 7905
rect 23940 7896 23992 7948
rect 29644 7939 29696 7948
rect 29644 7905 29653 7939
rect 29653 7905 29687 7939
rect 29687 7905 29696 7939
rect 29644 7896 29696 7905
rect 32220 7896 32272 7948
rect 34796 7896 34848 7948
rect 38476 7896 38528 7948
rect 41696 7939 41748 7948
rect 41696 7905 41705 7939
rect 41705 7905 41739 7939
rect 41739 7905 41748 7939
rect 41696 7896 41748 7905
rect 42340 7939 42392 7948
rect 42340 7905 42349 7939
rect 42349 7905 42383 7939
rect 42383 7905 42392 7939
rect 42340 7896 42392 7905
rect 43812 7939 43864 7948
rect 43812 7905 43821 7939
rect 43821 7905 43855 7939
rect 43855 7905 43864 7939
rect 43812 7896 43864 7905
rect 45928 7896 45980 7948
rect 47124 7896 47176 7948
rect 47400 7939 47452 7948
rect 47400 7905 47409 7939
rect 47409 7905 47443 7939
rect 47443 7905 47452 7939
rect 47400 7896 47452 7905
rect 22652 7828 22704 7880
rect 19156 7803 19208 7812
rect 19156 7769 19165 7803
rect 19165 7769 19199 7803
rect 19199 7769 19208 7803
rect 20720 7803 20772 7812
rect 19156 7760 19208 7769
rect 19800 7692 19852 7744
rect 20720 7769 20729 7803
rect 20729 7769 20763 7803
rect 20763 7769 20772 7803
rect 20720 7760 20772 7769
rect 21640 7760 21692 7812
rect 26700 7828 26752 7880
rect 28264 7828 28316 7880
rect 33324 7871 33376 7880
rect 33324 7837 33333 7871
rect 33333 7837 33367 7871
rect 33367 7837 33376 7871
rect 33324 7828 33376 7837
rect 35532 7828 35584 7880
rect 36728 7828 36780 7880
rect 39120 7828 39172 7880
rect 41512 7871 41564 7880
rect 41512 7837 41521 7871
rect 41521 7837 41555 7871
rect 41555 7837 41564 7871
rect 41512 7828 41564 7837
rect 42616 7828 42668 7880
rect 44456 7828 44508 7880
rect 47492 7828 47544 7880
rect 35440 7760 35492 7812
rect 40224 7760 40276 7812
rect 43904 7760 43956 7812
rect 46204 7760 46256 7812
rect 21732 7692 21784 7744
rect 26056 7735 26108 7744
rect 26056 7701 26065 7735
rect 26065 7701 26099 7735
rect 26099 7701 26108 7735
rect 26056 7692 26108 7701
rect 30656 7692 30708 7744
rect 30840 7735 30892 7744
rect 30840 7701 30849 7735
rect 30849 7701 30883 7735
rect 30883 7701 30892 7735
rect 30840 7692 30892 7701
rect 31300 7735 31352 7744
rect 31300 7701 31309 7735
rect 31309 7701 31343 7735
rect 31343 7701 31352 7735
rect 31300 7692 31352 7701
rect 35992 7735 36044 7744
rect 35992 7701 36001 7735
rect 36001 7701 36035 7735
rect 36035 7701 36044 7735
rect 35992 7692 36044 7701
rect 44456 7692 44508 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 22652 7531 22704 7540
rect 22652 7497 22661 7531
rect 22661 7497 22695 7531
rect 22695 7497 22704 7531
rect 22652 7488 22704 7497
rect 23940 7488 23992 7540
rect 24124 7531 24176 7540
rect 24124 7497 24133 7531
rect 24133 7497 24167 7531
rect 24167 7497 24176 7531
rect 24124 7488 24176 7497
rect 24952 7488 25004 7540
rect 26056 7488 26108 7540
rect 28172 7531 28224 7540
rect 28172 7497 28181 7531
rect 28181 7497 28215 7531
rect 28215 7497 28224 7531
rect 28172 7488 28224 7497
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 19800 7327 19852 7336
rect 19800 7293 19809 7327
rect 19809 7293 19843 7327
rect 19843 7293 19852 7327
rect 19800 7284 19852 7293
rect 21732 7216 21784 7268
rect 24400 7352 24452 7404
rect 25044 7352 25096 7404
rect 24124 7284 24176 7336
rect 27620 7284 27672 7336
rect 30472 7488 30524 7540
rect 32220 7531 32272 7540
rect 32220 7497 32229 7531
rect 32229 7497 32263 7531
rect 32263 7497 32272 7531
rect 32220 7488 32272 7497
rect 32588 7531 32640 7540
rect 32588 7497 32597 7531
rect 32597 7497 32631 7531
rect 32631 7497 32640 7531
rect 32588 7488 32640 7497
rect 33784 7531 33836 7540
rect 33784 7497 33793 7531
rect 33793 7497 33827 7531
rect 33827 7497 33836 7531
rect 33784 7488 33836 7497
rect 35716 7488 35768 7540
rect 37004 7531 37056 7540
rect 37004 7497 37013 7531
rect 37013 7497 37047 7531
rect 37047 7497 37056 7531
rect 37004 7488 37056 7497
rect 38476 7531 38528 7540
rect 38476 7497 38485 7531
rect 38485 7497 38519 7531
rect 38519 7497 38528 7531
rect 38476 7488 38528 7497
rect 39120 7531 39172 7540
rect 39120 7497 39129 7531
rect 39129 7497 39163 7531
rect 39163 7497 39172 7531
rect 39120 7488 39172 7497
rect 42340 7488 42392 7540
rect 42616 7488 42668 7540
rect 43812 7531 43864 7540
rect 43812 7497 43821 7531
rect 43821 7497 43855 7531
rect 43855 7497 43864 7531
rect 43812 7488 43864 7497
rect 44364 7531 44416 7540
rect 44364 7497 44373 7531
rect 44373 7497 44407 7531
rect 44407 7497 44416 7531
rect 44364 7488 44416 7497
rect 45008 7488 45060 7540
rect 46112 7488 46164 7540
rect 47124 7531 47176 7540
rect 47124 7497 47133 7531
rect 47133 7497 47167 7531
rect 47167 7497 47176 7531
rect 47124 7488 47176 7497
rect 30288 7463 30340 7472
rect 30288 7429 30297 7463
rect 30297 7429 30331 7463
rect 30331 7429 30340 7463
rect 30288 7420 30340 7429
rect 30840 7395 30892 7404
rect 30840 7361 30849 7395
rect 30849 7361 30883 7395
rect 30883 7361 30892 7395
rect 30840 7352 30892 7361
rect 31484 7395 31536 7404
rect 31484 7361 31493 7395
rect 31493 7361 31527 7395
rect 31527 7361 31536 7395
rect 31484 7352 31536 7361
rect 33324 7352 33376 7404
rect 35624 7395 35676 7404
rect 35624 7361 35633 7395
rect 35633 7361 35667 7395
rect 35667 7361 35676 7395
rect 35624 7352 35676 7361
rect 39580 7420 39632 7472
rect 40684 7352 40736 7404
rect 32588 7284 32640 7336
rect 32772 7284 32824 7336
rect 38660 7284 38712 7336
rect 28264 7216 28316 7268
rect 30932 7259 30984 7268
rect 22468 7148 22520 7200
rect 24584 7148 24636 7200
rect 25964 7191 26016 7200
rect 25964 7157 25973 7191
rect 25973 7157 26007 7191
rect 26007 7157 26016 7191
rect 25964 7148 26016 7157
rect 26424 7191 26476 7200
rect 26424 7157 26433 7191
rect 26433 7157 26467 7191
rect 26467 7157 26476 7191
rect 26424 7148 26476 7157
rect 26792 7148 26844 7200
rect 30564 7191 30616 7200
rect 30564 7157 30573 7191
rect 30573 7157 30607 7191
rect 30607 7157 30616 7191
rect 30564 7148 30616 7157
rect 30932 7225 30941 7259
rect 30941 7225 30975 7259
rect 30975 7225 30984 7259
rect 30932 7216 30984 7225
rect 35716 7259 35768 7268
rect 35716 7225 35725 7259
rect 35725 7225 35759 7259
rect 35759 7225 35768 7259
rect 35716 7216 35768 7225
rect 36268 7259 36320 7268
rect 36268 7225 36277 7259
rect 36277 7225 36311 7259
rect 36311 7225 36320 7259
rect 36268 7216 36320 7225
rect 38016 7216 38068 7268
rect 39028 7216 39080 7268
rect 31484 7148 31536 7200
rect 39856 7148 39908 7200
rect 40868 7148 40920 7200
rect 42156 7327 42208 7336
rect 42156 7293 42165 7327
rect 42165 7293 42199 7327
rect 42199 7293 42208 7327
rect 42156 7284 42208 7293
rect 43904 7420 43956 7472
rect 47400 7420 47452 7472
rect 45744 7352 45796 7404
rect 46388 7352 46440 7404
rect 44548 7259 44600 7268
rect 44548 7225 44557 7259
rect 44557 7225 44591 7259
rect 44591 7225 44600 7259
rect 44548 7216 44600 7225
rect 46204 7259 46256 7268
rect 41144 7148 41196 7200
rect 44364 7148 44416 7200
rect 46204 7225 46213 7259
rect 46213 7225 46247 7259
rect 46247 7225 46256 7259
rect 46204 7216 46256 7225
rect 46112 7148 46164 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 26700 6987 26752 6996
rect 26700 6953 26709 6987
rect 26709 6953 26743 6987
rect 26743 6953 26752 6987
rect 26700 6944 26752 6953
rect 29644 6944 29696 6996
rect 19892 6876 19944 6928
rect 21088 6919 21140 6928
rect 21088 6885 21097 6919
rect 21097 6885 21131 6919
rect 21131 6885 21140 6919
rect 21088 6876 21140 6885
rect 21640 6919 21692 6928
rect 21640 6885 21649 6919
rect 21649 6885 21683 6919
rect 21683 6885 21692 6919
rect 21640 6876 21692 6885
rect 23112 6876 23164 6928
rect 28172 6876 28224 6928
rect 29000 6919 29052 6928
rect 29000 6885 29009 6919
rect 29009 6885 29043 6919
rect 29043 6885 29052 6919
rect 29000 6876 29052 6885
rect 29184 6876 29236 6928
rect 32772 6944 32824 6996
rect 35256 6944 35308 6996
rect 35992 6944 36044 6996
rect 42156 6944 42208 6996
rect 42340 6944 42392 6996
rect 30104 6876 30156 6928
rect 30564 6876 30616 6928
rect 30932 6876 30984 6928
rect 34796 6876 34848 6928
rect 35440 6876 35492 6928
rect 35808 6876 35860 6928
rect 39028 6919 39080 6928
rect 39028 6885 39037 6919
rect 39037 6885 39071 6919
rect 39071 6885 39080 6919
rect 39028 6876 39080 6885
rect 39120 6919 39172 6928
rect 39120 6885 39129 6919
rect 39129 6885 39163 6919
rect 39163 6885 39172 6919
rect 39120 6876 39172 6885
rect 40224 6876 40276 6928
rect 40684 6919 40736 6928
rect 40684 6885 40693 6919
rect 40693 6885 40727 6919
rect 40727 6885 40736 6919
rect 43536 6919 43588 6928
rect 40684 6876 40736 6885
rect 43536 6885 43545 6919
rect 43545 6885 43579 6919
rect 43579 6885 43588 6919
rect 43536 6876 43588 6885
rect 44364 6876 44416 6928
rect 45192 6876 45244 6928
rect 46388 6876 46440 6928
rect 19432 6808 19484 6860
rect 24676 6808 24728 6860
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 32588 6808 32640 6860
rect 32956 6851 33008 6860
rect 32956 6817 32965 6851
rect 32965 6817 32999 6851
rect 32999 6817 33008 6851
rect 32956 6808 33008 6817
rect 33416 6808 33468 6860
rect 34612 6808 34664 6860
rect 35164 6808 35216 6860
rect 37740 6851 37792 6860
rect 37740 6817 37749 6851
rect 37749 6817 37783 6851
rect 37783 6817 37792 6851
rect 37740 6808 37792 6817
rect 42156 6808 42208 6860
rect 42708 6808 42760 6860
rect 46204 6851 46256 6860
rect 46204 6817 46213 6851
rect 46213 6817 46247 6851
rect 46247 6817 46256 6851
rect 46204 6808 46256 6817
rect 46296 6808 46348 6860
rect 21364 6740 21416 6792
rect 27988 6740 28040 6792
rect 27252 6672 27304 6724
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 22376 6647 22428 6656
rect 22376 6613 22385 6647
rect 22385 6613 22419 6647
rect 22419 6613 22428 6647
rect 22376 6604 22428 6613
rect 23388 6647 23440 6656
rect 23388 6613 23397 6647
rect 23397 6613 23431 6647
rect 23431 6613 23440 6647
rect 23388 6604 23440 6613
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 25320 6647 25372 6656
rect 25320 6613 25329 6647
rect 25329 6613 25363 6647
rect 25363 6613 25372 6647
rect 25320 6604 25372 6613
rect 25596 6647 25648 6656
rect 25596 6613 25605 6647
rect 25605 6613 25639 6647
rect 25639 6613 25648 6647
rect 25596 6604 25648 6613
rect 27160 6647 27212 6656
rect 27160 6613 27169 6647
rect 27169 6613 27203 6647
rect 27203 6613 27212 6647
rect 27160 6604 27212 6613
rect 28632 6647 28684 6656
rect 28632 6613 28641 6647
rect 28641 6613 28675 6647
rect 28675 6613 28684 6647
rect 31760 6740 31812 6792
rect 34704 6783 34756 6792
rect 34704 6749 34713 6783
rect 34713 6749 34747 6783
rect 34747 6749 34756 6783
rect 34704 6740 34756 6749
rect 36268 6783 36320 6792
rect 36268 6749 36277 6783
rect 36277 6749 36311 6783
rect 36311 6749 36320 6783
rect 36268 6740 36320 6749
rect 43444 6783 43496 6792
rect 28816 6672 28868 6724
rect 43444 6749 43453 6783
rect 43453 6749 43487 6783
rect 43487 6749 43496 6783
rect 43444 6740 43496 6749
rect 43904 6740 43956 6792
rect 42616 6672 42668 6724
rect 28632 6604 28684 6613
rect 33416 6604 33468 6656
rect 36268 6604 36320 6656
rect 38292 6604 38344 6656
rect 38476 6647 38528 6656
rect 38476 6613 38485 6647
rect 38485 6613 38519 6647
rect 38519 6613 38528 6647
rect 38476 6604 38528 6613
rect 41052 6604 41104 6656
rect 42340 6604 42392 6656
rect 44088 6604 44140 6656
rect 44548 6604 44600 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 19432 6400 19484 6452
rect 20352 6400 20404 6452
rect 21088 6400 21140 6452
rect 25412 6400 25464 6452
rect 28172 6400 28224 6452
rect 28448 6443 28500 6452
rect 28448 6409 28457 6443
rect 28457 6409 28491 6443
rect 28491 6409 28500 6443
rect 28448 6400 28500 6409
rect 29000 6400 29052 6452
rect 30288 6400 30340 6452
rect 31760 6443 31812 6452
rect 31760 6409 31769 6443
rect 31769 6409 31803 6443
rect 31803 6409 31812 6443
rect 31760 6400 31812 6409
rect 32956 6443 33008 6452
rect 32956 6409 32965 6443
rect 32965 6409 32999 6443
rect 32999 6409 33008 6443
rect 34612 6443 34664 6452
rect 32956 6400 33008 6409
rect 22468 6332 22520 6384
rect 22376 6264 22428 6316
rect 23756 6307 23808 6316
rect 23756 6273 23765 6307
rect 23765 6273 23799 6307
rect 23799 6273 23808 6307
rect 23756 6264 23808 6273
rect 24860 6264 24912 6316
rect 25320 6307 25372 6316
rect 25320 6273 25329 6307
rect 25329 6273 25363 6307
rect 25363 6273 25372 6307
rect 25320 6264 25372 6273
rect 27344 6332 27396 6384
rect 27988 6332 28040 6384
rect 28816 6332 28868 6384
rect 34612 6409 34621 6443
rect 34621 6409 34655 6443
rect 34655 6409 34664 6443
rect 34612 6400 34664 6409
rect 35624 6400 35676 6452
rect 38292 6443 38344 6452
rect 38292 6409 38301 6443
rect 38301 6409 38335 6443
rect 38335 6409 38344 6443
rect 38292 6400 38344 6409
rect 42156 6443 42208 6452
rect 42156 6409 42165 6443
rect 42165 6409 42199 6443
rect 42199 6409 42208 6443
rect 42156 6400 42208 6409
rect 42616 6443 42668 6452
rect 42616 6409 42625 6443
rect 42625 6409 42659 6443
rect 42659 6409 42668 6443
rect 42616 6400 42668 6409
rect 36084 6332 36136 6384
rect 37740 6375 37792 6384
rect 37740 6341 37749 6375
rect 37749 6341 37783 6375
rect 37783 6341 37792 6375
rect 37740 6332 37792 6341
rect 27160 6264 27212 6316
rect 27252 6307 27304 6316
rect 27252 6273 27261 6307
rect 27261 6273 27295 6307
rect 27295 6273 27304 6307
rect 27252 6264 27304 6273
rect 30472 6264 30524 6316
rect 19340 6196 19392 6248
rect 22100 6196 22152 6248
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 28448 6196 28500 6248
rect 30564 6239 30616 6248
rect 30564 6205 30573 6239
rect 30573 6205 30607 6239
rect 30607 6205 30616 6239
rect 30564 6196 30616 6205
rect 23940 6128 23992 6180
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 23112 6060 23164 6069
rect 24676 6103 24728 6112
rect 24676 6069 24685 6103
rect 24685 6069 24719 6103
rect 24719 6069 24728 6103
rect 24676 6060 24728 6069
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 26424 6128 26476 6180
rect 30288 6128 30340 6180
rect 33324 6264 33376 6316
rect 41052 6307 41104 6316
rect 41052 6273 41061 6307
rect 41061 6273 41095 6307
rect 41095 6273 41104 6307
rect 41052 6264 41104 6273
rect 41512 6307 41564 6316
rect 41512 6273 41521 6307
rect 41521 6273 41555 6307
rect 41555 6273 41564 6307
rect 41512 6264 41564 6273
rect 43444 6400 43496 6452
rect 45192 6443 45244 6452
rect 45192 6409 45201 6443
rect 45201 6409 45235 6443
rect 45235 6409 45244 6443
rect 45192 6400 45244 6409
rect 46296 6400 46348 6452
rect 43904 6307 43956 6316
rect 43904 6273 43913 6307
rect 43913 6273 43947 6307
rect 43947 6273 43956 6307
rect 43904 6264 43956 6273
rect 33416 6239 33468 6248
rect 33416 6205 33425 6239
rect 33425 6205 33459 6239
rect 33459 6205 33468 6239
rect 33416 6196 33468 6205
rect 35256 6196 35308 6248
rect 38292 6196 38344 6248
rect 38568 6196 38620 6248
rect 39120 6196 39172 6248
rect 44732 6239 44784 6248
rect 33968 6171 34020 6180
rect 33968 6137 33977 6171
rect 33977 6137 34011 6171
rect 34011 6137 34020 6171
rect 33968 6128 34020 6137
rect 36176 6171 36228 6180
rect 36176 6137 36185 6171
rect 36185 6137 36219 6171
rect 36219 6137 36228 6171
rect 36176 6128 36228 6137
rect 25136 6060 25188 6069
rect 29828 6060 29880 6112
rect 30104 6103 30156 6112
rect 30104 6069 30113 6103
rect 30113 6069 30147 6103
rect 30147 6069 30156 6103
rect 30104 6060 30156 6069
rect 31484 6103 31536 6112
rect 31484 6069 31493 6103
rect 31493 6069 31527 6103
rect 31527 6069 31536 6103
rect 31484 6060 31536 6069
rect 33416 6060 33468 6112
rect 35808 6060 35860 6112
rect 36452 6128 36504 6180
rect 36912 6128 36964 6180
rect 40132 6128 40184 6180
rect 44732 6205 44741 6239
rect 44741 6205 44775 6239
rect 44775 6205 44784 6239
rect 44732 6196 44784 6205
rect 46112 6196 46164 6248
rect 41696 6128 41748 6180
rect 41972 6128 42024 6180
rect 43444 6128 43496 6180
rect 43536 6128 43588 6180
rect 39764 6060 39816 6112
rect 40684 6060 40736 6112
rect 44732 6060 44784 6112
rect 45376 6060 45428 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 24676 5856 24728 5908
rect 27988 5899 28040 5908
rect 27988 5865 27997 5899
rect 27997 5865 28031 5899
rect 28031 5865 28040 5899
rect 27988 5856 28040 5865
rect 30564 5899 30616 5908
rect 30564 5865 30573 5899
rect 30573 5865 30607 5899
rect 30607 5865 30616 5899
rect 30564 5856 30616 5865
rect 31024 5856 31076 5908
rect 34796 5899 34848 5908
rect 34796 5865 34805 5899
rect 34805 5865 34839 5899
rect 34839 5865 34848 5899
rect 34796 5856 34848 5865
rect 35440 5856 35492 5908
rect 39028 5856 39080 5908
rect 39580 5856 39632 5908
rect 23112 5788 23164 5840
rect 24400 5788 24452 5840
rect 24860 5831 24912 5840
rect 24860 5797 24869 5831
rect 24869 5797 24903 5831
rect 24903 5797 24912 5831
rect 24860 5788 24912 5797
rect 27068 5788 27120 5840
rect 28172 5788 28224 5840
rect 28540 5788 28592 5840
rect 30288 5788 30340 5840
rect 21548 5720 21600 5772
rect 23388 5720 23440 5772
rect 30472 5763 30524 5772
rect 30472 5729 30481 5763
rect 30481 5729 30515 5763
rect 30515 5729 30524 5763
rect 30472 5720 30524 5729
rect 30840 5763 30892 5772
rect 30840 5729 30849 5763
rect 30849 5729 30883 5763
rect 30883 5729 30892 5763
rect 30840 5720 30892 5729
rect 32312 5720 32364 5772
rect 33048 5788 33100 5840
rect 38016 5788 38068 5840
rect 38936 5788 38988 5840
rect 40224 5856 40276 5908
rect 40868 5899 40920 5908
rect 40868 5865 40877 5899
rect 40877 5865 40911 5899
rect 40911 5865 40920 5899
rect 40868 5856 40920 5865
rect 41144 5856 41196 5908
rect 43904 5856 43956 5908
rect 46112 5899 46164 5908
rect 46112 5865 46121 5899
rect 46121 5865 46155 5899
rect 46155 5865 46164 5899
rect 46112 5856 46164 5865
rect 41880 5788 41932 5840
rect 43444 5788 43496 5840
rect 32680 5763 32732 5772
rect 32680 5729 32689 5763
rect 32689 5729 32723 5763
rect 32723 5729 32732 5763
rect 32680 5720 32732 5729
rect 33968 5720 34020 5772
rect 36360 5720 36412 5772
rect 45008 5763 45060 5772
rect 45008 5729 45017 5763
rect 45017 5729 45051 5763
rect 45051 5729 45060 5763
rect 45008 5720 45060 5729
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 24216 5695 24268 5704
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 27344 5695 27396 5704
rect 26332 5584 26384 5636
rect 27344 5661 27353 5695
rect 27353 5661 27387 5695
rect 27387 5661 27396 5695
rect 27344 5652 27396 5661
rect 28448 5652 28500 5704
rect 37464 5652 37516 5704
rect 39120 5652 39172 5704
rect 39304 5695 39356 5704
rect 39304 5661 39313 5695
rect 39313 5661 39347 5695
rect 39347 5661 39356 5695
rect 39304 5652 39356 5661
rect 40132 5652 40184 5704
rect 41512 5652 41564 5704
rect 43076 5652 43128 5704
rect 44088 5695 44140 5704
rect 44088 5661 44097 5695
rect 44097 5661 44131 5695
rect 44131 5661 44140 5695
rect 44088 5652 44140 5661
rect 29644 5584 29696 5636
rect 39028 5584 39080 5636
rect 39672 5584 39724 5636
rect 22468 5516 22520 5568
rect 23756 5559 23808 5568
rect 23756 5525 23765 5559
rect 23765 5525 23799 5559
rect 23799 5525 23808 5559
rect 23756 5516 23808 5525
rect 25320 5559 25372 5568
rect 25320 5525 25329 5559
rect 25329 5525 25363 5559
rect 25363 5525 25372 5559
rect 25320 5516 25372 5525
rect 26884 5559 26936 5568
rect 26884 5525 26893 5559
rect 26893 5525 26927 5559
rect 26927 5525 26936 5559
rect 26884 5516 26936 5525
rect 29460 5559 29512 5568
rect 29460 5525 29469 5559
rect 29469 5525 29503 5559
rect 29503 5525 29512 5559
rect 29460 5516 29512 5525
rect 33416 5516 33468 5568
rect 36820 5516 36872 5568
rect 37004 5559 37056 5568
rect 37004 5525 37013 5559
rect 37013 5525 37047 5559
rect 37047 5525 37056 5559
rect 37004 5516 37056 5525
rect 40224 5559 40276 5568
rect 40224 5525 40233 5559
rect 40233 5525 40267 5559
rect 40267 5525 40276 5559
rect 40224 5516 40276 5525
rect 43812 5516 43864 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 20352 5355 20404 5364
rect 20352 5321 20361 5355
rect 20361 5321 20395 5355
rect 20395 5321 20404 5355
rect 20352 5312 20404 5321
rect 21548 5355 21600 5364
rect 21548 5321 21557 5355
rect 21557 5321 21591 5355
rect 21591 5321 21600 5355
rect 21548 5312 21600 5321
rect 21916 5355 21968 5364
rect 21916 5321 21925 5355
rect 21925 5321 21959 5355
rect 21959 5321 21968 5355
rect 21916 5312 21968 5321
rect 23848 5312 23900 5364
rect 24400 5312 24452 5364
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 28172 5312 28224 5364
rect 28540 5355 28592 5364
rect 28540 5321 28549 5355
rect 28549 5321 28583 5355
rect 28583 5321 28592 5355
rect 28540 5312 28592 5321
rect 30472 5312 30524 5364
rect 32312 5355 32364 5364
rect 32312 5321 32321 5355
rect 32321 5321 32355 5355
rect 32355 5321 32364 5355
rect 32312 5312 32364 5321
rect 33968 5312 34020 5364
rect 36360 5355 36412 5364
rect 36360 5321 36369 5355
rect 36369 5321 36403 5355
rect 36403 5321 36412 5355
rect 36360 5312 36412 5321
rect 36452 5312 36504 5364
rect 37096 5312 37148 5364
rect 38016 5355 38068 5364
rect 38016 5321 38025 5355
rect 38025 5321 38059 5355
rect 38059 5321 38068 5355
rect 38016 5312 38068 5321
rect 38292 5355 38344 5364
rect 38292 5321 38301 5355
rect 38301 5321 38335 5355
rect 38335 5321 38344 5355
rect 38292 5312 38344 5321
rect 39580 5355 39632 5364
rect 39580 5321 39589 5355
rect 39589 5321 39623 5355
rect 39623 5321 39632 5355
rect 39580 5312 39632 5321
rect 40224 5312 40276 5364
rect 21364 5244 21416 5296
rect 20536 5219 20588 5228
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 21732 5176 21784 5228
rect 22376 5176 22428 5228
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 25320 5219 25372 5228
rect 24400 5176 24452 5185
rect 25320 5185 25329 5219
rect 25329 5185 25363 5219
rect 25363 5185 25372 5219
rect 25320 5176 25372 5185
rect 26884 5219 26936 5228
rect 26884 5185 26893 5219
rect 26893 5185 26927 5219
rect 26927 5185 26936 5219
rect 26884 5176 26936 5185
rect 21916 5108 21968 5160
rect 22100 5108 22152 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 34612 5244 34664 5296
rect 40684 5287 40736 5296
rect 40684 5253 40693 5287
rect 40693 5253 40727 5287
rect 40727 5253 40736 5287
rect 40684 5244 40736 5253
rect 40868 5244 40920 5296
rect 41512 5287 41564 5296
rect 31024 5219 31076 5228
rect 31024 5185 31033 5219
rect 31033 5185 31067 5219
rect 31067 5185 31076 5219
rect 31024 5176 31076 5185
rect 22468 5108 22520 5117
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 30840 5108 30892 5160
rect 33416 5176 33468 5228
rect 33600 5219 33652 5228
rect 33600 5185 33609 5219
rect 33609 5185 33643 5219
rect 33643 5185 33652 5219
rect 33600 5176 33652 5185
rect 34704 5176 34756 5228
rect 35532 5176 35584 5228
rect 37004 5219 37056 5228
rect 37004 5185 37013 5219
rect 37013 5185 37047 5219
rect 37047 5185 37056 5219
rect 37004 5176 37056 5185
rect 39304 5176 39356 5228
rect 40132 5176 40184 5228
rect 41512 5253 41521 5287
rect 41521 5253 41555 5287
rect 41555 5253 41564 5287
rect 41512 5244 41564 5253
rect 41880 5287 41932 5296
rect 41880 5253 41889 5287
rect 41889 5253 41923 5287
rect 41923 5253 41932 5287
rect 41880 5244 41932 5253
rect 20352 4972 20404 5024
rect 23112 5015 23164 5024
rect 23112 4981 23121 5015
rect 23121 4981 23155 5015
rect 23155 4981 23164 5015
rect 23112 4972 23164 4981
rect 23848 5083 23900 5092
rect 23848 5049 23857 5083
rect 23857 5049 23891 5083
rect 23891 5049 23900 5083
rect 25136 5083 25188 5092
rect 23848 5040 23900 5049
rect 25136 5049 25145 5083
rect 25145 5049 25179 5083
rect 25179 5049 25188 5083
rect 25136 5040 25188 5049
rect 27068 5040 27120 5092
rect 28448 5040 28500 5092
rect 24584 4972 24636 5024
rect 31024 5040 31076 5092
rect 33048 5040 33100 5092
rect 38292 5108 38344 5160
rect 39028 5151 39080 5160
rect 39028 5117 39037 5151
rect 39037 5117 39071 5151
rect 39071 5117 39080 5151
rect 39028 5108 39080 5117
rect 42340 5312 42392 5364
rect 43444 5355 43496 5364
rect 43444 5321 43453 5355
rect 43453 5321 43487 5355
rect 43487 5321 43496 5355
rect 43444 5312 43496 5321
rect 45008 5355 45060 5364
rect 45008 5321 45017 5355
rect 45017 5321 45051 5355
rect 45051 5321 45060 5355
rect 45008 5312 45060 5321
rect 43812 5219 43864 5228
rect 43812 5185 43821 5219
rect 43821 5185 43855 5219
rect 43855 5185 43864 5219
rect 43812 5176 43864 5185
rect 31944 5015 31996 5024
rect 31944 4981 31953 5015
rect 31953 4981 31987 5015
rect 31987 4981 31996 5015
rect 31944 4972 31996 4981
rect 33416 4972 33468 5024
rect 33692 4972 33744 5024
rect 34796 5040 34848 5092
rect 37096 5083 37148 5092
rect 37096 5049 37105 5083
rect 37105 5049 37139 5083
rect 37139 5049 37148 5083
rect 37096 5040 37148 5049
rect 37648 5083 37700 5092
rect 37648 5049 37657 5083
rect 37657 5049 37691 5083
rect 37691 5049 37700 5083
rect 37648 5040 37700 5049
rect 37740 5040 37792 5092
rect 40684 5040 40736 5092
rect 41604 5040 41656 5092
rect 43536 5040 43588 5092
rect 44456 5083 44508 5092
rect 44456 5049 44465 5083
rect 44465 5049 44499 5083
rect 44499 5049 44508 5083
rect 44456 5040 44508 5049
rect 36084 5015 36136 5024
rect 36084 4981 36093 5015
rect 36093 4981 36127 5015
rect 36127 4981 36136 5015
rect 36084 4972 36136 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 23664 4768 23716 4820
rect 24216 4768 24268 4820
rect 25964 4768 26016 4820
rect 27068 4768 27120 4820
rect 28264 4811 28316 4820
rect 28264 4777 28273 4811
rect 28273 4777 28307 4811
rect 28307 4777 28316 4811
rect 28264 4768 28316 4777
rect 29460 4768 29512 4820
rect 29828 4768 29880 4820
rect 31300 4768 31352 4820
rect 31760 4768 31812 4820
rect 32680 4811 32732 4820
rect 32680 4777 32689 4811
rect 32689 4777 32723 4811
rect 32723 4777 32732 4811
rect 32680 4768 32732 4777
rect 33048 4811 33100 4820
rect 33048 4777 33057 4811
rect 33057 4777 33091 4811
rect 33091 4777 33100 4811
rect 33048 4768 33100 4777
rect 35532 4811 35584 4820
rect 35532 4777 35541 4811
rect 35541 4777 35575 4811
rect 35575 4777 35584 4811
rect 35532 4768 35584 4777
rect 38844 4768 38896 4820
rect 43076 4811 43128 4820
rect 43076 4777 43085 4811
rect 43085 4777 43119 4811
rect 43119 4777 43128 4811
rect 43076 4768 43128 4777
rect 45008 4768 45060 4820
rect 23940 4700 23992 4752
rect 24400 4700 24452 4752
rect 24584 4743 24636 4752
rect 24584 4709 24593 4743
rect 24593 4709 24627 4743
rect 24627 4709 24636 4743
rect 24584 4700 24636 4709
rect 28448 4700 28500 4752
rect 30104 4700 30156 4752
rect 32588 4700 32640 4752
rect 33692 4700 33744 4752
rect 35716 4700 35768 4752
rect 36820 4700 36872 4752
rect 39488 4700 39540 4752
rect 39764 4743 39816 4752
rect 39764 4709 39773 4743
rect 39773 4709 39807 4743
rect 39807 4709 39816 4743
rect 39764 4700 39816 4709
rect 43444 4700 43496 4752
rect 44456 4700 44508 4752
rect 22928 4632 22980 4684
rect 25412 4675 25464 4684
rect 25412 4641 25421 4675
rect 25421 4641 25455 4675
rect 25455 4641 25464 4675
rect 25412 4632 25464 4641
rect 25596 4632 25648 4684
rect 26976 4632 27028 4684
rect 30656 4632 30708 4684
rect 31484 4632 31536 4684
rect 32128 4675 32180 4684
rect 32128 4641 32172 4675
rect 32172 4641 32180 4675
rect 38292 4675 38344 4684
rect 32128 4632 32180 4641
rect 38292 4641 38301 4675
rect 38301 4641 38335 4675
rect 38335 4641 38344 4675
rect 38292 4632 38344 4641
rect 23388 4564 23440 4616
rect 28080 4564 28132 4616
rect 29644 4564 29696 4616
rect 30840 4564 30892 4616
rect 32680 4564 32732 4616
rect 33600 4607 33652 4616
rect 33600 4573 33609 4607
rect 33609 4573 33643 4607
rect 33643 4573 33652 4607
rect 33600 4564 33652 4573
rect 35992 4564 36044 4616
rect 37648 4564 37700 4616
rect 37924 4496 37976 4548
rect 41328 4632 41380 4684
rect 42800 4632 42852 4684
rect 45376 4632 45428 4684
rect 38568 4607 38620 4616
rect 38568 4573 38577 4607
rect 38577 4573 38611 4607
rect 38611 4573 38620 4607
rect 38568 4564 38620 4573
rect 39120 4564 39172 4616
rect 43720 4607 43772 4616
rect 41788 4496 41840 4548
rect 43720 4573 43729 4607
rect 43729 4573 43763 4607
rect 43763 4573 43772 4607
rect 43720 4564 43772 4573
rect 43812 4496 43864 4548
rect 22468 4428 22520 4480
rect 34520 4471 34572 4480
rect 34520 4437 34529 4471
rect 34529 4437 34563 4471
rect 34563 4437 34572 4471
rect 34520 4428 34572 4437
rect 37464 4471 37516 4480
rect 37464 4437 37473 4471
rect 37473 4437 37507 4471
rect 37507 4437 37516 4471
rect 37464 4428 37516 4437
rect 40776 4471 40828 4480
rect 40776 4437 40785 4471
rect 40785 4437 40819 4471
rect 40819 4437 40828 4471
rect 40776 4428 40828 4437
rect 41696 4428 41748 4480
rect 41880 4471 41932 4480
rect 41880 4437 41889 4471
rect 41889 4437 41923 4471
rect 41923 4437 41932 4471
rect 41880 4428 41932 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 22928 4267 22980 4276
rect 22928 4233 22937 4267
rect 22937 4233 22971 4267
rect 22971 4233 22980 4267
rect 22928 4224 22980 4233
rect 25412 4267 25464 4276
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 26976 4267 27028 4276
rect 26976 4233 26985 4267
rect 26985 4233 27019 4267
rect 27019 4233 27028 4267
rect 26976 4224 27028 4233
rect 28632 4224 28684 4276
rect 29000 4267 29052 4276
rect 21732 4199 21784 4208
rect 21732 4165 21741 4199
rect 21741 4165 21775 4199
rect 21775 4165 21784 4199
rect 21732 4156 21784 4165
rect 23940 4199 23992 4208
rect 23940 4165 23949 4199
rect 23949 4165 23983 4199
rect 23983 4165 23992 4199
rect 23940 4156 23992 4165
rect 26148 4156 26200 4208
rect 29000 4233 29009 4267
rect 29009 4233 29043 4267
rect 29043 4233 29052 4267
rect 29000 4224 29052 4233
rect 29460 4224 29512 4276
rect 31300 4224 31352 4276
rect 32128 4267 32180 4276
rect 32128 4233 32137 4267
rect 32137 4233 32171 4267
rect 32171 4233 32180 4267
rect 32128 4224 32180 4233
rect 33600 4224 33652 4276
rect 37464 4224 37516 4276
rect 26424 4088 26476 4140
rect 28448 4088 28500 4140
rect 21732 4020 21784 4072
rect 22008 4020 22060 4072
rect 22468 4020 22520 4072
rect 24400 4063 24452 4072
rect 24400 4029 24409 4063
rect 24409 4029 24443 4063
rect 24443 4029 24452 4063
rect 24400 4020 24452 4029
rect 24492 4020 24544 4072
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 28356 4020 28408 4072
rect 22836 3952 22888 4004
rect 25136 3995 25188 4004
rect 25136 3961 25145 3995
rect 25145 3961 25179 3995
rect 25179 3961 25188 3995
rect 25136 3952 25188 3961
rect 26056 3995 26108 4004
rect 26056 3961 26065 3995
rect 26065 3961 26099 3995
rect 26099 3961 26108 3995
rect 26056 3952 26108 3961
rect 26148 3995 26200 4004
rect 26148 3961 26157 3995
rect 26157 3961 26191 3995
rect 26191 3961 26200 3995
rect 26148 3952 26200 3961
rect 26884 3952 26936 4004
rect 27160 3952 27212 4004
rect 29644 4131 29696 4140
rect 29644 4097 29653 4131
rect 29653 4097 29687 4131
rect 29687 4097 29696 4131
rect 29644 4088 29696 4097
rect 31024 4156 31076 4208
rect 33692 4199 33744 4208
rect 33692 4165 33701 4199
rect 33701 4165 33735 4199
rect 33735 4165 33744 4199
rect 33692 4156 33744 4165
rect 35716 4199 35768 4208
rect 35716 4165 35725 4199
rect 35725 4165 35759 4199
rect 35759 4165 35768 4199
rect 35716 4156 35768 4165
rect 36360 4156 36412 4208
rect 37924 4156 37976 4208
rect 38292 4224 38344 4276
rect 39488 4224 39540 4276
rect 41604 4267 41656 4276
rect 41604 4233 41613 4267
rect 41613 4233 41647 4267
rect 41647 4233 41656 4267
rect 41604 4224 41656 4233
rect 43444 4224 43496 4276
rect 39764 4156 39816 4208
rect 43996 4199 44048 4208
rect 43996 4165 44005 4199
rect 44005 4165 44039 4199
rect 44039 4165 44048 4199
rect 46204 4224 46256 4276
rect 45376 4199 45428 4208
rect 43996 4156 44048 4165
rect 45376 4165 45385 4199
rect 45385 4165 45419 4199
rect 45419 4165 45428 4199
rect 45376 4156 45428 4165
rect 42616 4088 42668 4140
rect 36084 4020 36136 4072
rect 36912 4063 36964 4072
rect 36912 4029 36921 4063
rect 36921 4029 36955 4063
rect 36955 4029 36964 4063
rect 36912 4020 36964 4029
rect 38292 4020 38344 4072
rect 38844 4020 38896 4072
rect 40776 4063 40828 4072
rect 40776 4029 40785 4063
rect 40785 4029 40819 4063
rect 40819 4029 40828 4063
rect 40776 4020 40828 4029
rect 45744 4063 45796 4072
rect 45744 4029 45753 4063
rect 45753 4029 45787 4063
rect 45787 4029 45796 4063
rect 45744 4020 45796 4029
rect 29368 3995 29420 4004
rect 29368 3961 29377 3995
rect 29377 3961 29411 3995
rect 29411 3961 29420 3995
rect 29368 3952 29420 3961
rect 29460 3995 29512 4004
rect 29460 3961 29469 3995
rect 29469 3961 29503 3995
rect 29503 3961 29512 3995
rect 29460 3952 29512 3961
rect 31208 3995 31260 4004
rect 31208 3961 31217 3995
rect 31217 3961 31251 3995
rect 31251 3961 31260 3995
rect 31208 3952 31260 3961
rect 31300 3995 31352 4004
rect 31300 3961 31309 3995
rect 31309 3961 31343 3995
rect 31343 3961 31352 3995
rect 32772 3995 32824 4004
rect 31300 3952 31352 3961
rect 32772 3961 32781 3995
rect 32781 3961 32815 3995
rect 32815 3961 32824 3995
rect 32772 3952 32824 3961
rect 36268 3995 36320 4004
rect 22560 3884 22612 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 28080 3927 28132 3936
rect 28080 3893 28089 3927
rect 28089 3893 28123 3927
rect 28123 3893 28132 3927
rect 28080 3884 28132 3893
rect 28448 3884 28500 3936
rect 32588 3927 32640 3936
rect 32588 3893 32597 3927
rect 32597 3893 32631 3927
rect 32631 3893 32640 3927
rect 36268 3961 36277 3995
rect 36277 3961 36311 3995
rect 36311 3961 36320 3995
rect 36268 3952 36320 3961
rect 36360 3995 36412 4004
rect 36360 3961 36369 3995
rect 36369 3961 36403 3995
rect 36403 3961 36412 3995
rect 39396 3995 39448 4004
rect 36360 3952 36412 3961
rect 39396 3961 39405 3995
rect 39405 3961 39439 3995
rect 39439 3961 39448 3995
rect 39396 3952 39448 3961
rect 41880 3995 41932 4004
rect 41880 3961 41889 3995
rect 41889 3961 41923 3995
rect 41923 3961 41932 3995
rect 41880 3952 41932 3961
rect 42524 3995 42576 4004
rect 32588 3884 32640 3893
rect 41052 3884 41104 3936
rect 41236 3927 41288 3936
rect 41236 3893 41245 3927
rect 41245 3893 41279 3927
rect 41279 3893 41288 3927
rect 41236 3884 41288 3893
rect 41604 3884 41656 3936
rect 42524 3961 42533 3995
rect 42533 3961 42567 3995
rect 42567 3961 42576 3995
rect 42524 3952 42576 3961
rect 43536 3995 43588 4004
rect 43536 3961 43545 3995
rect 43545 3961 43579 3995
rect 43579 3961 43588 3995
rect 43536 3952 43588 3961
rect 43904 3952 43956 4004
rect 42064 3884 42116 3936
rect 42800 3927 42852 3936
rect 42800 3893 42809 3927
rect 42809 3893 42843 3927
rect 42843 3893 42852 3927
rect 42800 3884 42852 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 22928 3680 22980 3732
rect 32772 3723 32824 3732
rect 32772 3689 32781 3723
rect 32781 3689 32815 3723
rect 32815 3689 32824 3723
rect 32772 3680 32824 3689
rect 36268 3680 36320 3732
rect 37832 3680 37884 3732
rect 23020 3612 23072 3664
rect 24584 3612 24636 3664
rect 26424 3612 26476 3664
rect 28632 3612 28684 3664
rect 30012 3612 30064 3664
rect 21364 3544 21416 3596
rect 24676 3587 24728 3596
rect 24676 3553 24685 3587
rect 24685 3553 24719 3587
rect 24719 3553 24728 3587
rect 24676 3544 24728 3553
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 29368 3587 29420 3596
rect 22836 3476 22888 3528
rect 24952 3476 25004 3528
rect 26608 3519 26660 3528
rect 26608 3485 26617 3519
rect 26617 3485 26651 3519
rect 26651 3485 26660 3519
rect 26608 3476 26660 3485
rect 26884 3519 26936 3528
rect 26884 3485 26893 3519
rect 26893 3485 26927 3519
rect 26927 3485 26936 3519
rect 26884 3476 26936 3485
rect 29368 3553 29377 3587
rect 29377 3553 29411 3587
rect 29411 3553 29420 3587
rect 29368 3544 29420 3553
rect 30288 3544 30340 3596
rect 30840 3587 30892 3596
rect 30840 3553 30849 3587
rect 30849 3553 30883 3587
rect 30883 3553 30892 3587
rect 30840 3544 30892 3553
rect 32036 3587 32088 3596
rect 32036 3553 32045 3587
rect 32045 3553 32079 3587
rect 32079 3553 32088 3587
rect 32036 3544 32088 3553
rect 33416 3587 33468 3596
rect 33416 3553 33425 3587
rect 33425 3553 33459 3587
rect 33459 3553 33468 3587
rect 33416 3544 33468 3553
rect 34612 3612 34664 3664
rect 37096 3655 37148 3664
rect 37096 3621 37105 3655
rect 37105 3621 37139 3655
rect 37139 3621 37148 3655
rect 37096 3612 37148 3621
rect 37556 3612 37608 3664
rect 38568 3680 38620 3732
rect 39396 3723 39448 3732
rect 35900 3544 35952 3596
rect 36544 3544 36596 3596
rect 38292 3587 38344 3596
rect 38292 3553 38301 3587
rect 38301 3553 38335 3587
rect 38335 3553 38344 3587
rect 38292 3544 38344 3553
rect 39396 3689 39405 3723
rect 39405 3689 39439 3723
rect 39439 3689 39448 3723
rect 39396 3680 39448 3689
rect 42800 3680 42852 3732
rect 43720 3680 43772 3732
rect 39580 3612 39632 3664
rect 39948 3612 40000 3664
rect 41788 3655 41840 3664
rect 41788 3621 41797 3655
rect 41797 3621 41831 3655
rect 41831 3621 41840 3655
rect 41788 3612 41840 3621
rect 41972 3612 42024 3664
rect 42524 3612 42576 3664
rect 40040 3544 40092 3596
rect 42616 3544 42668 3596
rect 30932 3519 30984 3528
rect 30932 3485 30941 3519
rect 30941 3485 30975 3519
rect 30975 3485 30984 3519
rect 30932 3476 30984 3485
rect 36084 3476 36136 3528
rect 39764 3476 39816 3528
rect 43628 3612 43680 3664
rect 43444 3519 43496 3528
rect 43444 3485 43453 3519
rect 43453 3485 43487 3519
rect 43487 3485 43496 3519
rect 43444 3476 43496 3485
rect 43996 3451 44048 3460
rect 43996 3417 44005 3451
rect 44005 3417 44039 3451
rect 44039 3417 44048 3451
rect 43996 3408 44048 3417
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 24032 3383 24084 3392
rect 24032 3349 24041 3383
rect 24041 3349 24075 3383
rect 24075 3349 24084 3383
rect 24032 3340 24084 3349
rect 24400 3340 24452 3392
rect 26056 3340 26108 3392
rect 27620 3383 27672 3392
rect 27620 3349 27629 3383
rect 27629 3349 27663 3383
rect 27663 3349 27672 3383
rect 27620 3340 27672 3349
rect 28172 3340 28224 3392
rect 29092 3383 29144 3392
rect 29092 3349 29101 3383
rect 29101 3349 29135 3383
rect 29135 3349 29144 3383
rect 29092 3340 29144 3349
rect 34704 3383 34756 3392
rect 34704 3349 34713 3383
rect 34713 3349 34747 3383
rect 34747 3349 34756 3383
rect 34704 3340 34756 3349
rect 35992 3340 36044 3392
rect 36176 3383 36228 3392
rect 36176 3349 36185 3383
rect 36185 3349 36219 3383
rect 36219 3349 36228 3383
rect 36176 3340 36228 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 22560 3136 22612 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 24400 3136 24452 3188
rect 24676 3136 24728 3188
rect 26424 3136 26476 3188
rect 26608 3136 26660 3188
rect 29092 3179 29144 3188
rect 29092 3145 29101 3179
rect 29101 3145 29135 3179
rect 29135 3145 29144 3179
rect 29092 3136 29144 3145
rect 30196 3136 30248 3188
rect 30840 3136 30892 3188
rect 32036 3136 32088 3188
rect 33692 3136 33744 3188
rect 34612 3179 34664 3188
rect 34612 3145 34621 3179
rect 34621 3145 34655 3179
rect 34655 3145 34664 3179
rect 34612 3136 34664 3145
rect 36544 3179 36596 3188
rect 36544 3145 36553 3179
rect 36553 3145 36587 3179
rect 36587 3145 36596 3179
rect 36544 3136 36596 3145
rect 41236 3136 41288 3188
rect 41972 3136 42024 3188
rect 42064 3179 42116 3188
rect 42064 3145 42073 3179
rect 42073 3145 42107 3179
rect 42107 3145 42116 3179
rect 42064 3136 42116 3145
rect 42432 3136 42484 3188
rect 43628 3179 43680 3188
rect 43628 3145 43637 3179
rect 43637 3145 43671 3179
rect 43671 3145 43680 3179
rect 43628 3136 43680 3145
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 28448 3068 28500 3120
rect 36084 3111 36136 3120
rect 24952 3043 25004 3052
rect 21364 3000 21416 3009
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 30932 3000 30984 3052
rect 22560 2932 22612 2984
rect 24032 2975 24084 2984
rect 24032 2941 24050 2975
rect 24050 2941 24084 2975
rect 24032 2932 24084 2941
rect 25044 2932 25096 2984
rect 27620 2932 27672 2984
rect 28264 2932 28316 2984
rect 29092 2932 29144 2984
rect 23112 2864 23164 2916
rect 24768 2864 24820 2916
rect 23388 2839 23440 2848
rect 23388 2805 23397 2839
rect 23397 2805 23431 2839
rect 23431 2805 23440 2839
rect 23388 2796 23440 2805
rect 25872 2839 25924 2848
rect 25872 2805 25881 2839
rect 25881 2805 25915 2839
rect 25915 2805 25924 2839
rect 25872 2796 25924 2805
rect 28356 2864 28408 2916
rect 28724 2864 28776 2916
rect 33416 2975 33468 2984
rect 33416 2941 33425 2975
rect 33425 2941 33459 2975
rect 33459 2941 33468 2975
rect 33416 2932 33468 2941
rect 36084 3077 36093 3111
rect 36093 3077 36127 3111
rect 36127 3077 36136 3111
rect 36084 3068 36136 3077
rect 39948 3111 40000 3120
rect 39948 3077 39957 3111
rect 39957 3077 39991 3111
rect 39991 3077 40000 3111
rect 39948 3068 40000 3077
rect 34336 2932 34388 2984
rect 34704 2932 34756 2984
rect 38292 3000 38344 3052
rect 39396 3000 39448 3052
rect 39764 3000 39816 3052
rect 40500 3043 40552 3052
rect 40500 3009 40509 3043
rect 40509 3009 40543 3043
rect 40543 3009 40552 3043
rect 40500 3000 40552 3009
rect 37556 2975 37608 2984
rect 37556 2941 37565 2975
rect 37565 2941 37599 2975
rect 37599 2941 37608 2975
rect 37556 2932 37608 2941
rect 28632 2839 28684 2848
rect 28632 2805 28641 2839
rect 28641 2805 28675 2839
rect 28675 2805 28684 2839
rect 31024 2864 31076 2916
rect 35072 2864 35124 2916
rect 37832 2907 37884 2916
rect 37832 2873 37841 2907
rect 37841 2873 37875 2907
rect 37875 2873 37884 2907
rect 37832 2864 37884 2873
rect 39948 2864 40000 2916
rect 41696 3000 41748 3052
rect 42340 3043 42392 3052
rect 42340 3009 42349 3043
rect 42349 3009 42383 3043
rect 42383 3009 42392 3043
rect 42340 3000 42392 3009
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 43904 3043 43956 3052
rect 43904 3009 43913 3043
rect 43913 3009 43947 3043
rect 43947 3009 43956 3043
rect 43904 3000 43956 3009
rect 44088 3000 44140 3052
rect 42064 2932 42116 2984
rect 42432 2907 42484 2916
rect 42432 2873 42441 2907
rect 42441 2873 42475 2907
rect 42475 2873 42484 2907
rect 42432 2864 42484 2873
rect 30288 2839 30340 2848
rect 28632 2796 28684 2805
rect 30288 2805 30297 2839
rect 30297 2805 30331 2839
rect 30331 2805 30340 2839
rect 30288 2796 30340 2805
rect 34612 2796 34664 2848
rect 38660 2796 38712 2848
rect 43628 2796 43680 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 21456 2592 21508 2644
rect 22836 2635 22888 2644
rect 22836 2601 22845 2635
rect 22845 2601 22879 2635
rect 22879 2601 22888 2635
rect 22836 2592 22888 2601
rect 24860 2592 24912 2644
rect 25044 2592 25096 2644
rect 26608 2592 26660 2644
rect 28172 2635 28224 2644
rect 28172 2601 28181 2635
rect 28181 2601 28215 2635
rect 28215 2601 28224 2635
rect 28172 2592 28224 2601
rect 28264 2592 28316 2644
rect 30932 2592 30984 2644
rect 31208 2592 31260 2644
rect 36176 2592 36228 2644
rect 37004 2592 37056 2644
rect 37832 2592 37884 2644
rect 22560 2567 22612 2576
rect 22560 2533 22569 2567
rect 22569 2533 22603 2567
rect 22603 2533 22612 2567
rect 22560 2524 22612 2533
rect 23388 2524 23440 2576
rect 24768 2567 24820 2576
rect 24768 2533 24777 2567
rect 24777 2533 24811 2567
rect 24811 2533 24820 2567
rect 24768 2524 24820 2533
rect 22008 2388 22060 2440
rect 25136 2456 25188 2508
rect 25872 2456 25924 2508
rect 28356 2499 28408 2508
rect 28356 2465 28365 2499
rect 28365 2465 28399 2499
rect 28399 2465 28408 2499
rect 28356 2456 28408 2465
rect 34336 2567 34388 2576
rect 34336 2533 34345 2567
rect 34345 2533 34379 2567
rect 34379 2533 34388 2567
rect 34336 2524 34388 2533
rect 34612 2524 34664 2576
rect 35992 2524 36044 2576
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 30196 2499 30248 2508
rect 30196 2465 30205 2499
rect 30205 2465 30239 2499
rect 30239 2465 30248 2499
rect 30196 2456 30248 2465
rect 31944 2456 31996 2508
rect 33416 2456 33468 2508
rect 34428 2456 34480 2508
rect 35072 2456 35124 2508
rect 38660 2635 38712 2644
rect 38660 2601 38669 2635
rect 38669 2601 38703 2635
rect 38703 2601 38712 2635
rect 40040 2635 40092 2644
rect 38660 2592 38712 2601
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 40500 2635 40552 2644
rect 40500 2601 40509 2635
rect 40509 2601 40543 2635
rect 40543 2601 40552 2635
rect 40500 2592 40552 2601
rect 41052 2592 41104 2644
rect 41972 2524 42024 2576
rect 43444 2524 43496 2576
rect 40776 2456 40828 2508
rect 42064 2388 42116 2440
rect 41880 2320 41932 2372
rect 30288 2252 30340 2304
rect 34428 2252 34480 2304
rect 42340 2252 42392 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 6182 49586 6238 50000
rect 6104 49558 6238 49586
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 6104 44169 6132 49558
rect 6182 49520 6238 49558
rect 18602 49586 18658 50000
rect 31114 49586 31170 50000
rect 43626 49586 43682 50000
rect 18602 49558 18920 49586
rect 18602 49520 18658 49558
rect 18892 45626 18920 49558
rect 31114 49558 31340 49586
rect 31114 49520 31170 49558
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 28172 46368 28224 46374
rect 28172 46310 28224 46316
rect 28448 46368 28500 46374
rect 28448 46310 28500 46316
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 25320 45824 25372 45830
rect 25320 45766 25372 45772
rect 18880 45620 18932 45626
rect 18880 45562 18932 45568
rect 21548 45620 21600 45626
rect 21548 45562 21600 45568
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 21560 44402 21588 45562
rect 22282 45384 22338 45393
rect 25332 45354 25360 45766
rect 22282 45319 22338 45328
rect 25320 45348 25372 45354
rect 22296 44538 22324 45319
rect 25320 45290 25372 45296
rect 25412 45348 25464 45354
rect 25412 45290 25464 45296
rect 27712 45348 27764 45354
rect 27712 45290 27764 45296
rect 25136 45280 25188 45286
rect 25136 45222 25188 45228
rect 25148 45014 25176 45222
rect 25136 45008 25188 45014
rect 25136 44950 25188 44956
rect 23848 44940 23900 44946
rect 23848 44882 23900 44888
rect 22284 44532 22336 44538
rect 22284 44474 22336 44480
rect 21548 44396 21600 44402
rect 21548 44338 21600 44344
rect 19156 44328 19208 44334
rect 19156 44270 19208 44276
rect 6090 44160 6146 44169
rect 6090 44095 6146 44104
rect 19062 44160 19118 44169
rect 19062 44095 19118 44104
rect 18052 43716 18104 43722
rect 18052 43658 18104 43664
rect 16488 43648 16540 43654
rect 16488 43590 16540 43596
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 16500 43314 16528 43590
rect 18064 43382 18092 43658
rect 18052 43376 18104 43382
rect 18052 43318 18104 43324
rect 16488 43308 16540 43314
rect 16488 43250 16540 43256
rect 17224 43308 17276 43314
rect 17224 43250 17276 43256
rect 16500 42906 16528 43250
rect 16580 43172 16632 43178
rect 16580 43114 16632 43120
rect 16488 42900 16540 42906
rect 16488 42842 16540 42848
rect 16592 42838 16620 43114
rect 16304 42832 16356 42838
rect 16304 42774 16356 42780
rect 16580 42832 16632 42838
rect 16580 42774 16632 42780
rect 15936 42764 15988 42770
rect 15936 42706 15988 42712
rect 15948 42566 15976 42706
rect 16212 42696 16264 42702
rect 16212 42638 16264 42644
rect 15936 42560 15988 42566
rect 15936 42502 15988 42508
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 15568 42152 15620 42158
rect 15568 42094 15620 42100
rect 14924 42016 14976 42022
rect 14924 41958 14976 41964
rect 14936 41585 14964 41958
rect 14922 41576 14978 41585
rect 14922 41511 14978 41520
rect 15384 41540 15436 41546
rect 13912 41472 13964 41478
rect 13912 41414 13964 41420
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 13924 38962 13952 41414
rect 14004 40928 14056 40934
rect 14004 40870 14056 40876
rect 13912 38956 13964 38962
rect 13912 38898 13964 38904
rect 13636 38888 13688 38894
rect 13636 38830 13688 38836
rect 13820 38888 13872 38894
rect 13820 38830 13872 38836
rect 13544 38752 13596 38758
rect 13544 38694 13596 38700
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 13268 35760 13320 35766
rect 13268 35702 13320 35708
rect 13280 35630 13308 35702
rect 13268 35624 13320 35630
rect 13268 35566 13320 35572
rect 13280 34950 13308 35566
rect 13268 34944 13320 34950
rect 13268 34886 13320 34892
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 13280 30802 13308 34886
rect 13556 34542 13584 38694
rect 13648 36242 13676 38830
rect 13832 38486 13860 38830
rect 13820 38480 13872 38486
rect 13820 38422 13872 38428
rect 14016 37330 14044 40870
rect 14004 37324 14056 37330
rect 14004 37266 14056 37272
rect 14016 36582 14044 37266
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14004 36576 14056 36582
rect 14004 36518 14056 36524
rect 13636 36236 13688 36242
rect 13636 36178 13688 36184
rect 13648 34950 13676 36178
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13636 34944 13688 34950
rect 13636 34886 13688 34892
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13556 34202 13584 34478
rect 13360 34196 13412 34202
rect 13360 34138 13412 34144
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 12728 30054 12756 30738
rect 13280 30394 13308 30738
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 12728 29753 12756 29990
rect 12714 29744 12770 29753
rect 12714 29679 12770 29688
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 13096 28762 13124 29990
rect 13372 29306 13400 34138
rect 13648 32978 13676 34886
rect 13832 34542 13860 35566
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13832 33590 13860 34478
rect 13820 33584 13872 33590
rect 13820 33526 13872 33532
rect 13820 33040 13872 33046
rect 13820 32982 13872 32988
rect 13636 32972 13688 32978
rect 13636 32914 13688 32920
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13372 29102 13400 29242
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 13372 27334 13400 29038
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 13556 25809 13584 32302
rect 13648 32230 13676 32914
rect 13832 32570 13860 32982
rect 13912 32972 13964 32978
rect 13912 32914 13964 32920
rect 13820 32564 13872 32570
rect 13820 32506 13872 32512
rect 13820 32428 13872 32434
rect 13924 32416 13952 32914
rect 14016 32570 14044 36518
rect 14568 36310 14596 36654
rect 14648 36644 14700 36650
rect 14648 36586 14700 36592
rect 14556 36304 14608 36310
rect 14556 36246 14608 36252
rect 14188 36236 14240 36242
rect 14188 36178 14240 36184
rect 14200 35698 14228 36178
rect 14660 35834 14688 36586
rect 14936 36242 14964 41511
rect 15384 41482 15436 41488
rect 15396 40934 15424 41482
rect 15580 41478 15608 42094
rect 15568 41472 15620 41478
rect 15568 41414 15620 41420
rect 15384 40928 15436 40934
rect 15384 40870 15436 40876
rect 15948 40633 15976 42502
rect 16224 42362 16252 42638
rect 16316 42362 16344 42774
rect 17132 42628 17184 42634
rect 17132 42570 17184 42576
rect 16212 42356 16264 42362
rect 16212 42298 16264 42304
rect 16304 42356 16356 42362
rect 16304 42298 16356 42304
rect 16672 42356 16724 42362
rect 16672 42298 16724 42304
rect 16212 42084 16264 42090
rect 16212 42026 16264 42032
rect 16224 40662 16252 42026
rect 16684 41750 16712 42298
rect 16672 41744 16724 41750
rect 16672 41686 16724 41692
rect 16684 41274 16712 41686
rect 16672 41268 16724 41274
rect 16672 41210 16724 41216
rect 17144 41138 17172 42570
rect 17236 41750 17264 43250
rect 17224 41744 17276 41750
rect 17224 41686 17276 41692
rect 17132 41132 17184 41138
rect 17132 41074 17184 41080
rect 16396 40928 16448 40934
rect 16396 40870 16448 40876
rect 16408 40730 16436 40870
rect 17144 40730 17172 41074
rect 16396 40724 16448 40730
rect 16396 40666 16448 40672
rect 17132 40724 17184 40730
rect 17132 40666 17184 40672
rect 16212 40656 16264 40662
rect 15934 40624 15990 40633
rect 16212 40598 16264 40604
rect 15934 40559 15990 40568
rect 15292 40520 15344 40526
rect 15292 40462 15344 40468
rect 15304 39846 15332 40462
rect 15292 39840 15344 39846
rect 15292 39782 15344 39788
rect 15304 38962 15332 39782
rect 15292 38956 15344 38962
rect 15292 38898 15344 38904
rect 15752 38752 15804 38758
rect 15752 38694 15804 38700
rect 15568 38480 15620 38486
rect 15568 38422 15620 38428
rect 15200 37800 15252 37806
rect 15200 37742 15252 37748
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14660 35562 14688 35770
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14648 35556 14700 35562
rect 14648 35498 14700 35504
rect 14660 34746 14688 35498
rect 14752 35290 14780 35566
rect 14936 35494 14964 36178
rect 14924 35488 14976 35494
rect 14924 35430 14976 35436
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14648 34740 14700 34746
rect 14648 34682 14700 34688
rect 14660 34474 14688 34682
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14648 34468 14700 34474
rect 14648 34410 14700 34416
rect 14660 33658 14688 34410
rect 14844 34202 14872 34478
rect 14832 34196 14884 34202
rect 14832 34138 14884 34144
rect 14648 33652 14700 33658
rect 14648 33594 14700 33600
rect 14660 33134 14688 33594
rect 14740 33448 14792 33454
rect 14740 33390 14792 33396
rect 14568 33106 14688 33134
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 14384 32434 14412 32846
rect 14568 32570 14596 33106
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 13872 32388 13952 32416
rect 14372 32428 14424 32434
rect 13820 32370 13872 32376
rect 14372 32370 14424 32376
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13648 28014 13676 32166
rect 13728 31816 13780 31822
rect 13728 31758 13780 31764
rect 13740 31482 13768 31758
rect 13728 31476 13780 31482
rect 13728 31418 13780 31424
rect 13832 30784 13860 32370
rect 14384 32026 14412 32370
rect 14568 32298 14596 32506
rect 14556 32292 14608 32298
rect 14556 32234 14608 32240
rect 14372 32020 14424 32026
rect 14372 31962 14424 31968
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 13912 30796 13964 30802
rect 13832 30756 13912 30784
rect 13912 30738 13964 30744
rect 13924 29714 13952 30738
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 13912 29708 13964 29714
rect 13832 29668 13912 29696
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13740 28762 13768 29582
rect 13832 29102 13860 29668
rect 13912 29650 13964 29656
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13832 28694 13860 29038
rect 13820 28688 13872 28694
rect 13820 28630 13872 28636
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 13728 27940 13780 27946
rect 13728 27882 13780 27888
rect 13740 27130 13768 27882
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 14108 26518 14136 29990
rect 14384 29850 14412 31758
rect 14568 30870 14596 32234
rect 14752 32026 14780 33390
rect 14740 32020 14792 32026
rect 14740 31962 14792 31968
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14556 29776 14608 29782
rect 14660 29764 14688 31622
rect 14740 31136 14792 31142
rect 14936 31124 14964 35430
rect 15212 31346 15240 37742
rect 15476 37732 15528 37738
rect 15476 37674 15528 37680
rect 15292 37664 15344 37670
rect 15292 37606 15344 37612
rect 15304 37398 15332 37606
rect 15292 37392 15344 37398
rect 15292 37334 15344 37340
rect 15304 36378 15332 37334
rect 15384 37120 15436 37126
rect 15384 37062 15436 37068
rect 15396 36786 15424 37062
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15488 36378 15516 37674
rect 15580 37466 15608 38422
rect 15660 38412 15712 38418
rect 15660 38354 15712 38360
rect 15672 38010 15700 38354
rect 15660 38004 15712 38010
rect 15660 37946 15712 37952
rect 15568 37460 15620 37466
rect 15568 37402 15620 37408
rect 15292 36372 15344 36378
rect 15292 36314 15344 36320
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15672 34202 15700 37946
rect 15764 35766 15792 38694
rect 15948 37942 15976 40559
rect 16120 40384 16172 40390
rect 16120 40326 16172 40332
rect 16132 39982 16160 40326
rect 16120 39976 16172 39982
rect 16120 39918 16172 39924
rect 16132 38486 16160 39918
rect 16224 39914 16252 40598
rect 17236 40508 17264 41686
rect 17408 41608 17460 41614
rect 17408 41550 17460 41556
rect 17420 41274 17448 41550
rect 17408 41268 17460 41274
rect 17408 41210 17460 41216
rect 17960 40996 18012 41002
rect 17960 40938 18012 40944
rect 17408 40656 17460 40662
rect 17408 40598 17460 40604
rect 17316 40520 17368 40526
rect 17236 40480 17316 40508
rect 17316 40462 17368 40468
rect 17328 40118 17356 40462
rect 17420 40186 17448 40598
rect 17972 40526 18000 40938
rect 17960 40520 18012 40526
rect 17960 40462 18012 40468
rect 17408 40180 17460 40186
rect 17408 40122 17460 40128
rect 17316 40112 17368 40118
rect 17316 40054 17368 40060
rect 16212 39908 16264 39914
rect 16212 39850 16264 39856
rect 16224 39574 16252 39850
rect 17960 39636 18012 39642
rect 17960 39578 18012 39584
rect 16212 39568 16264 39574
rect 16212 39510 16264 39516
rect 16224 39098 16252 39510
rect 16764 39432 16816 39438
rect 16764 39374 16816 39380
rect 16212 39092 16264 39098
rect 16212 39034 16264 39040
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16500 38554 16528 38830
rect 16776 38758 16804 39374
rect 16764 38752 16816 38758
rect 16764 38694 16816 38700
rect 16776 38554 16804 38694
rect 17972 38554 18000 39578
rect 18064 39574 18092 43318
rect 18972 43172 19024 43178
rect 18972 43114 19024 43120
rect 18420 43104 18472 43110
rect 18420 43046 18472 43052
rect 18604 43104 18656 43110
rect 18604 43046 18656 43052
rect 18880 43104 18932 43110
rect 18880 43046 18932 43052
rect 18432 42906 18460 43046
rect 18420 42900 18472 42906
rect 18420 42842 18472 42848
rect 18616 42129 18644 43046
rect 18892 42838 18920 43046
rect 18984 42906 19012 43114
rect 19076 42945 19104 44095
rect 19168 43790 19196 44270
rect 21364 44260 21416 44266
rect 21364 44202 21416 44208
rect 19248 44192 19300 44198
rect 19248 44134 19300 44140
rect 19156 43784 19208 43790
rect 19260 43761 19288 44134
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19340 43920 19392 43926
rect 19340 43862 19392 43868
rect 19156 43726 19208 43732
rect 19246 43752 19302 43761
rect 19168 43450 19196 43726
rect 19246 43687 19302 43696
rect 19156 43444 19208 43450
rect 19156 43386 19208 43392
rect 19352 43092 19380 43862
rect 19306 43064 19380 43092
rect 21180 43104 21232 43110
rect 19062 42936 19118 42945
rect 18972 42900 19024 42906
rect 19306 42922 19334 43064
rect 21180 43046 21232 43052
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19062 42871 19118 42880
rect 19260 42894 19334 42922
rect 19430 42936 19486 42945
rect 18972 42842 19024 42848
rect 18880 42832 18932 42838
rect 18880 42774 18932 42780
rect 18972 42764 19024 42770
rect 18972 42706 19024 42712
rect 18602 42120 18658 42129
rect 18524 42078 18602 42106
rect 18144 40724 18196 40730
rect 18144 40666 18196 40672
rect 18052 39568 18104 39574
rect 18052 39510 18104 39516
rect 18064 39098 18092 39510
rect 18052 39092 18104 39098
rect 18052 39034 18104 39040
rect 18052 38820 18104 38826
rect 18052 38762 18104 38768
rect 16488 38548 16540 38554
rect 16488 38490 16540 38496
rect 16764 38548 16816 38554
rect 16764 38490 16816 38496
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 16120 38480 16172 38486
rect 16120 38422 16172 38428
rect 17868 38412 17920 38418
rect 17868 38354 17920 38360
rect 17040 38208 17092 38214
rect 17040 38150 17092 38156
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 15936 37936 15988 37942
rect 15936 37878 15988 37884
rect 16580 37936 16632 37942
rect 16580 37878 16632 37884
rect 16120 37732 16172 37738
rect 16120 37674 16172 37680
rect 16132 37398 16160 37674
rect 16120 37392 16172 37398
rect 16120 37334 16172 37340
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15844 35760 15896 35766
rect 15844 35702 15896 35708
rect 15856 35290 15884 35702
rect 15844 35284 15896 35290
rect 15844 35226 15896 35232
rect 16040 35154 16068 37062
rect 16132 36922 16160 37334
rect 16396 37188 16448 37194
rect 16396 37130 16448 37136
rect 16120 36916 16172 36922
rect 16120 36858 16172 36864
rect 16132 36582 16160 36858
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 16132 36378 16160 36518
rect 16120 36372 16172 36378
rect 16120 36314 16172 36320
rect 16408 36174 16436 37130
rect 16592 36582 16620 37878
rect 17052 37670 17080 38150
rect 17040 37664 17092 37670
rect 17040 37606 17092 37612
rect 17788 37398 17816 38150
rect 17880 37738 17908 38354
rect 18064 38010 18092 38762
rect 18052 38004 18104 38010
rect 18052 37946 18104 37952
rect 17868 37732 17920 37738
rect 17868 37674 17920 37680
rect 17776 37392 17828 37398
rect 17776 37334 17828 37340
rect 17684 36848 17736 36854
rect 17684 36790 17736 36796
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 16488 36304 16540 36310
rect 16488 36246 16540 36252
rect 16396 36168 16448 36174
rect 16396 36110 16448 36116
rect 16408 35290 16436 36110
rect 16500 35834 16528 36246
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 16488 35216 16540 35222
rect 16488 35158 16540 35164
rect 16028 35148 16080 35154
rect 16028 35090 16080 35096
rect 16040 34678 16068 35090
rect 16500 34746 16528 35158
rect 16592 35086 16620 36518
rect 16684 35834 16712 36722
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 17052 35086 17080 36110
rect 17500 35624 17552 35630
rect 17498 35592 17500 35601
rect 17552 35592 17554 35601
rect 17498 35527 17554 35536
rect 17512 35494 17540 35527
rect 17500 35488 17552 35494
rect 17500 35430 17552 35436
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 17040 35080 17092 35086
rect 17040 35022 17092 35028
rect 16592 34746 16620 35022
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 16488 34740 16540 34746
rect 16488 34682 16540 34688
rect 16580 34740 16632 34746
rect 16580 34682 16632 34688
rect 16028 34672 16080 34678
rect 16028 34614 16080 34620
rect 16396 34672 16448 34678
rect 16396 34614 16448 34620
rect 16408 34202 16436 34614
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 16396 34196 16448 34202
rect 16396 34138 16448 34144
rect 15672 33454 15700 34138
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16040 33522 16068 33934
rect 16408 33658 16436 34138
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16028 33516 16080 33522
rect 16028 33458 16080 33464
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15660 33448 15712 33454
rect 15660 33390 15712 33396
rect 15304 31686 15332 33390
rect 15384 33040 15436 33046
rect 15384 32982 15436 32988
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15396 32570 15424 32982
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15580 32502 15608 32982
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 15568 32496 15620 32502
rect 15568 32438 15620 32444
rect 15580 31958 15608 32438
rect 15568 31952 15620 31958
rect 15856 31929 15884 32846
rect 16408 32502 16436 33594
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 16868 32570 16896 33322
rect 17236 33046 17264 34886
rect 17512 33658 17540 35430
rect 17696 34134 17724 36790
rect 17788 36378 17816 37334
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17880 36242 17908 37674
rect 18052 37664 18104 37670
rect 18156 37652 18184 40666
rect 18104 37624 18184 37652
rect 18420 37664 18472 37670
rect 18052 37606 18104 37612
rect 18420 37606 18472 37612
rect 17960 37392 18012 37398
rect 17960 37334 18012 37340
rect 17972 36650 18000 37334
rect 17960 36644 18012 36650
rect 17960 36586 18012 36592
rect 17868 36236 17920 36242
rect 17868 36178 17920 36184
rect 17880 34950 17908 36178
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 18064 34542 18092 37606
rect 18432 37466 18460 37606
rect 18420 37460 18472 37466
rect 18420 37402 18472 37408
rect 18432 36786 18460 37402
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18524 36564 18552 42078
rect 18602 42055 18658 42064
rect 18984 42022 19012 42706
rect 18972 42016 19024 42022
rect 18972 41958 19024 41964
rect 18696 41744 18748 41750
rect 18696 41686 18748 41692
rect 18708 41274 18736 41686
rect 18880 41608 18932 41614
rect 18880 41550 18932 41556
rect 18696 41268 18748 41274
rect 18696 41210 18748 41216
rect 18892 40934 18920 41550
rect 18880 40928 18932 40934
rect 18880 40870 18932 40876
rect 18604 40588 18656 40594
rect 18604 40530 18656 40536
rect 18616 40186 18644 40530
rect 18696 40520 18748 40526
rect 18696 40462 18748 40468
rect 18604 40180 18656 40186
rect 18604 40122 18656 40128
rect 18616 39098 18644 40122
rect 18708 39574 18736 40462
rect 18696 39568 18748 39574
rect 18696 39510 18748 39516
rect 18604 39092 18656 39098
rect 18604 39034 18656 39040
rect 18788 38888 18840 38894
rect 18788 38830 18840 38836
rect 18696 37936 18748 37942
rect 18696 37878 18748 37884
rect 18524 36536 18644 36564
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 18432 35766 18460 36178
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18420 35760 18472 35766
rect 18420 35702 18472 35708
rect 18420 35488 18472 35494
rect 18420 35430 18472 35436
rect 18432 34610 18460 35430
rect 18524 35154 18552 36110
rect 18616 35834 18644 36536
rect 18604 35828 18656 35834
rect 18604 35770 18656 35776
rect 18616 35630 18644 35770
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18512 35148 18564 35154
rect 18512 35090 18564 35096
rect 18524 34746 18552 35090
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18616 34785 18644 35022
rect 18602 34776 18658 34785
rect 18512 34740 18564 34746
rect 18602 34711 18658 34720
rect 18512 34682 18564 34688
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 18064 34202 18092 34478
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18512 34400 18564 34406
rect 18512 34342 18564 34348
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17684 34128 17736 34134
rect 17684 34070 17736 34076
rect 17960 34128 18012 34134
rect 17960 34070 18012 34076
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17512 33454 17540 33594
rect 17500 33448 17552 33454
rect 17500 33390 17552 33396
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17224 33040 17276 33046
rect 17224 32982 17276 32988
rect 17132 32972 17184 32978
rect 17132 32914 17184 32920
rect 16856 32564 16908 32570
rect 16856 32506 16908 32512
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 16868 32366 16896 32506
rect 16856 32360 16908 32366
rect 16856 32302 16908 32308
rect 17144 32230 17172 32914
rect 17236 32881 17264 32982
rect 17222 32872 17278 32881
rect 17222 32807 17278 32816
rect 17236 32570 17264 32807
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 16396 32224 16448 32230
rect 16396 32166 16448 32172
rect 17132 32224 17184 32230
rect 17132 32166 17184 32172
rect 15568 31894 15620 31900
rect 15842 31920 15898 31929
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15396 31482 15424 31758
rect 15580 31482 15608 31894
rect 15842 31855 15898 31864
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15016 31340 15068 31346
rect 15016 31282 15068 31288
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 14792 31096 14964 31124
rect 14740 31078 14792 31084
rect 14608 29736 14688 29764
rect 14556 29718 14608 29724
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14384 29170 14412 29582
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 14568 28966 14596 29718
rect 14752 29696 14780 31078
rect 14660 29668 14780 29696
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 14370 28656 14426 28665
rect 14370 28591 14426 28600
rect 14384 28558 14412 28591
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 28218 14412 28494
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 14200 26790 14228 27474
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 26926 14412 27270
rect 14372 26920 14424 26926
rect 14372 26862 14424 26868
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 13542 25800 13598 25809
rect 13542 25735 13598 25744
rect 14200 25265 14228 26726
rect 14384 26246 14412 26862
rect 14372 26240 14424 26246
rect 14372 26182 14424 26188
rect 14384 26081 14412 26182
rect 14370 26072 14426 26081
rect 14370 26007 14426 26016
rect 14186 25256 14242 25265
rect 14186 25191 14242 25200
rect 14278 25120 14334 25129
rect 4220 25052 4516 25072
rect 14278 25055 14334 25064
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 14108 23866 14136 24142
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14108 23769 14136 23802
rect 14094 23760 14150 23769
rect 14094 23695 14150 23704
rect 14292 23633 14320 25055
rect 14476 23730 14504 27814
rect 14568 27538 14596 28902
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14660 24041 14688 29668
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14752 26926 14780 27066
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14752 26586 14780 26862
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 14844 25906 14872 26930
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14844 25498 14872 25842
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 14936 24954 14964 25298
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14646 24032 14702 24041
rect 14646 23967 14702 23976
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14278 23624 14334 23633
rect 14278 23559 14334 23568
rect 14292 23186 14320 23559
rect 14476 23322 14504 23666
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 14292 22778 14320 23122
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14660 22574 14688 23967
rect 15028 23474 15056 31282
rect 15396 30938 15424 31418
rect 15672 31346 15700 31690
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15304 30394 15332 30806
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15108 30388 15160 30394
rect 15108 30330 15160 30336
rect 15292 30388 15344 30394
rect 15292 30330 15344 30336
rect 15120 26926 15148 30330
rect 15304 29782 15332 30330
rect 15488 30122 15516 30534
rect 15476 30116 15528 30122
rect 15476 30058 15528 30064
rect 15752 30116 15804 30122
rect 15752 30058 15804 30064
rect 15488 29850 15516 30058
rect 15764 29850 15792 30058
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15292 29776 15344 29782
rect 15212 29736 15292 29764
rect 15212 29306 15240 29736
rect 15292 29718 15344 29724
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15212 28966 15240 29242
rect 15304 29102 15332 29582
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15200 28960 15252 28966
rect 15200 28902 15252 28908
rect 15304 28762 15332 29038
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15856 28558 15884 31855
rect 16304 31680 16356 31686
rect 16304 31622 16356 31628
rect 16120 31204 16172 31210
rect 16316 31192 16344 31622
rect 16172 31164 16344 31192
rect 16120 31146 16172 31152
rect 16316 30938 16344 31164
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15948 28694 15976 28902
rect 16408 28762 16436 32166
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16868 31414 16896 31826
rect 16856 31408 16908 31414
rect 16856 31350 16908 31356
rect 16488 31204 16540 31210
rect 16488 31146 16540 31152
rect 16500 30122 16528 31146
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16592 30394 16620 30670
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16500 29578 16528 30058
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16396 28756 16448 28762
rect 16396 28698 16448 28704
rect 15936 28688 15988 28694
rect 15936 28630 15988 28636
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15488 28218 15516 28494
rect 15948 28218 15976 28630
rect 16500 28558 16528 29514
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 15384 27668 15436 27674
rect 15384 27610 15436 27616
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15396 26450 15424 27610
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15764 26790 15792 27474
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16118 27024 16174 27033
rect 16118 26959 16174 26968
rect 16132 26926 16160 26959
rect 16408 26926 16436 27406
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15568 26512 15620 26518
rect 15488 26472 15568 26500
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15396 26042 15424 26386
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15488 25702 15516 26472
rect 15568 26454 15620 26460
rect 15764 25945 15792 26726
rect 15750 25936 15806 25945
rect 15750 25871 15806 25880
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15488 25430 15516 25638
rect 15764 25498 15792 25638
rect 15752 25492 15804 25498
rect 15752 25434 15804 25440
rect 15476 25424 15528 25430
rect 15476 25366 15528 25372
rect 15488 24614 15516 25366
rect 15948 25362 15976 26726
rect 16408 26586 16436 26862
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16212 25492 16264 25498
rect 16212 25434 16264 25440
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 16132 24682 16160 25162
rect 16224 24682 16252 25434
rect 16408 25430 16436 26182
rect 16396 25424 16448 25430
rect 16396 25366 16448 25372
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16120 24676 16172 24682
rect 16120 24618 16172 24624
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 15488 23594 15516 24550
rect 16040 24138 16068 24550
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15200 23520 15252 23526
rect 15028 23468 15200 23474
rect 15028 23462 15252 23468
rect 15028 23446 15240 23462
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 15212 22098 15240 23446
rect 15856 23254 15884 23598
rect 16132 23254 16160 24618
rect 16316 24342 16344 25094
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16316 23866 16344 24278
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16500 23474 16528 28494
rect 16592 26926 16620 29990
rect 16960 29850 16988 29990
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 17236 29238 17264 32506
rect 17328 31346 17356 33254
rect 17972 33114 18000 34070
rect 18064 33522 18092 34138
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 18156 32978 18184 34342
rect 18524 34105 18552 34342
rect 18616 34134 18644 34711
rect 18604 34128 18656 34134
rect 18510 34096 18566 34105
rect 18604 34070 18656 34076
rect 18510 34031 18566 34040
rect 18604 33448 18656 33454
rect 18708 33436 18736 37878
rect 18800 36174 18828 38830
rect 18892 38486 18920 40870
rect 18984 40497 19012 41958
rect 19076 40730 19104 42871
rect 19260 42838 19288 42894
rect 19580 42928 19876 42948
rect 19430 42871 19486 42880
rect 19444 42838 19472 42871
rect 21192 42838 21220 43046
rect 19248 42832 19300 42838
rect 19432 42832 19484 42838
rect 19300 42780 19380 42794
rect 19248 42774 19380 42780
rect 19432 42774 19484 42780
rect 21180 42832 21232 42838
rect 21180 42774 21232 42780
rect 19260 42766 19380 42774
rect 21376 42770 21404 44202
rect 19156 42696 19208 42702
rect 19156 42638 19208 42644
rect 19168 42362 19196 42638
rect 19156 42356 19208 42362
rect 19156 42298 19208 42304
rect 19352 42022 19380 42766
rect 21364 42764 21416 42770
rect 21364 42706 21416 42712
rect 21376 42362 21404 42706
rect 21364 42356 21416 42362
rect 21364 42298 21416 42304
rect 21560 42158 21588 44338
rect 22296 44334 22324 44474
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22008 44192 22060 44198
rect 22008 44134 22060 44140
rect 21916 43784 21968 43790
rect 21916 43726 21968 43732
rect 21928 43382 21956 43726
rect 21916 43376 21968 43382
rect 21916 43318 21968 43324
rect 21732 43172 21784 43178
rect 21732 43114 21784 43120
rect 21744 42566 21772 43114
rect 21928 42906 21956 43318
rect 21916 42900 21968 42906
rect 21916 42842 21968 42848
rect 21824 42832 21876 42838
rect 21824 42774 21876 42780
rect 21732 42560 21784 42566
rect 21732 42502 21784 42508
rect 21744 42294 21772 42502
rect 21836 42294 21864 42774
rect 21732 42288 21784 42294
rect 21732 42230 21784 42236
rect 21824 42288 21876 42294
rect 21824 42230 21876 42236
rect 22020 42226 22048 44134
rect 22100 43920 22152 43926
rect 22100 43862 22152 43868
rect 22112 43178 22140 43862
rect 22100 43172 22152 43178
rect 22100 43114 22152 43120
rect 22112 42838 22140 43114
rect 22100 42832 22152 42838
rect 22100 42774 22152 42780
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 20168 42152 20220 42158
rect 20168 42094 20220 42100
rect 21548 42152 21600 42158
rect 21548 42094 21600 42100
rect 19892 42084 19944 42090
rect 19892 42026 19944 42032
rect 19340 42016 19392 42022
rect 19340 41958 19392 41964
rect 19352 41818 19380 41958
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19904 41138 19932 42026
rect 19892 41132 19944 41138
rect 19892 41074 19944 41080
rect 19432 40996 19484 41002
rect 19432 40938 19484 40944
rect 19064 40724 19116 40730
rect 19064 40666 19116 40672
rect 18970 40488 19026 40497
rect 18970 40423 19026 40432
rect 19156 40384 19208 40390
rect 19156 40326 19208 40332
rect 19064 39976 19116 39982
rect 19064 39918 19116 39924
rect 19076 39302 19104 39918
rect 19064 39296 19116 39302
rect 19064 39238 19116 39244
rect 19076 38962 19104 39238
rect 19064 38956 19116 38962
rect 19064 38898 19116 38904
rect 19168 38894 19196 40326
rect 19444 40186 19472 40938
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19904 40662 19932 41074
rect 19892 40656 19944 40662
rect 19892 40598 19944 40604
rect 19432 40180 19484 40186
rect 19432 40122 19484 40128
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19616 39500 19668 39506
rect 19616 39442 19668 39448
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 19156 38888 19208 38894
rect 19156 38830 19208 38836
rect 18880 38480 18932 38486
rect 18880 38422 18932 38428
rect 19168 38418 19196 38830
rect 19444 38554 19472 39238
rect 19628 38894 19656 39442
rect 19616 38888 19668 38894
rect 19616 38830 19668 38836
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19432 38548 19484 38554
rect 19432 38490 19484 38496
rect 19156 38412 19208 38418
rect 19156 38354 19208 38360
rect 19444 37874 19472 38490
rect 20180 38010 20208 42094
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 20536 40996 20588 41002
rect 20536 40938 20588 40944
rect 20260 39976 20312 39982
rect 20260 39918 20312 39924
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 19432 37868 19484 37874
rect 19432 37810 19484 37816
rect 19892 37868 19944 37874
rect 19892 37810 19944 37816
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19444 37398 19472 37606
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19432 37392 19484 37398
rect 19432 37334 19484 37340
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19352 36922 19380 37198
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19352 36378 19380 36858
rect 19444 36854 19472 37334
rect 19616 37256 19668 37262
rect 19616 37198 19668 37204
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19628 36786 19656 37198
rect 19904 37194 19932 37810
rect 19892 37188 19944 37194
rect 19892 37130 19944 37136
rect 19904 36904 19932 37130
rect 19904 36876 20024 36904
rect 19616 36780 19668 36786
rect 19616 36722 19668 36728
rect 19892 36780 19944 36786
rect 19892 36722 19944 36728
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 18788 36168 18840 36174
rect 18788 36110 18840 36116
rect 19248 36032 19300 36038
rect 19248 35974 19300 35980
rect 19260 35698 19288 35974
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19340 35556 19392 35562
rect 19340 35498 19392 35504
rect 18972 35488 19024 35494
rect 18972 35430 19024 35436
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18892 34678 18920 35226
rect 18880 34672 18932 34678
rect 18880 34614 18932 34620
rect 18656 33408 18736 33436
rect 18604 33390 18656 33396
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18064 32434 18092 32846
rect 18616 32774 18644 33390
rect 18984 33289 19012 35430
rect 19352 34950 19380 35498
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19352 34474 19380 34886
rect 19904 34610 19932 36722
rect 19996 35698 20024 36876
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 19076 34202 19104 34342
rect 19352 34202 19380 34410
rect 19444 34202 19472 34546
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19064 34196 19116 34202
rect 19064 34138 19116 34144
rect 19340 34196 19392 34202
rect 19340 34138 19392 34144
rect 19432 34196 19484 34202
rect 19432 34138 19484 34144
rect 19076 33697 19104 34138
rect 20180 34066 20208 37946
rect 20272 36242 20300 39918
rect 20548 39506 20576 40938
rect 21192 40934 21220 41550
rect 21284 41206 21312 41754
rect 22020 41750 22048 42162
rect 22112 42090 22140 42774
rect 22100 42084 22152 42090
rect 22100 42026 22152 42032
rect 22112 41818 22140 42026
rect 22100 41812 22152 41818
rect 22100 41754 22152 41760
rect 22008 41744 22060 41750
rect 22008 41686 22060 41692
rect 22192 41268 22244 41274
rect 22192 41210 22244 41216
rect 21272 41200 21324 41206
rect 21272 41142 21324 41148
rect 22204 41002 22232 41210
rect 21732 40996 21784 41002
rect 21732 40938 21784 40944
rect 22192 40996 22244 41002
rect 22192 40938 22244 40944
rect 21180 40928 21232 40934
rect 21180 40870 21232 40876
rect 20628 39908 20680 39914
rect 20628 39850 20680 39856
rect 20640 39574 20668 39850
rect 20628 39568 20680 39574
rect 20628 39510 20680 39516
rect 20536 39500 20588 39506
rect 20536 39442 20588 39448
rect 21088 39296 21140 39302
rect 21088 39238 21140 39244
rect 20352 38752 20404 38758
rect 20352 38694 20404 38700
rect 20260 36236 20312 36242
rect 20260 36178 20312 36184
rect 20272 35834 20300 36178
rect 20260 35828 20312 35834
rect 20260 35770 20312 35776
rect 20272 34610 20300 35770
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 19800 33856 19852 33862
rect 19800 33798 19852 33804
rect 19062 33688 19118 33697
rect 19062 33623 19118 33632
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19064 33380 19116 33386
rect 19064 33322 19116 33328
rect 18970 33280 19026 33289
rect 18970 33215 19026 33224
rect 18970 33144 19026 33153
rect 18892 33106 18970 33134
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 18234 31920 18290 31929
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17316 31340 17368 31346
rect 17316 31282 17368 31288
rect 17696 30938 17724 31758
rect 18064 31482 18092 31894
rect 18234 31855 18290 31864
rect 18248 31822 18276 31855
rect 18892 31822 18920 33106
rect 18970 33079 19026 33088
rect 19076 32910 19104 33322
rect 19340 33040 19392 33046
rect 19340 32982 19392 32988
rect 19064 32904 19116 32910
rect 19064 32846 19116 32852
rect 19076 32570 19104 32846
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18972 32224 19024 32230
rect 18972 32166 19024 32172
rect 18984 31958 19012 32166
rect 18972 31952 19024 31958
rect 18972 31894 19024 31900
rect 18236 31816 18288 31822
rect 18236 31758 18288 31764
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 18052 31476 18104 31482
rect 18052 31418 18104 31424
rect 18064 31142 18092 31418
rect 18800 31278 18828 31622
rect 18788 31272 18840 31278
rect 18788 31214 18840 31220
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 18064 30870 18092 31078
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 18064 30394 18092 30806
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 18432 30394 18460 30602
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 18420 30388 18472 30394
rect 18420 30330 18472 30336
rect 18064 30104 18092 30330
rect 18236 30116 18288 30122
rect 18064 30076 18236 30104
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17788 29850 17816 29990
rect 18064 29850 18092 30076
rect 18236 30058 18288 30064
rect 18788 30116 18840 30122
rect 18788 30058 18840 30064
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18420 29776 18472 29782
rect 18420 29718 18472 29724
rect 18432 29306 18460 29718
rect 18800 29646 18828 30058
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 16672 29232 16724 29238
rect 16672 29174 16724 29180
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 16684 28014 16712 29174
rect 18052 29096 18104 29102
rect 18052 29038 18104 29044
rect 17592 28960 17644 28966
rect 17592 28902 17644 28908
rect 17224 28620 17276 28626
rect 17224 28562 17276 28568
rect 17236 28422 17264 28562
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16684 27674 16712 27950
rect 17132 27940 17184 27946
rect 17132 27882 17184 27888
rect 16672 27668 16724 27674
rect 16672 27610 16724 27616
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 17144 26586 17172 27882
rect 17236 27878 17264 28358
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 17236 27538 17264 27814
rect 17512 27538 17540 27950
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17236 26994 17264 27474
rect 17512 27130 17540 27474
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26897 17264 26930
rect 17222 26888 17278 26897
rect 17222 26823 17278 26832
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17236 25770 17264 26386
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17132 25424 17184 25430
rect 17132 25366 17184 25372
rect 17144 24954 17172 25366
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 16764 24880 16816 24886
rect 16764 24822 16816 24828
rect 16776 24342 16804 24822
rect 16764 24336 16816 24342
rect 16764 24278 16816 24284
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17052 23798 17080 24142
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16408 23446 16528 23474
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15672 22506 15700 22918
rect 15856 22778 15884 23190
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 15856 22488 15884 22714
rect 16132 22642 16160 23054
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 15936 22500 15988 22506
rect 15856 22460 15936 22488
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 15212 21350 15240 22034
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 3790 2000 3846 2009
rect 3790 1935 3846 1944
rect 3514 82 3570 480
rect 3804 82 3832 1935
rect 3514 54 3832 82
rect 10598 82 10654 480
rect 10980 82 11008 9386
rect 13832 8945 13860 21286
rect 15304 21146 15332 22374
rect 15856 22234 15884 22460
rect 15936 22442 15988 22448
rect 16132 22234 16160 22578
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 16408 13814 16436 23446
rect 16684 22982 16712 23666
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22166 16712 22918
rect 17236 22681 17264 25706
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17328 25430 17356 25638
rect 17316 25424 17368 25430
rect 17316 25366 17368 25372
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17420 24954 17448 25230
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17604 23905 17632 28902
rect 18064 28694 18092 29038
rect 18432 28762 18460 29242
rect 18800 29238 18828 29582
rect 18892 29560 18920 31758
rect 18972 29572 19024 29578
rect 18892 29532 18972 29560
rect 18972 29514 19024 29520
rect 18788 29232 18840 29238
rect 18788 29174 18840 29180
rect 18420 28756 18472 28762
rect 18420 28698 18472 28704
rect 19156 28756 19208 28762
rect 19156 28698 19208 28704
rect 18052 28688 18104 28694
rect 18052 28630 18104 28636
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 28218 17816 28562
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 18248 27538 18276 27814
rect 19168 27538 19196 28698
rect 19260 28626 19288 32710
rect 19352 32298 19380 32982
rect 19340 32292 19392 32298
rect 19340 32234 19392 32240
rect 19444 31890 19472 33594
rect 19812 33454 19840 33798
rect 20180 33658 20208 34002
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 20088 33386 20116 33458
rect 20272 33402 20300 34546
rect 20364 34406 20392 38694
rect 20536 38412 20588 38418
rect 20536 38354 20588 38360
rect 20904 38412 20956 38418
rect 20904 38354 20956 38360
rect 20548 37670 20576 38354
rect 20720 38208 20772 38214
rect 20720 38150 20772 38156
rect 20536 37664 20588 37670
rect 20536 37606 20588 37612
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20076 33380 20128 33386
rect 20076 33322 20128 33328
rect 20180 33374 20300 33402
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 20088 32978 20116 33322
rect 19892 32972 19944 32978
rect 19892 32914 19944 32920
rect 20076 32972 20128 32978
rect 20076 32914 20128 32920
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19904 31958 19932 32914
rect 20180 32858 20208 33374
rect 20260 33312 20312 33318
rect 20260 33254 20312 33260
rect 20088 32830 20208 32858
rect 19892 31952 19944 31958
rect 19892 31894 19944 31900
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19430 31512 19486 31521
rect 19904 31482 19932 31894
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19430 31447 19486 31456
rect 19892 31476 19944 31482
rect 19444 31414 19472 31447
rect 19892 31418 19944 31424
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19260 28529 19288 28562
rect 19246 28520 19302 28529
rect 19246 28455 19302 28464
rect 19260 28150 19288 28455
rect 19352 28218 19380 28562
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 19156 27532 19208 27538
rect 19156 27474 19208 27480
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18064 26994 18092 27406
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 17788 25838 17816 26726
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17972 25974 18000 26182
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 18064 25906 18092 26522
rect 18880 26512 18932 26518
rect 18984 26500 19012 26726
rect 19168 26586 19196 27474
rect 19352 26858 19380 27542
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 18932 26472 19012 26500
rect 18880 26454 18932 26460
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18432 26042 18460 26318
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17590 23896 17646 23905
rect 17590 23831 17646 23840
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17512 22778 17540 23530
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17222 22672 17278 22681
rect 17144 22630 17222 22658
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 21457 16528 21490
rect 16486 21448 16542 21457
rect 16486 21383 16542 21392
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16960 20534 16988 20810
rect 17144 20602 17172 22630
rect 17222 22607 17278 22616
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21350 17264 22034
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 21146 17264 21286
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17512 20602 17540 20878
rect 17788 20602 17816 25774
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17880 24886 17908 25298
rect 18432 25294 18460 25978
rect 18524 25362 18552 26318
rect 18984 26042 19012 26472
rect 18972 26036 19024 26042
rect 18972 25978 19024 25984
rect 18972 25696 19024 25702
rect 18972 25638 19024 25644
rect 18984 25430 19012 25638
rect 18696 25424 18748 25430
rect 18696 25366 18748 25372
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 18432 24682 18460 25094
rect 18708 24954 18736 25366
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18616 24818 18644 24890
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 24410 18184 24550
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17880 23866 17908 24210
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 18156 23730 18184 24006
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18156 23474 18184 23666
rect 18248 23594 18276 24346
rect 18236 23588 18288 23594
rect 18288 23548 18368 23576
rect 18236 23530 18288 23536
rect 18156 23446 18276 23474
rect 18248 23118 18276 23446
rect 18340 23254 18368 23548
rect 18328 23248 18380 23254
rect 18328 23190 18380 23196
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17972 21690 18000 22442
rect 18156 22234 18184 23054
rect 18340 22506 18368 23190
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 18156 21350 18184 22034
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18064 20942 18092 21286
rect 18892 21010 18920 24822
rect 18984 24410 19012 25366
rect 19444 25362 19472 31350
rect 19996 31142 20024 31826
rect 20088 31192 20116 32830
rect 20272 32774 20300 33254
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20272 32026 20300 32710
rect 20364 32366 20392 34342
rect 20548 32502 20576 37606
rect 20732 36786 20760 38150
rect 20916 37942 20944 38354
rect 20904 37936 20956 37942
rect 20904 37878 20956 37884
rect 20916 37466 20944 37878
rect 20904 37460 20956 37466
rect 20904 37402 20956 37408
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 21008 36922 21036 37198
rect 20996 36916 21048 36922
rect 20996 36858 21048 36864
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20732 36378 20760 36722
rect 20812 36644 20864 36650
rect 20812 36586 20864 36592
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20824 36310 20852 36586
rect 20812 36304 20864 36310
rect 20812 36246 20864 36252
rect 20628 35556 20680 35562
rect 20628 35498 20680 35504
rect 20640 34950 20668 35498
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20640 34746 20668 34886
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20640 34406 20668 34682
rect 20812 34468 20864 34474
rect 20812 34410 20864 34416
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20824 34202 20852 34410
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 20732 33318 20760 34002
rect 20720 33312 20772 33318
rect 20640 33272 20720 33300
rect 20640 32774 20668 33272
rect 20720 33254 20772 33260
rect 21100 33134 21128 39238
rect 21192 38554 21220 40870
rect 21744 40730 21772 40938
rect 22204 40730 22232 40938
rect 21732 40724 21784 40730
rect 21732 40666 21784 40672
rect 22192 40724 22244 40730
rect 22192 40666 22244 40672
rect 21548 40588 21600 40594
rect 21548 40530 21600 40536
rect 21560 39846 21588 40530
rect 22204 39914 22232 40666
rect 22192 39908 22244 39914
rect 22192 39850 22244 39856
rect 21548 39840 21600 39846
rect 21548 39782 21600 39788
rect 22204 39642 22232 39850
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22008 39568 22060 39574
rect 22008 39510 22060 39516
rect 21456 39432 21508 39438
rect 21456 39374 21508 39380
rect 21364 39364 21416 39370
rect 21364 39306 21416 39312
rect 21376 38894 21404 39306
rect 21468 38962 21496 39374
rect 22020 39030 22048 39510
rect 22008 39024 22060 39030
rect 22008 38966 22060 38972
rect 21456 38956 21508 38962
rect 21456 38898 21508 38904
rect 21364 38888 21416 38894
rect 21364 38830 21416 38836
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 21376 38418 21404 38830
rect 22008 38820 22060 38826
rect 22008 38762 22060 38768
rect 21364 38412 21416 38418
rect 21364 38354 21416 38360
rect 21376 38010 21404 38354
rect 21364 38004 21416 38010
rect 21364 37946 21416 37952
rect 22020 37806 22048 38762
rect 22296 38554 22324 44270
rect 23860 44266 23888 44882
rect 24952 44872 25004 44878
rect 24952 44814 25004 44820
rect 24964 44538 24992 44814
rect 24952 44532 25004 44538
rect 24952 44474 25004 44480
rect 23848 44260 23900 44266
rect 23848 44202 23900 44208
rect 25228 44260 25280 44266
rect 25228 44202 25280 44208
rect 25240 43926 25268 44202
rect 25332 43994 25360 45290
rect 25424 45014 25452 45290
rect 27620 45280 27672 45286
rect 27620 45222 27672 45228
rect 27632 45082 27660 45222
rect 27620 45076 27672 45082
rect 27620 45018 27672 45024
rect 25412 45008 25464 45014
rect 25412 44950 25464 44956
rect 25424 44266 25452 44950
rect 27068 44940 27120 44946
rect 27068 44882 27120 44888
rect 25872 44872 25924 44878
rect 25872 44814 25924 44820
rect 25688 44396 25740 44402
rect 25688 44338 25740 44344
rect 25412 44260 25464 44266
rect 25412 44202 25464 44208
rect 25424 43994 25452 44202
rect 25320 43988 25372 43994
rect 25320 43930 25372 43936
rect 25412 43988 25464 43994
rect 25412 43930 25464 43936
rect 25228 43920 25280 43926
rect 25228 43862 25280 43868
rect 24768 43852 24820 43858
rect 24768 43794 24820 43800
rect 25320 43852 25372 43858
rect 25320 43794 25372 43800
rect 23388 43784 23440 43790
rect 23388 43726 23440 43732
rect 22376 43308 22428 43314
rect 22376 43250 22428 43256
rect 22388 40118 22416 43250
rect 22928 43104 22980 43110
rect 22928 43046 22980 43052
rect 22940 42838 22968 43046
rect 22928 42832 22980 42838
rect 22928 42774 22980 42780
rect 22560 42628 22612 42634
rect 22560 42570 22612 42576
rect 22572 41138 22600 42570
rect 22940 42362 22968 42774
rect 22928 42356 22980 42362
rect 22928 42298 22980 42304
rect 22652 42084 22704 42090
rect 22652 42026 22704 42032
rect 22560 41132 22612 41138
rect 22560 41074 22612 41080
rect 22468 40996 22520 41002
rect 22468 40938 22520 40944
rect 22480 40186 22508 40938
rect 22664 40662 22692 42026
rect 23400 41750 23428 43726
rect 24780 43450 24808 43794
rect 24768 43444 24820 43450
rect 24768 43386 24820 43392
rect 24768 43172 24820 43178
rect 24768 43114 24820 43120
rect 24216 43104 24268 43110
rect 24216 43046 24268 43052
rect 24492 43104 24544 43110
rect 24492 43046 24544 43052
rect 23848 42764 23900 42770
rect 23848 42706 23900 42712
rect 23860 42022 23888 42706
rect 24228 42702 24256 43046
rect 24216 42696 24268 42702
rect 24216 42638 24268 42644
rect 23848 42016 23900 42022
rect 23848 41958 23900 41964
rect 22836 41744 22888 41750
rect 22836 41686 22888 41692
rect 23388 41744 23440 41750
rect 23388 41686 23440 41692
rect 22848 41274 22876 41686
rect 23388 41608 23440 41614
rect 23388 41550 23440 41556
rect 22836 41268 22888 41274
rect 22836 41210 22888 41216
rect 22652 40656 22704 40662
rect 22652 40598 22704 40604
rect 22744 40520 22796 40526
rect 22744 40462 22796 40468
rect 22468 40180 22520 40186
rect 22468 40122 22520 40128
rect 22376 40112 22428 40118
rect 22376 40054 22428 40060
rect 22652 39840 22704 39846
rect 22652 39782 22704 39788
rect 22284 38548 22336 38554
rect 22284 38490 22336 38496
rect 22008 37800 22060 37806
rect 22008 37742 22060 37748
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21732 37392 21784 37398
rect 21732 37334 21784 37340
rect 21364 37256 21416 37262
rect 21364 37198 21416 37204
rect 21376 36650 21404 37198
rect 21744 36650 21772 37334
rect 21836 37126 21864 37606
rect 22020 37126 22048 37742
rect 21824 37120 21876 37126
rect 21824 37062 21876 37068
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 21836 36854 21864 37062
rect 21824 36848 21876 36854
rect 21824 36790 21876 36796
rect 21364 36644 21416 36650
rect 21364 36586 21416 36592
rect 21732 36644 21784 36650
rect 21732 36586 21784 36592
rect 21272 36032 21324 36038
rect 21272 35974 21324 35980
rect 21284 35698 21312 35974
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 21284 35290 21312 35634
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21376 34678 21404 36586
rect 21732 36236 21784 36242
rect 21732 36178 21784 36184
rect 21916 36236 21968 36242
rect 21916 36178 21968 36184
rect 21744 36106 21772 36178
rect 21732 36100 21784 36106
rect 21732 36042 21784 36048
rect 21744 35698 21772 36042
rect 21928 35766 21956 36178
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21364 34672 21416 34678
rect 21364 34614 21416 34620
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21928 33454 21956 33798
rect 21916 33448 21968 33454
rect 21916 33390 21968 33396
rect 22020 33386 22048 37062
rect 22664 36718 22692 39782
rect 22756 39642 22784 40462
rect 22848 40186 22876 41210
rect 23020 41132 23072 41138
rect 23020 41074 23072 41080
rect 22836 40180 22888 40186
rect 22836 40122 22888 40128
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 23032 38962 23060 41074
rect 23400 40934 23428 41550
rect 23388 40928 23440 40934
rect 23388 40870 23440 40876
rect 23112 40112 23164 40118
rect 23112 40054 23164 40060
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 23032 38486 23060 38898
rect 23020 38480 23072 38486
rect 23020 38422 23072 38428
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 22756 37874 22784 38150
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 23032 37670 23060 38422
rect 23020 37664 23072 37670
rect 23020 37606 23072 37612
rect 22744 37324 22796 37330
rect 23124 37312 23152 40054
rect 23296 39500 23348 39506
rect 23296 39442 23348 39448
rect 23308 39030 23336 39442
rect 23400 39098 23428 40870
rect 23756 39976 23808 39982
rect 23756 39918 23808 39924
rect 23388 39092 23440 39098
rect 23388 39034 23440 39040
rect 23296 39024 23348 39030
rect 23296 38966 23348 38972
rect 23664 37800 23716 37806
rect 23664 37742 23716 37748
rect 23676 37466 23704 37742
rect 23664 37460 23716 37466
rect 23664 37402 23716 37408
rect 23204 37324 23256 37330
rect 23124 37284 23204 37312
rect 22744 37266 22796 37272
rect 23204 37266 23256 37272
rect 22756 36922 22784 37266
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 23216 36854 23244 37266
rect 23204 36848 23256 36854
rect 23204 36790 23256 36796
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22664 36582 22692 36654
rect 22652 36576 22704 36582
rect 22652 36518 22704 36524
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22204 35154 22232 36110
rect 22664 35329 22692 36518
rect 23112 36304 23164 36310
rect 23112 36246 23164 36252
rect 23124 35834 23152 36246
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23492 35834 23520 36110
rect 23112 35828 23164 35834
rect 23112 35770 23164 35776
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 22836 35488 22888 35494
rect 22836 35430 22888 35436
rect 22650 35320 22706 35329
rect 22560 35284 22612 35290
rect 22650 35255 22706 35264
rect 22560 35226 22612 35232
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 22204 34746 22232 35090
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22572 34678 22600 35226
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 21364 33380 21416 33386
rect 21364 33322 21416 33328
rect 22008 33380 22060 33386
rect 22008 33322 22060 33328
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 21008 33106 21128 33134
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20536 32496 20588 32502
rect 20536 32438 20588 32444
rect 20352 32360 20404 32366
rect 20352 32302 20404 32308
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20456 31414 20484 32166
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20260 31204 20312 31210
rect 20088 31164 20208 31192
rect 19984 31136 20036 31142
rect 20036 31096 20116 31124
rect 19984 31078 20036 31084
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19904 29034 19932 29650
rect 19996 29646 20024 29990
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19996 29306 20024 29582
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 20088 29050 20116 31096
rect 20180 30938 20208 31164
rect 20260 31146 20312 31152
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20180 30394 20208 30874
rect 20272 30598 20300 31146
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 20180 30190 20208 30330
rect 20272 30326 20300 30534
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 20364 29850 20392 30670
rect 20456 30054 20484 30738
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 29170 20208 29446
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 19892 29028 19944 29034
rect 20088 29022 20208 29050
rect 19892 28970 19944 28976
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19904 28393 19932 28970
rect 19890 28384 19946 28393
rect 19890 28319 19946 28328
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19892 27328 19944 27334
rect 19892 27270 19944 27276
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19904 26042 19932 27270
rect 19996 26994 20024 27814
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26586 20024 26930
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 20076 26240 20128 26246
rect 20076 26182 20128 26188
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19904 24954 19932 25978
rect 20088 25906 20116 26182
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25498 20116 25842
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19076 24313 19104 24346
rect 19062 24304 19118 24313
rect 19062 24239 19118 24248
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19076 21622 19104 23666
rect 19168 23202 19196 24754
rect 19996 24682 20024 25094
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20088 24682 20116 24890
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 19984 24676 20036 24682
rect 19984 24618 20036 24624
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19352 24342 19380 24618
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 20088 24342 20116 24618
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19260 23322 19288 24142
rect 19352 23866 19380 24278
rect 20180 24206 20208 29022
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 20272 25770 20300 26726
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20364 25770 20392 25842
rect 20260 25764 20312 25770
rect 20260 25706 20312 25712
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19720 23730 19748 24006
rect 19996 23798 20024 24142
rect 20272 23866 20300 25706
rect 20364 25294 20392 25706
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19444 23526 19472 23591
rect 19708 23588 19760 23594
rect 19812 23576 19840 23666
rect 19760 23548 19840 23576
rect 19708 23530 19760 23536
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19444 23202 19472 23462
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19168 23174 19472 23202
rect 19616 23180 19668 23186
rect 19168 22642 19196 23174
rect 19616 23122 19668 23128
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19628 22506 19656 23122
rect 19616 22500 19668 22506
rect 19616 22442 19668 22448
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19996 22166 20024 23734
rect 20168 23588 20220 23594
rect 20272 23576 20300 23802
rect 20456 23769 20484 29990
rect 20442 23760 20498 23769
rect 20442 23695 20498 23704
rect 20220 23548 20300 23576
rect 20168 23530 20220 23536
rect 20180 22982 20208 23530
rect 20548 23474 20576 32302
rect 20640 29753 20668 32710
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20732 30802 20760 32438
rect 20720 30796 20772 30802
rect 20720 30738 20772 30744
rect 20720 30116 20772 30122
rect 20720 30058 20772 30064
rect 20626 29744 20682 29753
rect 20626 29679 20682 29688
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20272 23446 20576 23474
rect 20168 22976 20220 22982
rect 20168 22918 20220 22924
rect 20180 22506 20208 22918
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19246 21720 19302 21729
rect 19352 21690 19380 21966
rect 19246 21655 19302 21664
rect 19340 21684 19392 21690
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 19260 21146 19288 21655
rect 19340 21626 19392 21632
rect 19444 21554 19472 22102
rect 20088 21962 20116 22442
rect 20180 22234 20208 22442
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 20272 21690 20300 23446
rect 20640 23254 20668 24618
rect 20732 23474 20760 30058
rect 20824 29714 20852 33050
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20902 28792 20958 28801
rect 20902 28727 20958 28736
rect 20916 28626 20944 28727
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20916 28218 20944 28562
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 21008 23474 21036 33106
rect 21088 33040 21140 33046
rect 21376 33017 21404 33322
rect 21732 33312 21784 33318
rect 21732 33254 21784 33260
rect 21088 32982 21140 32988
rect 21362 33008 21418 33017
rect 21100 32230 21128 32982
rect 21362 32943 21418 32952
rect 21640 32836 21692 32842
rect 21640 32778 21692 32784
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 21100 30122 21128 32166
rect 21652 31958 21680 32778
rect 21744 32366 21772 33254
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21928 32026 21956 32302
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21640 31952 21692 31958
rect 21640 31894 21692 31900
rect 21652 31346 21680 31894
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21744 31482 21772 31758
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 22284 31272 22336 31278
rect 22284 31214 22336 31220
rect 21272 31204 21324 31210
rect 21272 31146 21324 31152
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 21192 30870 21220 31078
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 21192 30394 21220 30806
rect 21180 30388 21232 30394
rect 21180 30330 21232 30336
rect 21284 30326 21312 31146
rect 22296 30938 22324 31214
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 21088 30116 21140 30122
rect 21088 30058 21140 30064
rect 21100 29782 21128 30058
rect 21088 29776 21140 29782
rect 21088 29718 21140 29724
rect 21100 29306 21128 29718
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 21100 29034 21128 29242
rect 21376 29238 21404 30602
rect 22388 30394 22416 33390
rect 22376 30388 22428 30394
rect 22376 30330 22428 30336
rect 21364 29232 21416 29238
rect 21364 29174 21416 29180
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 21284 28762 21312 29106
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21100 28014 21128 28358
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21468 27946 21496 28358
rect 21836 28014 21864 28970
rect 21824 28008 21876 28014
rect 21824 27950 21876 27956
rect 21456 27940 21508 27946
rect 21456 27882 21508 27888
rect 21468 27538 21496 27882
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 21456 27532 21508 27538
rect 21456 27474 21508 27480
rect 21100 27130 21128 27474
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21100 26450 21128 26862
rect 21468 26586 21496 27474
rect 21732 27464 21784 27470
rect 21732 27406 21784 27412
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21744 26450 21772 27406
rect 21928 26994 21956 27814
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21928 26586 21956 26930
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 22020 26518 22048 26794
rect 22008 26512 22060 26518
rect 22008 26454 22060 26460
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21100 25702 21128 26386
rect 21732 26036 21784 26042
rect 21732 25978 21784 25984
rect 21744 25770 21772 25978
rect 22020 25906 22048 26454
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22204 25974 22232 26182
rect 22192 25968 22244 25974
rect 22192 25910 22244 25916
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22020 25777 22048 25842
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 22468 25764 22520 25770
rect 22468 25706 22520 25712
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21100 25430 21128 25638
rect 21088 25424 21140 25430
rect 21088 25366 21140 25372
rect 21916 25424 21968 25430
rect 21916 25366 21968 25372
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21456 24676 21508 24682
rect 21456 24618 21508 24624
rect 21468 23866 21496 24618
rect 21560 24614 21588 25298
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21364 23656 21416 23662
rect 21284 23633 21364 23644
rect 21270 23624 21364 23633
rect 21326 23616 21364 23624
rect 21364 23598 21416 23604
rect 21270 23559 21326 23568
rect 20732 23446 20852 23474
rect 21008 23446 21128 23474
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20640 22710 20668 23190
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 22098 20392 22374
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 20536 21480 20588 21486
rect 20824 21457 20852 23446
rect 20536 21422 20588 21428
rect 20810 21448 20866 21457
rect 20548 21350 20576 21422
rect 20810 21383 20866 21392
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 17788 20330 17816 20538
rect 18708 20534 18736 20878
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17776 20324 17828 20330
rect 17776 20266 17828 20272
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16500 18970 16528 19246
rect 16868 18970 16896 19858
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 17144 18834 17172 19178
rect 17512 19174 17540 19858
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17144 18426 17172 18770
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16868 17338 16896 17682
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16960 15910 16988 16594
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16316 13786 16436 13814
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 12986 16160 13262
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 10810 16160 12922
rect 16224 12646 16252 13738
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16132 10130 16160 10746
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16132 9722 16160 10066
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16224 9518 16252 12582
rect 16316 10538 16344 13786
rect 16960 13326 16988 15846
rect 17420 14618 17448 18906
rect 17512 16658 17540 19110
rect 17788 18970 17816 20266
rect 18064 20058 18092 20334
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18248 19922 18276 20198
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17788 18426 17816 18906
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17788 17814 17816 18362
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17788 17270 17816 17750
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17512 16250 17540 16594
rect 18064 16538 18092 19382
rect 18524 19310 18552 19858
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 17746 18184 19110
rect 18524 18970 18552 19246
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18154 18368 18566
rect 18708 18358 18736 20470
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18524 17542 18552 18226
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16794 18184 17138
rect 18248 17066 18276 17478
rect 18524 17338 18552 17478
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18236 16584 18288 16590
rect 18142 16552 18198 16561
rect 18064 16510 18142 16538
rect 18236 16526 18288 16532
rect 18142 16487 18198 16496
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 18156 15570 18184 16487
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18156 15162 18184 15506
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17604 14414 17632 14758
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 14074 17632 14350
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17958 13832 18014 13841
rect 17040 13728 17092 13734
rect 17092 13688 17172 13716
rect 17040 13670 17092 13676
rect 17144 13462 17172 13688
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16960 12646 16988 13262
rect 17144 13190 17172 13398
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12714 17172 13126
rect 17880 12986 17908 13806
rect 17958 13767 17960 13776
rect 18012 13767 18014 13776
rect 17960 13738 18012 13744
rect 17972 13394 18000 13738
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 18248 12986 18276 16526
rect 18432 13530 18460 16934
rect 18616 16726 18644 17274
rect 18708 17270 18736 18294
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18800 17082 18828 20742
rect 18984 20602 19012 21014
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19514 19380 19858
rect 20088 19718 20116 20334
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17202 18920 17478
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18800 17054 18920 17082
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18524 16046 18552 16594
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 15570 18552 15982
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18524 15162 18552 15506
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 17144 9382 17172 12650
rect 17880 12442 17908 12922
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 17868 12436 17920 12442
rect 17788 12396 17868 12424
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17420 11558 17448 12242
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 13818 8936 13874 8945
rect 13818 8871 13874 8880
rect 17144 2009 17172 9318
rect 17130 2000 17186 2009
rect 17130 1935 17186 1944
rect 10598 54 11008 82
rect 17420 82 17448 11494
rect 17788 10742 17816 12396
rect 17868 12378 17920 12384
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17880 10470 17908 11154
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17512 10266 17540 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17880 10062 17908 10406
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17880 9722 17908 9998
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17880 9178 17908 9658
rect 17972 9178 18000 12582
rect 18524 11898 18552 12582
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 11762 18644 16050
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18708 13814 18736 14486
rect 18708 13802 18828 13814
rect 18708 13796 18840 13802
rect 18708 13786 18788 13796
rect 18788 13738 18840 13744
rect 18800 13190 18828 13738
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 11354 18644 11698
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18144 9444 18196 9450
rect 18248 9432 18276 10134
rect 18196 9404 18276 9432
rect 18144 9386 18196 9392
rect 18800 9382 18828 10406
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18616 9110 18644 9318
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18800 9042 18828 9318
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18708 8498 18736 8978
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18892 7954 18920 17054
rect 19260 16658 19288 19246
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 18086 19472 18770
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19996 18086 20024 18158
rect 20088 18154 20116 19654
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20272 19242 20300 19314
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16250 19288 16594
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 12306 19012 15438
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 13938 19104 14894
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19076 13705 19104 13874
rect 19062 13696 19118 13705
rect 19062 13631 19118 13640
rect 19076 13530 19104 13631
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19168 12696 19196 15030
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19260 13852 19288 14418
rect 19444 14346 19472 18022
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19536 17066 19564 17682
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19720 16250 19748 16594
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19904 15026 19932 17614
rect 19996 17048 20024 18022
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20364 17338 20392 17614
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20076 17060 20128 17066
rect 19996 17020 20076 17048
rect 20076 17002 20128 17008
rect 19984 16584 20036 16590
rect 20088 16561 20116 17002
rect 19984 16526 20036 16532
rect 20074 16552 20130 16561
rect 19996 16114 20024 16526
rect 20364 16522 20392 17070
rect 20074 16487 20130 16496
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 15706 20484 16050
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19904 14550 19932 14962
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19340 13864 19392 13870
rect 19260 13841 19340 13852
rect 19246 13832 19340 13841
rect 19302 13824 19340 13832
rect 19340 13806 19392 13812
rect 19246 13767 19302 13776
rect 19292 13696 19348 13705
rect 19348 13654 19472 13682
rect 19292 13631 19348 13640
rect 19444 13433 19472 13654
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19430 13424 19486 13433
rect 19430 13359 19486 13368
rect 19248 12708 19300 12714
rect 19168 12668 19248 12696
rect 19248 12650 19300 12656
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 12442 19380 12650
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11898 19012 12242
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18984 10810 19012 11086
rect 19168 10810 19196 11222
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19444 10470 19472 11494
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19904 11286 19932 12038
rect 20548 11898 20576 21286
rect 20904 20324 20956 20330
rect 20904 20266 20956 20272
rect 20916 19854 20944 20266
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19514 20944 19790
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20640 17338 20668 19178
rect 20732 18630 20760 19314
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18290 20760 18566
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20640 17066 20668 17274
rect 21008 17202 21036 17818
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20640 16250 20668 17002
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 15978 20668 16186
rect 21100 16182 21128 23446
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21376 22710 21404 23122
rect 21560 22817 21588 24550
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21836 23322 21864 24278
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 21928 23050 21956 25366
rect 22204 24682 22232 25366
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22204 24342 22232 24618
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 22204 23866 22232 24278
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21546 22808 21602 22817
rect 21546 22743 21602 22752
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21560 21486 21588 22743
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21652 21350 21680 21830
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21284 20602 21312 20878
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21284 19242 21312 19994
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18902 21404 19110
rect 21560 18902 21588 20198
rect 21836 20058 21864 20266
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 21928 19938 21956 22986
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22204 22506 22232 22714
rect 22388 22642 22416 24754
rect 22480 24410 22508 25706
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22112 22234 22140 22442
rect 22480 22234 22508 23054
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 21350 22048 22034
rect 22480 21690 22508 22170
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 21836 19910 21956 19938
rect 22388 19922 22416 20198
rect 22376 19916 22428 19922
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21376 18426 21404 18838
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21560 18426 21588 18702
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21192 16794 21220 17682
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21560 16726 21588 16934
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21468 16114 21496 16526
rect 21560 16250 21588 16662
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20640 14890 20668 15914
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21376 15638 21404 15846
rect 21744 15638 21772 16526
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20640 14006 20668 14826
rect 20732 14618 20760 15574
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 15162 21128 15438
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20824 14550 20852 14758
rect 21100 14600 21128 15098
rect 21180 14612 21232 14618
rect 21100 14572 21180 14600
rect 21180 14554 21232 14560
rect 21744 14550 21772 15574
rect 21836 15434 21864 19910
rect 22376 19858 22428 19864
rect 22572 18222 22600 34342
rect 22664 33114 22692 35255
rect 22848 34746 22876 35430
rect 23570 34776 23626 34785
rect 22836 34740 22888 34746
rect 23570 34711 23626 34720
rect 22836 34682 22888 34688
rect 22848 34542 22876 34682
rect 23112 34672 23164 34678
rect 23112 34614 23164 34620
rect 22836 34536 22888 34542
rect 22834 34504 22836 34513
rect 22888 34504 22890 34513
rect 22834 34439 22890 34448
rect 22928 34400 22980 34406
rect 22928 34342 22980 34348
rect 22940 34202 22968 34342
rect 22928 34196 22980 34202
rect 22928 34138 22980 34144
rect 22744 34060 22796 34066
rect 22744 34002 22796 34008
rect 22756 33658 22784 34002
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22652 33108 22704 33114
rect 22652 33050 22704 33056
rect 22652 32904 22704 32910
rect 22756 32881 22784 33594
rect 22836 33380 22888 33386
rect 22836 33322 22888 33328
rect 22652 32846 22704 32852
rect 22742 32872 22798 32881
rect 22664 32570 22692 32846
rect 22742 32807 22798 32816
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22848 30326 22876 33322
rect 23124 33046 23152 34614
rect 23584 34542 23612 34711
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23204 34060 23256 34066
rect 23204 34002 23256 34008
rect 23216 33658 23244 34002
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23112 33040 23164 33046
rect 23112 32982 23164 32988
rect 23124 32298 23152 32982
rect 23112 32292 23164 32298
rect 23112 32234 23164 32240
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 23032 31278 23060 31826
rect 23020 31272 23072 31278
rect 23020 31214 23072 31220
rect 23124 30734 23152 32234
rect 23216 31890 23244 33594
rect 23308 32978 23336 33934
rect 23768 33017 23796 39918
rect 23860 39846 23888 41958
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 24412 40730 24440 41550
rect 24504 40769 24532 43046
rect 24780 42906 24808 43114
rect 24768 42900 24820 42906
rect 24768 42842 24820 42848
rect 24952 42832 25004 42838
rect 24952 42774 25004 42780
rect 24676 42696 24728 42702
rect 24676 42638 24728 42644
rect 24584 42016 24636 42022
rect 24584 41958 24636 41964
rect 24490 40760 24546 40769
rect 24400 40724 24452 40730
rect 24490 40695 24546 40704
rect 24400 40666 24452 40672
rect 24490 40624 24546 40633
rect 24308 40588 24360 40594
rect 24490 40559 24546 40568
rect 24308 40530 24360 40536
rect 24320 39846 24348 40530
rect 23848 39840 23900 39846
rect 23848 39782 23900 39788
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24124 39500 24176 39506
rect 24124 39442 24176 39448
rect 24136 38826 24164 39442
rect 24124 38820 24176 38826
rect 24124 38762 24176 38768
rect 23940 38208 23992 38214
rect 23940 38150 23992 38156
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 23860 36310 23888 37606
rect 23952 36650 23980 38150
rect 24124 37120 24176 37126
rect 24124 37062 24176 37068
rect 24136 36786 24164 37062
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24216 36780 24268 36786
rect 24216 36722 24268 36728
rect 23940 36644 23992 36650
rect 23940 36586 23992 36592
rect 23952 36378 23980 36586
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 23848 36304 23900 36310
rect 23848 36246 23900 36252
rect 24136 35834 24164 36722
rect 24228 36242 24256 36722
rect 24216 36236 24268 36242
rect 24216 36178 24268 36184
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 24228 35562 24256 36178
rect 24320 35766 24348 39782
rect 24504 38894 24532 40559
rect 24596 39506 24624 41958
rect 24688 41818 24716 42638
rect 24964 42294 24992 42774
rect 24952 42288 25004 42294
rect 24952 42230 25004 42236
rect 24676 41812 24728 41818
rect 24676 41754 24728 41760
rect 24964 41750 24992 42230
rect 25136 42084 25188 42090
rect 25136 42026 25188 42032
rect 25044 42016 25096 42022
rect 25044 41958 25096 41964
rect 24952 41744 25004 41750
rect 24952 41686 25004 41692
rect 24964 41206 24992 41686
rect 24952 41200 25004 41206
rect 24952 41142 25004 41148
rect 24768 41132 24820 41138
rect 24768 41074 24820 41080
rect 24674 40760 24730 40769
rect 24780 40730 24808 41074
rect 24674 40695 24730 40704
rect 24768 40724 24820 40730
rect 24584 39500 24636 39506
rect 24584 39442 24636 39448
rect 24492 38888 24544 38894
rect 24492 38830 24544 38836
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24492 38548 24544 38554
rect 24492 38490 24544 38496
rect 24504 36854 24532 38490
rect 24596 38350 24624 38694
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 24688 37330 24716 40695
rect 24768 40666 24820 40672
rect 25056 40662 25084 41958
rect 25148 41478 25176 42026
rect 25136 41472 25188 41478
rect 25136 41414 25188 41420
rect 25148 41274 25176 41414
rect 25136 41268 25188 41274
rect 25136 41210 25188 41216
rect 25136 40996 25188 41002
rect 25136 40938 25188 40944
rect 25044 40656 25096 40662
rect 25044 40598 25096 40604
rect 24952 40520 25004 40526
rect 24952 40462 25004 40468
rect 24964 39914 24992 40462
rect 25056 40186 25084 40598
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 24952 39908 25004 39914
rect 24952 39850 25004 39856
rect 24964 39642 24992 39850
rect 24952 39636 25004 39642
rect 24952 39578 25004 39584
rect 24952 39296 25004 39302
rect 24952 39238 25004 39244
rect 24860 38820 24912 38826
rect 24860 38762 24912 38768
rect 24676 37324 24728 37330
rect 24676 37266 24728 37272
rect 24688 36922 24716 37266
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24492 36848 24544 36854
rect 24492 36790 24544 36796
rect 24504 36242 24532 36790
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 24504 35834 24532 36178
rect 24492 35828 24544 35834
rect 24492 35770 24544 35776
rect 24308 35760 24360 35766
rect 24308 35702 24360 35708
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24032 35556 24084 35562
rect 24032 35498 24084 35504
rect 24216 35556 24268 35562
rect 24216 35498 24268 35504
rect 24044 35086 24072 35498
rect 24124 35216 24176 35222
rect 24124 35158 24176 35164
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24044 34678 24072 35022
rect 24136 34746 24164 35158
rect 24308 35080 24360 35086
rect 24308 35022 24360 35028
rect 24124 34740 24176 34746
rect 24124 34682 24176 34688
rect 24032 34672 24084 34678
rect 24032 34614 24084 34620
rect 24320 34542 24348 35022
rect 24308 34536 24360 34542
rect 24308 34478 24360 34484
rect 24124 34196 24176 34202
rect 24124 34138 24176 34144
rect 24136 33522 24164 34138
rect 24596 33590 24624 35566
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24688 33658 24716 33934
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 24780 33522 24808 33934
rect 24872 33590 24900 38762
rect 24964 38486 24992 39238
rect 25148 39030 25176 40938
rect 25136 39024 25188 39030
rect 25136 38966 25188 38972
rect 25148 38826 25176 38966
rect 25136 38820 25188 38826
rect 25136 38762 25188 38768
rect 24952 38480 25004 38486
rect 24952 38422 25004 38428
rect 24964 37466 24992 38422
rect 24952 37460 25004 37466
rect 24952 37402 25004 37408
rect 25332 37330 25360 43794
rect 25596 43172 25648 43178
rect 25596 43114 25648 43120
rect 25608 42770 25636 43114
rect 25596 42764 25648 42770
rect 25596 42706 25648 42712
rect 25700 42140 25728 44338
rect 25780 42152 25832 42158
rect 25700 42112 25780 42140
rect 25780 42094 25832 42100
rect 25884 41750 25912 44814
rect 27080 44198 27108 44882
rect 27436 44736 27488 44742
rect 27436 44678 27488 44684
rect 27448 44402 27476 44678
rect 27436 44396 27488 44402
rect 27436 44338 27488 44344
rect 27068 44192 27120 44198
rect 27068 44134 27120 44140
rect 27160 44192 27212 44198
rect 27160 44134 27212 44140
rect 26792 43852 26844 43858
rect 26792 43794 26844 43800
rect 26608 43648 26660 43654
rect 26608 43590 26660 43596
rect 26620 43450 26648 43590
rect 26608 43444 26660 43450
rect 26608 43386 26660 43392
rect 26804 43110 26832 43794
rect 27080 43761 27108 44134
rect 27172 43994 27200 44134
rect 27448 43994 27476 44338
rect 27632 44266 27660 45018
rect 27724 44470 27752 45290
rect 28184 45014 28212 46310
rect 28460 45393 28488 46310
rect 30196 46164 30248 46170
rect 30196 46106 30248 46112
rect 28724 46096 28776 46102
rect 28724 46038 28776 46044
rect 28632 45960 28684 45966
rect 28632 45902 28684 45908
rect 28644 45626 28672 45902
rect 28736 45626 28764 46038
rect 29000 45960 29052 45966
rect 29000 45902 29052 45908
rect 28632 45620 28684 45626
rect 28632 45562 28684 45568
rect 28724 45620 28776 45626
rect 28724 45562 28776 45568
rect 28724 45484 28776 45490
rect 28724 45426 28776 45432
rect 28446 45384 28502 45393
rect 28446 45319 28502 45328
rect 28172 45008 28224 45014
rect 28172 44950 28224 44956
rect 28448 45008 28500 45014
rect 28448 44950 28500 44956
rect 27804 44872 27856 44878
rect 27804 44814 27856 44820
rect 27712 44464 27764 44470
rect 27712 44406 27764 44412
rect 27816 44402 27844 44814
rect 28184 44538 28212 44950
rect 28172 44532 28224 44538
rect 28172 44474 28224 44480
rect 27804 44396 27856 44402
rect 27804 44338 27856 44344
rect 27620 44260 27672 44266
rect 27620 44202 27672 44208
rect 27160 43988 27212 43994
rect 27160 43930 27212 43936
rect 27436 43988 27488 43994
rect 27436 43930 27488 43936
rect 27632 43858 27660 44202
rect 28460 44198 28488 44950
rect 28448 44192 28500 44198
rect 28448 44134 28500 44140
rect 28448 43920 28500 43926
rect 28448 43862 28500 43868
rect 27436 43852 27488 43858
rect 27436 43794 27488 43800
rect 27620 43852 27672 43858
rect 27620 43794 27672 43800
rect 27066 43752 27122 43761
rect 27066 43687 27122 43696
rect 25964 43104 26016 43110
rect 25964 43046 26016 43052
rect 26792 43104 26844 43110
rect 26792 43046 26844 43052
rect 25976 42838 26004 43046
rect 25964 42832 26016 42838
rect 25964 42774 26016 42780
rect 25976 42022 26004 42774
rect 26804 42673 26832 43046
rect 26884 42900 26936 42906
rect 26884 42842 26936 42848
rect 26790 42664 26846 42673
rect 26790 42599 26846 42608
rect 26516 42152 26568 42158
rect 26804 42129 26832 42599
rect 26516 42094 26568 42100
rect 26790 42120 26846 42129
rect 26528 42022 26556 42094
rect 26790 42055 26846 42064
rect 25964 42016 26016 42022
rect 25964 41958 26016 41964
rect 26516 42016 26568 42022
rect 26516 41958 26568 41964
rect 25872 41744 25924 41750
rect 25872 41686 25924 41692
rect 25884 41274 25912 41686
rect 26516 41676 26568 41682
rect 26516 41618 26568 41624
rect 25872 41268 25924 41274
rect 25872 41210 25924 41216
rect 25884 40662 25912 41210
rect 26528 40934 26556 41618
rect 26792 41540 26844 41546
rect 26792 41482 26844 41488
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 25872 40656 25924 40662
rect 26528 40633 26556 40870
rect 25872 40598 25924 40604
rect 26514 40624 26570 40633
rect 26514 40559 26570 40568
rect 26528 40361 26556 40559
rect 26514 40352 26570 40361
rect 26514 40287 26570 40296
rect 26804 39982 26832 41482
rect 26896 41138 26924 42842
rect 27080 42634 27108 43687
rect 27448 43178 27476 43794
rect 28356 43784 28408 43790
rect 28356 43726 28408 43732
rect 28368 43450 28396 43726
rect 28356 43444 28408 43450
rect 28356 43386 28408 43392
rect 28460 43314 28488 43862
rect 28632 43444 28684 43450
rect 28632 43386 28684 43392
rect 27620 43308 27672 43314
rect 27620 43250 27672 43256
rect 28448 43308 28500 43314
rect 28448 43250 28500 43256
rect 27436 43172 27488 43178
rect 27436 43114 27488 43120
rect 27160 42764 27212 42770
rect 27160 42706 27212 42712
rect 27344 42764 27396 42770
rect 27344 42706 27396 42712
rect 27068 42628 27120 42634
rect 27068 42570 27120 42576
rect 27172 42294 27200 42706
rect 27356 42362 27384 42706
rect 27344 42356 27396 42362
rect 27344 42298 27396 42304
rect 27160 42288 27212 42294
rect 27160 42230 27212 42236
rect 26976 42084 27028 42090
rect 26976 42026 27028 42032
rect 26988 41818 27016 42026
rect 26976 41812 27028 41818
rect 26976 41754 27028 41760
rect 26884 41132 26936 41138
rect 26884 41074 26936 41080
rect 26976 40588 27028 40594
rect 26976 40530 27028 40536
rect 26988 40118 27016 40530
rect 27172 40458 27200 42230
rect 27356 40594 27384 42298
rect 27632 42158 27660 43250
rect 28460 42838 28488 43250
rect 28448 42832 28500 42838
rect 28448 42774 28500 42780
rect 28356 42764 28408 42770
rect 28356 42706 28408 42712
rect 28080 42628 28132 42634
rect 28080 42570 28132 42576
rect 27620 42152 27672 42158
rect 27620 42094 27672 42100
rect 27896 42084 27948 42090
rect 27896 42026 27948 42032
rect 27908 41614 27936 42026
rect 27988 41744 28040 41750
rect 27988 41686 28040 41692
rect 27896 41608 27948 41614
rect 27896 41550 27948 41556
rect 27620 41472 27672 41478
rect 27620 41414 27672 41420
rect 27632 41070 27660 41414
rect 27620 41064 27672 41070
rect 27620 41006 27672 41012
rect 27344 40588 27396 40594
rect 27344 40530 27396 40536
rect 27160 40452 27212 40458
rect 27160 40394 27212 40400
rect 26976 40112 27028 40118
rect 27028 40072 27108 40100
rect 26976 40054 27028 40060
rect 26792 39976 26844 39982
rect 26792 39918 26844 39924
rect 26056 39908 26108 39914
rect 26056 39850 26108 39856
rect 25504 39840 25556 39846
rect 25504 39782 25556 39788
rect 25516 39302 25544 39782
rect 25964 39636 26016 39642
rect 25964 39578 26016 39584
rect 25504 39296 25556 39302
rect 25504 39238 25556 39244
rect 25516 38962 25544 39238
rect 25504 38956 25556 38962
rect 25504 38898 25556 38904
rect 25976 38894 26004 39578
rect 25964 38888 26016 38894
rect 25964 38830 26016 38836
rect 25976 38554 26004 38830
rect 25964 38548 26016 38554
rect 25964 38490 26016 38496
rect 25688 37732 25740 37738
rect 25688 37674 25740 37680
rect 25320 37324 25372 37330
rect 25320 37266 25372 37272
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 24952 35488 25004 35494
rect 24952 35430 25004 35436
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24124 33380 24176 33386
rect 24124 33322 24176 33328
rect 24136 33114 24164 33322
rect 24124 33108 24176 33114
rect 24124 33050 24176 33056
rect 23754 33008 23810 33017
rect 23296 32972 23348 32978
rect 23754 32943 23810 32952
rect 23296 32914 23348 32920
rect 23308 32570 23336 32914
rect 23296 32564 23348 32570
rect 23296 32506 23348 32512
rect 24584 32564 24636 32570
rect 24584 32506 24636 32512
rect 24492 32428 24544 32434
rect 24412 32388 24492 32416
rect 23204 31884 23256 31890
rect 23204 31826 23256 31832
rect 23216 31346 23244 31826
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 24032 31816 24084 31822
rect 24032 31758 24084 31764
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23124 30394 23152 30670
rect 23112 30388 23164 30394
rect 23112 30330 23164 30336
rect 22836 30320 22888 30326
rect 22742 30288 22798 30297
rect 22836 30262 22888 30268
rect 22742 30223 22798 30232
rect 22756 30190 22784 30223
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22652 28960 22704 28966
rect 22652 28902 22704 28908
rect 22664 28014 22692 28902
rect 22848 28762 22876 30262
rect 23216 29714 23244 31282
rect 23308 30938 23336 31758
rect 24044 31414 24072 31758
rect 24412 31686 24440 32388
rect 24492 32370 24544 32376
rect 24596 32298 24624 32506
rect 24780 32434 24808 33458
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 24584 32292 24636 32298
rect 24584 32234 24636 32240
rect 24596 31958 24624 32234
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24412 31482 24440 31622
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24032 31408 24084 31414
rect 24032 31350 24084 31356
rect 24780 31346 24808 32370
rect 24964 31346 24992 35430
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25148 34134 25176 34342
rect 25136 34128 25188 34134
rect 25136 34070 25188 34076
rect 25148 33318 25176 34070
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 25148 33046 25176 33254
rect 25136 33040 25188 33046
rect 25136 32982 25188 32988
rect 24768 31340 24820 31346
rect 24952 31340 25004 31346
rect 24768 31282 24820 31288
rect 24872 31300 24952 31328
rect 23940 31272 23992 31278
rect 23940 31214 23992 31220
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23676 29782 23704 30126
rect 23768 30122 23796 30330
rect 23756 30116 23808 30122
rect 23756 30058 23808 30064
rect 23768 29850 23796 30058
rect 23756 29844 23808 29850
rect 23756 29786 23808 29792
rect 23664 29776 23716 29782
rect 23664 29718 23716 29724
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 23204 29708 23256 29714
rect 23204 29650 23256 29656
rect 22940 29034 22968 29650
rect 23216 29306 23244 29650
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 22928 29028 22980 29034
rect 22928 28970 22980 28976
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22664 27470 22692 27950
rect 22756 27538 22784 28494
rect 22848 28218 22876 28698
rect 22836 28212 22888 28218
rect 22836 28154 22888 28160
rect 22744 27532 22796 27538
rect 22744 27474 22796 27480
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22756 27130 22784 27474
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22940 27062 22968 28970
rect 23216 28490 23244 29242
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23492 28626 23520 28902
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23478 28520 23534 28529
rect 23204 28484 23256 28490
rect 23478 28455 23534 28464
rect 23204 28426 23256 28432
rect 23492 28014 23520 28455
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 23032 26858 23060 27542
rect 23848 27396 23900 27402
rect 23848 27338 23900 27344
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22756 25430 22784 26726
rect 22928 26444 22980 26450
rect 22928 26386 22980 26392
rect 22940 26042 22968 26386
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 22834 25800 22890 25809
rect 22834 25735 22890 25744
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22664 24410 22692 25230
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22664 23866 22692 24346
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22756 23118 22784 24142
rect 22848 23866 22876 25735
rect 23308 24954 23336 26182
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23308 24682 23336 24890
rect 23296 24676 23348 24682
rect 23296 24618 23348 24624
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22940 23798 22968 24074
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 23308 23254 23336 24618
rect 23492 24342 23520 27270
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 23866 23428 24142
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23400 23322 23428 23802
rect 23492 23730 23520 24278
rect 23676 24041 23704 25774
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23768 24818 23796 25434
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23662 24032 23718 24041
rect 23662 23967 23718 23976
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 23308 22778 23336 23190
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22940 22030 22968 22578
rect 23308 22234 23336 22714
rect 23492 22506 23520 23666
rect 23860 23594 23888 27338
rect 23952 26450 23980 31214
rect 24584 31204 24636 31210
rect 24584 31146 24636 31152
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24124 30592 24176 30598
rect 24124 30534 24176 30540
rect 24136 29782 24164 30534
rect 24412 30394 24440 31078
rect 24596 30938 24624 31146
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24400 30388 24452 30394
rect 24400 30330 24452 30336
rect 24124 29776 24176 29782
rect 24124 29718 24176 29724
rect 24136 29306 24164 29718
rect 24780 29646 24808 31282
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24688 29306 24716 29514
rect 24780 29306 24808 29582
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24688 29102 24716 29242
rect 24676 29096 24728 29102
rect 24676 29038 24728 29044
rect 24124 28960 24176 28966
rect 24044 28920 24124 28948
rect 23940 26444 23992 26450
rect 23940 26386 23992 26392
rect 23952 25945 23980 26386
rect 23938 25936 23994 25945
rect 23938 25871 23994 25880
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 23952 24818 23980 25230
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23952 24138 23980 24754
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23848 23588 23900 23594
rect 23848 23530 23900 23536
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22756 21418 22784 21966
rect 23032 21690 23060 22102
rect 23662 21856 23718 21865
rect 23662 21791 23718 21800
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 23572 21412 23624 21418
rect 23572 21354 23624 21360
rect 22756 21146 22784 21354
rect 23584 21146 23612 21354
rect 23676 21350 23704 21791
rect 23768 21350 23796 22646
rect 23860 22642 23888 22918
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23952 21418 23980 22170
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22664 20602 22692 20946
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 23676 20516 23704 21286
rect 23584 20488 23704 20516
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22664 18714 22692 19314
rect 23112 19304 23164 19310
rect 23110 19272 23112 19281
rect 23164 19272 23166 19281
rect 23308 19242 23336 19926
rect 23492 19854 23520 20266
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23110 19207 23166 19216
rect 23296 19236 23348 19242
rect 23124 19174 23152 19207
rect 23296 19178 23348 19184
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 23112 19168 23164 19174
rect 23400 19145 23428 19450
rect 23112 19110 23164 19116
rect 23386 19136 23442 19145
rect 22756 18834 22784 19110
rect 23386 19071 23442 19080
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 22664 18698 22784 18714
rect 22664 18692 22796 18698
rect 22664 18686 22744 18692
rect 22744 18634 22796 18640
rect 22756 18426 22784 18634
rect 23124 18426 23152 18770
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 21928 17746 21956 18022
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 22296 17610 22324 18022
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22756 17338 22784 17614
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22940 16182 22968 16594
rect 23124 16425 23152 16934
rect 23110 16416 23166 16425
rect 23110 16351 23166 16360
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22480 16046 22508 16118
rect 23308 16046 23336 17478
rect 23400 17338 23428 17682
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23400 16794 23428 17274
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22664 15570 22692 15846
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 22664 15162 22692 15506
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 20824 14074 20852 14486
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20640 11830 20668 13942
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20916 13394 20944 13670
rect 21008 13530 21036 14350
rect 21836 13938 21864 14758
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 12986 20944 13330
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21008 12238 21036 13262
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12374 21128 12582
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20456 11354 20484 11630
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20640 11286 20668 11766
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 21008 11218 21036 12174
rect 21100 11354 21128 12310
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11694 21312 12174
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10674 19564 10950
rect 20088 10742 20116 11154
rect 21284 10810 21312 11222
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19996 10266 20024 10610
rect 21652 10606 21680 11086
rect 21744 10674 21772 11494
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21652 10266 21680 10542
rect 21744 10266 21772 10610
rect 21836 10305 21864 11630
rect 21822 10296 21878 10305
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21732 10260 21784 10266
rect 21822 10231 21878 10240
rect 21732 10202 21784 10208
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 19168 9586 19196 10066
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19444 8362 19472 9522
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19996 8537 20024 9318
rect 20180 9178 20208 9454
rect 21468 9382 21496 10066
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8634 20116 8978
rect 20904 8968 20956 8974
rect 21468 8945 21496 9318
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 20904 8910 20956 8916
rect 21454 8936 21510 8945
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19982 8528 20038 8537
rect 19982 8463 20038 8472
rect 20916 8362 20944 8910
rect 21454 8871 21510 8880
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 19168 7818 19196 8298
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19444 7546 19472 7890
rect 20732 7818 20760 8298
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19444 6866 19472 7482
rect 19812 7342 19840 7686
rect 21100 7410 21128 7958
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 19800 7336 19852 7342
rect 19852 7296 19932 7324
rect 19800 7278 19852 7284
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19904 6934 19932 7296
rect 19892 6928 19944 6934
rect 19892 6870 19944 6876
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6254 19380 6598
rect 19444 6458 19472 6802
rect 21100 6458 21128 6870
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 20364 5370 20392 6394
rect 21376 6118 21404 6734
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 20534 5672 20590 5681
rect 20534 5607 20590 5616
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20364 5030 20392 5306
rect 20548 5234 20576 5607
rect 21376 5302 21404 6054
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 20548 4826 20576 5170
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21376 3058 21404 3538
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 21468 2650 21496 8871
rect 21652 8634 21680 8978
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21652 6934 21680 7754
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21744 7274 21772 7686
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21560 5370 21588 5714
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21744 5234 21772 7210
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21836 5114 21864 10231
rect 21928 5370 21956 14894
rect 22020 13190 22048 14962
rect 23308 14550 23336 15982
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23400 15162 23428 15438
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23400 14890 23428 15098
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23296 14544 23348 14550
rect 23216 14504 23296 14532
rect 23216 14074 23244 14504
rect 23296 14486 23348 14492
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23308 14074 23336 14350
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13462 22232 13738
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22020 12714 22048 13126
rect 22204 12850 22232 13262
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 22020 11694 22048 12650
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 22020 10062 22048 11630
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22020 9722 22048 9998
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22112 6254 22140 12718
rect 22204 12442 22232 12786
rect 22756 12782 22784 13670
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22848 12986 22876 13398
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 23216 12374 23244 14010
rect 23308 12850 23336 14010
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 11354 23060 12174
rect 23216 11898 23244 12310
rect 23400 11898 23428 14826
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23400 11626 23428 11834
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23400 10810 23428 11154
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 10130 22692 10406
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22664 9722 22692 10066
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 23492 9518 23520 15030
rect 23584 14618 23612 20488
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23664 19304 23716 19310
rect 23768 19281 23796 19314
rect 23664 19246 23716 19252
rect 23754 19272 23810 19281
rect 23676 18970 23704 19246
rect 23754 19207 23810 19216
rect 23938 19272 23994 19281
rect 23938 19207 23994 19216
rect 23952 19174 23980 19207
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 23952 17338 23980 18022
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 23952 17134 23980 17274
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 15026 23796 15302
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23860 11014 23888 11698
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8634 22784 8978
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22940 8022 22968 9318
rect 23124 8634 23152 9318
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23584 8362 23612 10474
rect 23860 10266 23888 10950
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23860 9518 23888 9862
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23768 9217 23796 9454
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23754 9208 23810 9217
rect 23754 9143 23810 9152
rect 23860 8498 23888 9318
rect 24044 9042 24072 28920
rect 24124 28902 24176 28908
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 24228 28490 24256 28698
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24308 28484 24360 28490
rect 24308 28426 24360 28432
rect 24320 28014 24348 28426
rect 24504 28082 24532 28494
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 24308 28008 24360 28014
rect 24308 27950 24360 27956
rect 24136 27849 24164 27950
rect 24122 27840 24178 27849
rect 24122 27775 24178 27784
rect 24320 27674 24348 27950
rect 24308 27668 24360 27674
rect 24308 27610 24360 27616
rect 24872 27538 24900 31300
rect 24952 31282 25004 31288
rect 24952 30796 25004 30802
rect 24952 30738 25004 30744
rect 24964 30054 24992 30738
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24872 26994 24900 27474
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24872 26897 24900 26930
rect 24858 26888 24914 26897
rect 24858 26823 24914 26832
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24780 26042 24808 26386
rect 24768 26036 24820 26042
rect 24768 25978 24820 25984
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 24136 21457 24164 23530
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24412 22710 24440 23054
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 24320 22166 24348 22442
rect 24308 22160 24360 22166
rect 24308 22102 24360 22108
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24122 21448 24178 21457
rect 24122 21383 24178 21392
rect 24228 21146 24256 21966
rect 24320 21690 24348 22102
rect 24412 22030 24440 22646
rect 24504 22506 24532 23054
rect 24780 23050 24808 25978
rect 24964 25809 24992 29990
rect 25044 26920 25096 26926
rect 25044 26862 25096 26868
rect 25056 26081 25084 26862
rect 25042 26072 25098 26081
rect 25042 26007 25098 26016
rect 24950 25800 25006 25809
rect 24950 25735 25006 25744
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 25056 24886 25084 25366
rect 25148 24954 25176 25706
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25148 24682 25176 24890
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24964 23798 24992 24142
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24964 23322 24992 23734
rect 25240 23474 25268 37130
rect 25332 36922 25360 37266
rect 25700 37262 25728 37674
rect 25688 37256 25740 37262
rect 25688 37198 25740 37204
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25332 32978 25360 36858
rect 25964 36644 26016 36650
rect 25964 36586 26016 36592
rect 25976 36378 26004 36586
rect 25964 36372 26016 36378
rect 25964 36314 26016 36320
rect 25976 35562 26004 36314
rect 25872 35556 25924 35562
rect 25872 35498 25924 35504
rect 25964 35556 26016 35562
rect 25964 35498 26016 35504
rect 25884 34950 25912 35498
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25872 34944 25924 34950
rect 25872 34886 25924 34892
rect 25608 34474 25636 34886
rect 25596 34468 25648 34474
rect 25596 34410 25648 34416
rect 25608 34105 25636 34410
rect 25594 34096 25650 34105
rect 25594 34031 25650 34040
rect 25884 33658 25912 34886
rect 26068 34048 26096 39850
rect 27080 39030 27108 40072
rect 27172 39574 27200 40394
rect 27356 40186 27384 40530
rect 27344 40180 27396 40186
rect 27344 40122 27396 40128
rect 27632 39846 27660 41006
rect 27908 40730 27936 41550
rect 28000 41274 28028 41686
rect 27988 41268 28040 41274
rect 27988 41210 28040 41216
rect 27896 40724 27948 40730
rect 27896 40666 27948 40672
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 27436 39840 27488 39846
rect 27436 39782 27488 39788
rect 27620 39840 27672 39846
rect 27620 39782 27672 39788
rect 27160 39568 27212 39574
rect 27160 39510 27212 39516
rect 27172 39098 27200 39510
rect 27252 39500 27304 39506
rect 27252 39442 27304 39448
rect 27160 39092 27212 39098
rect 27160 39034 27212 39040
rect 27068 39024 27120 39030
rect 27068 38966 27120 38972
rect 26148 38752 26200 38758
rect 26148 38694 26200 38700
rect 26160 38486 26188 38694
rect 26148 38480 26200 38486
rect 26148 38422 26200 38428
rect 26608 38480 26660 38486
rect 26608 38422 26660 38428
rect 26160 37738 26188 38422
rect 26240 38276 26292 38282
rect 26240 38218 26292 38224
rect 26148 37732 26200 37738
rect 26148 37674 26200 37680
rect 26252 36786 26280 38218
rect 26620 38010 26648 38422
rect 26976 38344 27028 38350
rect 26976 38286 27028 38292
rect 26988 38010 27016 38286
rect 27080 38010 27108 38966
rect 27264 38826 27292 39442
rect 27448 38894 27476 39782
rect 27724 39642 27752 39986
rect 27712 39636 27764 39642
rect 27712 39578 27764 39584
rect 27436 38888 27488 38894
rect 27436 38830 27488 38836
rect 27896 38888 27948 38894
rect 27896 38830 27948 38836
rect 27252 38820 27304 38826
rect 27252 38762 27304 38768
rect 27908 38321 27936 38830
rect 27894 38312 27950 38321
rect 27894 38247 27950 38256
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 26976 38004 27028 38010
rect 26976 37946 27028 37952
rect 27068 38004 27120 38010
rect 27068 37946 27120 37952
rect 27620 38004 27672 38010
rect 27620 37946 27672 37952
rect 26792 37936 26844 37942
rect 26792 37878 26844 37884
rect 26804 37330 26832 37878
rect 27632 37806 27660 37946
rect 27620 37800 27672 37806
rect 27620 37742 27672 37748
rect 26884 37732 26936 37738
rect 26884 37674 26936 37680
rect 26792 37324 26844 37330
rect 26792 37266 26844 37272
rect 26332 37120 26384 37126
rect 26332 37062 26384 37068
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26160 36038 26188 36722
rect 26252 36106 26280 36722
rect 26344 36310 26372 37062
rect 26804 36922 26832 37266
rect 26792 36916 26844 36922
rect 26792 36858 26844 36864
rect 26896 36786 26924 37674
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 26884 36780 26936 36786
rect 26884 36722 26936 36728
rect 26332 36304 26384 36310
rect 26332 36246 26384 36252
rect 26792 36304 26844 36310
rect 26792 36246 26844 36252
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26160 35834 26188 35974
rect 26148 35828 26200 35834
rect 26148 35770 26200 35776
rect 26344 35290 26372 36246
rect 26804 35816 26832 36246
rect 26896 36174 26924 36722
rect 27724 36582 27752 37198
rect 28092 36922 28120 42570
rect 28368 42226 28396 42706
rect 28356 42220 28408 42226
rect 28356 42162 28408 42168
rect 28460 41206 28488 42774
rect 28644 42362 28672 43386
rect 28736 42702 28764 45426
rect 29012 45014 29040 45902
rect 30208 45490 30236 46106
rect 30380 46028 30432 46034
rect 30380 45970 30432 45976
rect 31208 46028 31260 46034
rect 31208 45970 31260 45976
rect 30392 45626 30420 45970
rect 30380 45620 30432 45626
rect 30380 45562 30432 45568
rect 29368 45484 29420 45490
rect 29368 45426 29420 45432
rect 30196 45484 30248 45490
rect 30196 45426 30248 45432
rect 29380 45082 29408 45426
rect 30196 45348 30248 45354
rect 30196 45290 30248 45296
rect 29368 45076 29420 45082
rect 29368 45018 29420 45024
rect 29000 45008 29052 45014
rect 29000 44950 29052 44956
rect 29012 43926 29040 44950
rect 30208 44266 30236 45290
rect 30392 45082 30420 45562
rect 31220 45286 31248 45970
rect 31312 45286 31340 49558
rect 43626 49558 43760 49586
rect 43626 49520 43682 49558
rect 41052 47116 41104 47122
rect 41052 47058 41104 47064
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 41064 46646 41092 47058
rect 41512 46912 41564 46918
rect 41512 46854 41564 46860
rect 36084 46640 36136 46646
rect 36084 46582 36136 46588
rect 41052 46640 41104 46646
rect 41052 46582 41104 46588
rect 34704 46368 34756 46374
rect 34704 46310 34756 46316
rect 34152 46096 34204 46102
rect 34152 46038 34204 46044
rect 32864 45824 32916 45830
rect 32864 45766 32916 45772
rect 33324 45824 33376 45830
rect 33324 45766 33376 45772
rect 32876 45422 32904 45766
rect 32864 45416 32916 45422
rect 32864 45358 32916 45364
rect 31208 45280 31260 45286
rect 31208 45222 31260 45228
rect 31300 45280 31352 45286
rect 31300 45222 31352 45228
rect 32220 45280 32272 45286
rect 32220 45222 32272 45228
rect 30380 45076 30432 45082
rect 30380 45018 30432 45024
rect 31220 44946 31248 45222
rect 30380 44940 30432 44946
rect 30380 44882 30432 44888
rect 31208 44940 31260 44946
rect 31208 44882 31260 44888
rect 30392 44538 30420 44882
rect 30748 44872 30800 44878
rect 30748 44814 30800 44820
rect 30380 44532 30432 44538
rect 30380 44474 30432 44480
rect 30196 44260 30248 44266
rect 30196 44202 30248 44208
rect 30208 43926 30236 44202
rect 29000 43920 29052 43926
rect 29000 43862 29052 43868
rect 30196 43920 30248 43926
rect 30196 43862 30248 43868
rect 29012 43314 29040 43862
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 29644 43308 29696 43314
rect 29644 43250 29696 43256
rect 29656 42838 29684 43250
rect 30208 43110 30236 43862
rect 30392 43382 30420 44474
rect 30760 43858 30788 44814
rect 30840 44396 30892 44402
rect 30840 44338 30892 44344
rect 30748 43852 30800 43858
rect 30748 43794 30800 43800
rect 30760 43450 30788 43794
rect 30748 43444 30800 43450
rect 30748 43386 30800 43392
rect 30380 43376 30432 43382
rect 30380 43318 30432 43324
rect 30196 43104 30248 43110
rect 30196 43046 30248 43052
rect 30208 42838 30236 43046
rect 28816 42832 28868 42838
rect 28816 42774 28868 42780
rect 29644 42832 29696 42838
rect 29644 42774 29696 42780
rect 30196 42832 30248 42838
rect 30196 42774 30248 42780
rect 28724 42696 28776 42702
rect 28724 42638 28776 42644
rect 28632 42356 28684 42362
rect 28632 42298 28684 42304
rect 28736 41818 28764 42638
rect 28828 42566 28856 42774
rect 28816 42560 28868 42566
rect 28816 42502 28868 42508
rect 29092 42560 29144 42566
rect 29092 42502 29144 42508
rect 29104 42362 29132 42502
rect 29092 42356 29144 42362
rect 29092 42298 29144 42304
rect 28816 42016 28868 42022
rect 28816 41958 28868 41964
rect 28724 41812 28776 41818
rect 28724 41754 28776 41760
rect 28448 41200 28500 41206
rect 28448 41142 28500 41148
rect 28540 40996 28592 41002
rect 28540 40938 28592 40944
rect 28552 40730 28580 40938
rect 28540 40724 28592 40730
rect 28540 40666 28592 40672
rect 28552 40186 28580 40666
rect 28828 40633 28856 41958
rect 29552 41744 29604 41750
rect 29552 41686 29604 41692
rect 29460 41608 29512 41614
rect 29460 41550 29512 41556
rect 29472 41138 29500 41550
rect 29564 41274 29592 41686
rect 29656 41614 29684 42774
rect 30208 42022 30236 42774
rect 30748 42696 30800 42702
rect 30748 42638 30800 42644
rect 30760 42022 30788 42638
rect 30196 42016 30248 42022
rect 30196 41958 30248 41964
rect 30748 42016 30800 42022
rect 30748 41958 30800 41964
rect 29644 41608 29696 41614
rect 29644 41550 29696 41556
rect 29552 41268 29604 41274
rect 29552 41210 29604 41216
rect 29460 41132 29512 41138
rect 29460 41074 29512 41080
rect 29564 40730 29592 41210
rect 30208 41002 30236 41958
rect 30760 41818 30788 41958
rect 30748 41812 30800 41818
rect 30748 41754 30800 41760
rect 30564 41064 30616 41070
rect 30564 41006 30616 41012
rect 30196 40996 30248 41002
rect 30196 40938 30248 40944
rect 30576 40730 30604 41006
rect 29552 40724 29604 40730
rect 29552 40666 29604 40672
rect 30564 40724 30616 40730
rect 30564 40666 30616 40672
rect 28814 40624 28870 40633
rect 28814 40559 28870 40568
rect 30564 40588 30616 40594
rect 30564 40530 30616 40536
rect 28908 40520 28960 40526
rect 28908 40462 28960 40468
rect 29826 40488 29882 40497
rect 28920 40186 28948 40462
rect 29826 40423 29882 40432
rect 28540 40180 28592 40186
rect 28540 40122 28592 40128
rect 28908 40180 28960 40186
rect 28908 40122 28960 40128
rect 28552 39642 28580 40122
rect 28540 39636 28592 39642
rect 28540 39578 28592 39584
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 28172 38888 28224 38894
rect 28172 38830 28224 38836
rect 28184 38214 28212 38830
rect 28276 38554 28304 39374
rect 28552 39098 28580 39578
rect 28632 39296 28684 39302
rect 28632 39238 28684 39244
rect 29184 39296 29236 39302
rect 29184 39238 29236 39244
rect 29460 39296 29512 39302
rect 29460 39238 29512 39244
rect 28540 39092 28592 39098
rect 28540 39034 28592 39040
rect 28356 38956 28408 38962
rect 28356 38898 28408 38904
rect 28264 38548 28316 38554
rect 28264 38490 28316 38496
rect 28172 38208 28224 38214
rect 28172 38150 28224 38156
rect 28184 37806 28212 38150
rect 28276 37874 28304 38490
rect 28368 38350 28396 38898
rect 28540 38820 28592 38826
rect 28540 38762 28592 38768
rect 28552 38350 28580 38762
rect 28356 38344 28408 38350
rect 28356 38286 28408 38292
rect 28540 38344 28592 38350
rect 28540 38286 28592 38292
rect 28264 37868 28316 37874
rect 28264 37810 28316 37816
rect 28172 37800 28224 37806
rect 28172 37742 28224 37748
rect 28184 37466 28212 37742
rect 28172 37460 28224 37466
rect 28172 37402 28224 37408
rect 28368 37262 28396 38286
rect 28552 37466 28580 38286
rect 28540 37460 28592 37466
rect 28540 37402 28592 37408
rect 28448 37392 28500 37398
rect 28448 37334 28500 37340
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28080 36916 28132 36922
rect 28080 36858 28132 36864
rect 28092 36718 28120 36858
rect 28080 36712 28132 36718
rect 28080 36654 28132 36660
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 27160 36032 27212 36038
rect 27160 35974 27212 35980
rect 26884 35828 26936 35834
rect 26804 35788 26884 35816
rect 26884 35770 26936 35776
rect 26896 35737 26924 35770
rect 26882 35728 26938 35737
rect 26882 35663 26938 35672
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26884 34468 26936 34474
rect 26884 34410 26936 34416
rect 26700 34400 26752 34406
rect 26700 34342 26752 34348
rect 26608 34128 26660 34134
rect 26608 34070 26660 34076
rect 25976 34020 26096 34048
rect 25872 33652 25924 33658
rect 25872 33594 25924 33600
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 25332 32502 25360 32914
rect 25412 32768 25464 32774
rect 25412 32710 25464 32716
rect 25320 32496 25372 32502
rect 25320 32438 25372 32444
rect 25424 32366 25452 32710
rect 25412 32360 25464 32366
rect 25412 32302 25464 32308
rect 25412 31952 25464 31958
rect 25412 31894 25464 31900
rect 25424 31482 25452 31894
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25688 31204 25740 31210
rect 25688 31146 25740 31152
rect 25700 30394 25728 31146
rect 25688 30388 25740 30394
rect 25688 30330 25740 30336
rect 25872 29028 25924 29034
rect 25872 28970 25924 28976
rect 25884 28762 25912 28970
rect 25872 28756 25924 28762
rect 25872 28698 25924 28704
rect 25412 28416 25464 28422
rect 25412 28358 25464 28364
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25332 24818 25360 26318
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25332 24410 25360 24754
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 25424 24342 25452 28358
rect 25688 28008 25740 28014
rect 25688 27950 25740 27956
rect 25700 27606 25728 27950
rect 25688 27600 25740 27606
rect 25688 27542 25740 27548
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25516 26926 25544 27406
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25516 26450 25544 26862
rect 25504 26444 25556 26450
rect 25504 26386 25556 26392
rect 25516 25498 25544 26386
rect 25608 25906 25636 26930
rect 25596 25900 25648 25906
rect 25596 25842 25648 25848
rect 25608 25498 25636 25842
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25608 24818 25636 25230
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 25424 23866 25452 24278
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25884 23866 25912 24142
rect 25412 23860 25464 23866
rect 25872 23860 25924 23866
rect 25412 23802 25464 23808
rect 25792 23820 25872 23848
rect 25148 23446 25268 23474
rect 25424 23474 25452 23802
rect 25424 23446 25636 23474
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24872 22817 24900 23122
rect 24858 22808 24914 22817
rect 25056 22778 25084 23122
rect 24858 22743 24914 22752
rect 25044 22772 25096 22778
rect 24872 22642 24900 22743
rect 25044 22714 25096 22720
rect 25056 22681 25084 22714
rect 25042 22672 25098 22681
rect 24860 22636 24912 22642
rect 25042 22607 25098 22616
rect 24860 22578 24912 22584
rect 24492 22500 24544 22506
rect 24492 22442 24544 22448
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24308 21684 24360 21690
rect 24308 21626 24360 21632
rect 24504 21554 24532 22442
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 25148 20398 25176 23446
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25424 22506 25452 22986
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25412 22500 25464 22506
rect 25412 22442 25464 22448
rect 25424 22166 25452 22442
rect 25516 22234 25544 22918
rect 25608 22506 25636 23446
rect 25792 22710 25820 23820
rect 25872 23802 25924 23808
rect 25976 23474 26004 34020
rect 26054 33688 26110 33697
rect 26054 33623 26110 33632
rect 26068 33454 26096 33623
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 26068 28082 26096 33390
rect 26620 33386 26648 34070
rect 26712 33998 26740 34342
rect 26896 33998 26924 34410
rect 26700 33992 26752 33998
rect 26700 33934 26752 33940
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26608 33380 26660 33386
rect 26608 33322 26660 33328
rect 26608 33108 26660 33114
rect 26712 33096 26740 33934
rect 26792 33516 26844 33522
rect 26792 33458 26844 33464
rect 26660 33068 26740 33096
rect 26608 33050 26660 33056
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26160 32570 26188 32710
rect 26804 32570 26832 33458
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26792 32564 26844 32570
rect 26792 32506 26844 32512
rect 26896 31822 26924 33934
rect 27068 33040 27120 33046
rect 27068 32982 27120 32988
rect 27080 32570 27108 32982
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 27068 32224 27120 32230
rect 27172 32212 27200 35974
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 27264 34610 27292 35090
rect 27724 34678 27752 36518
rect 27816 36378 27844 36518
rect 27804 36372 27856 36378
rect 27804 36314 27856 36320
rect 27816 35698 27844 36314
rect 27804 35692 27856 35698
rect 27804 35634 27856 35640
rect 28092 35601 28120 36654
rect 28078 35592 28134 35601
rect 28368 35562 28396 37198
rect 28460 36582 28488 37334
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28078 35527 28134 35536
rect 28356 35556 28408 35562
rect 27804 34944 27856 34950
rect 27804 34886 27856 34892
rect 27816 34746 27844 34886
rect 27804 34740 27856 34746
rect 27804 34682 27856 34688
rect 27712 34672 27764 34678
rect 27712 34614 27764 34620
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 28092 34406 28120 35527
rect 28356 35498 28408 35504
rect 28262 35320 28318 35329
rect 28262 35255 28318 35264
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33522 27568 33798
rect 28184 33658 28212 33934
rect 28172 33652 28224 33658
rect 28172 33594 28224 33600
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27436 33380 27488 33386
rect 27436 33322 27488 33328
rect 27448 32910 27476 33322
rect 28184 33134 28212 33594
rect 28092 33106 28212 33134
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27528 32768 27580 32774
rect 27528 32710 27580 32716
rect 27540 32298 27568 32710
rect 27724 32298 27752 32846
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27712 32292 27764 32298
rect 27712 32234 27764 32240
rect 27120 32184 27200 32212
rect 27068 32166 27120 32172
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26240 31204 26292 31210
rect 26240 31146 26292 31152
rect 26252 30598 26280 31146
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26712 30870 26740 31078
rect 26896 30870 26924 31758
rect 26700 30864 26752 30870
rect 26700 30806 26752 30812
rect 26884 30864 26936 30870
rect 26884 30806 26936 30812
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26148 30116 26200 30122
rect 26148 30058 26200 30064
rect 26160 28694 26188 30058
rect 26252 28762 26280 30534
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 26344 29510 26372 30126
rect 26896 29646 26924 30806
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26344 29170 26372 29446
rect 26896 29170 26924 29582
rect 27080 29186 27108 32166
rect 27448 32026 27476 32234
rect 27436 32020 27488 32026
rect 27436 31962 27488 31968
rect 27448 31482 27476 31962
rect 27540 31890 27568 32234
rect 28092 31958 28120 33106
rect 28080 31952 28132 31958
rect 28080 31894 28132 31900
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27436 31476 27488 31482
rect 27436 31418 27488 31424
rect 28276 31414 28304 35255
rect 28460 35222 28488 36518
rect 28540 36304 28592 36310
rect 28540 36246 28592 36252
rect 28552 35766 28580 36246
rect 28540 35760 28592 35766
rect 28540 35702 28592 35708
rect 28448 35216 28500 35222
rect 28448 35158 28500 35164
rect 28460 34728 28488 35158
rect 28460 34700 28580 34728
rect 28552 34610 28580 34700
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28460 34513 28488 34546
rect 28644 34542 28672 39238
rect 29196 39098 29224 39238
rect 28724 39092 28776 39098
rect 28724 39034 28776 39040
rect 29184 39092 29236 39098
rect 29184 39034 29236 39040
rect 28736 38486 28764 39034
rect 29196 38758 29224 39034
rect 29472 38962 29500 39238
rect 29460 38956 29512 38962
rect 29460 38898 29512 38904
rect 29644 38956 29696 38962
rect 29644 38898 29696 38904
rect 29184 38752 29236 38758
rect 29184 38694 29236 38700
rect 28724 38480 28776 38486
rect 28724 38422 28776 38428
rect 28736 38010 28764 38422
rect 29460 38208 29512 38214
rect 29460 38150 29512 38156
rect 28724 38004 28776 38010
rect 28724 37946 28776 37952
rect 29184 37800 29236 37806
rect 29236 37760 29316 37788
rect 29184 37742 29236 37748
rect 29288 37466 29316 37760
rect 29472 37738 29500 38150
rect 29656 38010 29684 38898
rect 29644 38004 29696 38010
rect 29644 37946 29696 37952
rect 29368 37732 29420 37738
rect 29368 37674 29420 37680
rect 29460 37732 29512 37738
rect 29460 37674 29512 37680
rect 29276 37460 29328 37466
rect 29276 37402 29328 37408
rect 29380 37126 29408 37674
rect 29840 37330 29868 40423
rect 30576 39846 30604 40530
rect 30852 39846 30880 44338
rect 31220 43654 31248 44882
rect 31312 43994 31340 45222
rect 32232 45082 32260 45222
rect 32220 45076 32272 45082
rect 32220 45018 32272 45024
rect 32876 45014 32904 45358
rect 32864 45008 32916 45014
rect 32864 44950 32916 44956
rect 32128 44940 32180 44946
rect 32128 44882 32180 44888
rect 32220 44940 32272 44946
rect 32220 44882 32272 44888
rect 31392 44736 31444 44742
rect 31392 44678 31444 44684
rect 31404 44402 31432 44678
rect 31392 44396 31444 44402
rect 31392 44338 31444 44344
rect 32140 43994 32168 44882
rect 32232 44538 32260 44882
rect 33336 44538 33364 45766
rect 34164 45354 34192 46038
rect 34716 45626 34744 46310
rect 35624 46028 35676 46034
rect 35624 45970 35676 45976
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34704 45620 34756 45626
rect 34704 45562 34756 45568
rect 34152 45348 34204 45354
rect 34152 45290 34204 45296
rect 35256 45348 35308 45354
rect 35256 45290 35308 45296
rect 33416 45280 33468 45286
rect 33416 45222 33468 45228
rect 32220 44532 32272 44538
rect 32220 44474 32272 44480
rect 33324 44532 33376 44538
rect 33324 44474 33376 44480
rect 31300 43988 31352 43994
rect 31300 43930 31352 43936
rect 32128 43988 32180 43994
rect 32128 43930 32180 43936
rect 30932 43648 30984 43654
rect 30932 43590 30984 43596
rect 31208 43648 31260 43654
rect 31208 43590 31260 43596
rect 30944 43178 30972 43590
rect 30932 43172 30984 43178
rect 30932 43114 30984 43120
rect 31220 42158 31248 43590
rect 32232 43314 32260 44474
rect 32956 44328 33008 44334
rect 32956 44270 33008 44276
rect 32968 43897 32996 44270
rect 33428 43994 33456 45222
rect 34164 45014 34192 45290
rect 34152 45008 34204 45014
rect 34152 44950 34204 44956
rect 34796 45008 34848 45014
rect 34796 44950 34848 44956
rect 34060 44872 34112 44878
rect 34060 44814 34112 44820
rect 34072 44538 34100 44814
rect 34060 44532 34112 44538
rect 34060 44474 34112 44480
rect 33416 43988 33468 43994
rect 33416 43930 33468 43936
rect 32954 43888 33010 43897
rect 32954 43823 33010 43832
rect 32220 43308 32272 43314
rect 32220 43250 32272 43256
rect 32036 43240 32088 43246
rect 32036 43182 32088 43188
rect 31208 42152 31260 42158
rect 31208 42094 31260 42100
rect 31220 41818 31248 42094
rect 31208 41812 31260 41818
rect 31208 41754 31260 41760
rect 31392 41676 31444 41682
rect 31392 41618 31444 41624
rect 31404 40934 31432 41618
rect 31392 40928 31444 40934
rect 31392 40870 31444 40876
rect 31404 40594 31432 40870
rect 31392 40588 31444 40594
rect 31392 40530 31444 40536
rect 31404 39982 31432 40530
rect 30932 39976 30984 39982
rect 30932 39918 30984 39924
rect 31392 39976 31444 39982
rect 31392 39918 31444 39924
rect 30196 39840 30248 39846
rect 30196 39782 30248 39788
rect 30564 39840 30616 39846
rect 30564 39782 30616 39788
rect 30840 39840 30892 39846
rect 30840 39782 30892 39788
rect 30208 39574 30236 39782
rect 30196 39568 30248 39574
rect 30196 39510 30248 39516
rect 30288 38820 30340 38826
rect 30288 38762 30340 38768
rect 30300 38486 30328 38762
rect 30288 38480 30340 38486
rect 30288 38422 30340 38428
rect 30380 38480 30432 38486
rect 30380 38422 30432 38428
rect 30392 38010 30420 38422
rect 30472 38276 30524 38282
rect 30472 38218 30524 38224
rect 30380 38004 30432 38010
rect 30380 37946 30432 37952
rect 29828 37324 29880 37330
rect 29828 37266 29880 37272
rect 29368 37120 29420 37126
rect 29368 37062 29420 37068
rect 28908 36168 28960 36174
rect 28960 36128 29040 36156
rect 28908 36110 28960 36116
rect 29012 35494 29040 36128
rect 29380 36106 29408 37062
rect 29840 36922 29868 37266
rect 30484 37126 30512 38218
rect 30576 37670 30604 39782
rect 30944 39642 30972 39918
rect 30932 39636 30984 39642
rect 30932 39578 30984 39584
rect 30944 39302 30972 39578
rect 31404 39574 31432 39918
rect 31392 39568 31444 39574
rect 31392 39510 31444 39516
rect 31024 39500 31076 39506
rect 31024 39442 31076 39448
rect 30932 39296 30984 39302
rect 30932 39238 30984 39244
rect 31036 39098 31064 39442
rect 31024 39092 31076 39098
rect 31076 39052 31156 39080
rect 31024 39034 31076 39040
rect 30564 37664 30616 37670
rect 30564 37606 30616 37612
rect 31024 37324 31076 37330
rect 31024 37266 31076 37272
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 29748 36378 29776 36586
rect 29736 36372 29788 36378
rect 29736 36314 29788 36320
rect 29368 36100 29420 36106
rect 29368 36042 29420 36048
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 29012 34746 29040 35430
rect 29380 35222 29408 36042
rect 29748 35834 29776 36314
rect 29840 36038 29868 36858
rect 30300 36310 30328 37062
rect 30484 36786 30512 37062
rect 30472 36780 30524 36786
rect 30472 36722 30524 36728
rect 30288 36304 30340 36310
rect 30288 36246 30340 36252
rect 30380 36304 30432 36310
rect 30380 36246 30432 36252
rect 29828 36032 29880 36038
rect 29828 35974 29880 35980
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29748 35329 29776 35566
rect 29734 35320 29790 35329
rect 30300 35290 30328 36246
rect 30392 35834 30420 36246
rect 30484 36174 30512 36722
rect 30932 36644 30984 36650
rect 30932 36586 30984 36592
rect 30944 36242 30972 36586
rect 31036 36582 31064 37266
rect 31128 37194 31156 39052
rect 31208 38344 31260 38350
rect 31208 38286 31260 38292
rect 31220 37806 31248 38286
rect 31208 37800 31260 37806
rect 31208 37742 31260 37748
rect 31300 37800 31352 37806
rect 31300 37742 31352 37748
rect 31312 37466 31340 37742
rect 31300 37460 31352 37466
rect 31220 37420 31300 37448
rect 31116 37188 31168 37194
rect 31116 37130 31168 37136
rect 31024 36576 31076 36582
rect 31024 36518 31076 36524
rect 30932 36236 30984 36242
rect 30932 36178 30984 36184
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 29734 35255 29790 35264
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 29368 35216 29420 35222
rect 29368 35158 29420 35164
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29840 34746 29868 34954
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29828 34740 29880 34746
rect 29828 34682 29880 34688
rect 29552 34672 29604 34678
rect 29552 34614 29604 34620
rect 28632 34536 28684 34542
rect 28446 34504 28502 34513
rect 28632 34478 28684 34484
rect 28446 34439 28502 34448
rect 29092 33924 29144 33930
rect 29092 33866 29144 33872
rect 28632 33040 28684 33046
rect 28632 32982 28684 32988
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28448 32292 28500 32298
rect 28448 32234 28500 32240
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28264 31408 28316 31414
rect 28264 31350 28316 31356
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 30394 27476 30670
rect 27436 30388 27488 30394
rect 27436 30330 27488 30336
rect 27160 30048 27212 30054
rect 27160 29990 27212 29996
rect 27172 29782 27200 29990
rect 27160 29776 27212 29782
rect 27160 29718 27212 29724
rect 27172 29306 27200 29718
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 26884 29164 26936 29170
rect 27080 29158 27200 29186
rect 26884 29106 26936 29112
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26148 28688 26200 28694
rect 26148 28630 26200 28636
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26160 27946 26188 28630
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26148 27940 26200 27946
rect 26148 27882 26200 27888
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 25884 23446 26004 23474
rect 25780 22704 25832 22710
rect 25780 22646 25832 22652
rect 25596 22500 25648 22506
rect 25596 22442 25648 22448
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24964 19514 24992 19858
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24964 18426 24992 19450
rect 25056 18834 25084 20198
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 18358 25084 18770
rect 25148 18426 25176 20334
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25148 18222 25176 18362
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24228 17746 24256 18022
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 16658 24624 17478
rect 25056 17338 25084 17682
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24596 16250 24624 16594
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24228 15094 24256 15506
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24412 14414 24440 14826
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24308 14000 24360 14006
rect 24308 13942 24360 13948
rect 24320 13734 24348 13942
rect 24492 13796 24544 13802
rect 24492 13738 24544 13744
rect 24308 13728 24360 13734
rect 24308 13670 24360 13676
rect 24504 13530 24532 13738
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24504 12170 24532 13466
rect 24596 12986 24624 14826
rect 24780 13394 24808 14894
rect 24872 14890 24900 15506
rect 24860 14884 24912 14890
rect 24860 14826 24912 14832
rect 24964 14550 24992 17002
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25240 16114 25268 16390
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25240 15638 25268 16050
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 14958 25268 15302
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24872 14074 24900 14350
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24964 14006 24992 14486
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24596 12782 24624 12922
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24504 11762 24532 12106
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24492 11552 24544 11558
rect 24596 11540 24624 12242
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24688 11762 24716 12038
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24544 11512 24624 11540
rect 24492 11494 24544 11500
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23676 8090 23704 8230
rect 23860 8090 23888 8434
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 22928 8016 22980 8022
rect 22928 7958 22980 7964
rect 23952 7954 23980 8774
rect 24044 8566 24072 8978
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22664 7546 22692 7822
rect 23952 7546 23980 7890
rect 24136 7546 24164 9454
rect 24228 9178 24256 10066
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24136 7342 24164 7482
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22388 6322 22416 6598
rect 22480 6390 22508 7142
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21928 5166 21956 5306
rect 21744 5086 21864 5114
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21744 4214 21772 5086
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21744 4078 21772 4150
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22020 3398 22048 4014
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 22020 2446 22048 3334
rect 22112 3097 22140 5102
rect 22296 4865 22324 6190
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 5234 22416 5646
rect 22480 5574 22508 6190
rect 23124 6118 23152 6870
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5846 23152 6054
rect 23112 5840 23164 5846
rect 23112 5782 23164 5788
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22282 4856 22338 4865
rect 22388 4826 22416 5170
rect 22480 5166 22508 5510
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22282 4791 22338 4800
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22480 4486 22508 5102
rect 23124 5030 23152 5782
rect 23400 5778 23428 6598
rect 23768 6322 23796 6598
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23768 5234 23796 5510
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 4078 22508 4422
rect 22940 4282 22968 4626
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22836 4004 22888 4010
rect 22836 3946 22888 3952
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22572 3194 22600 3878
rect 22848 3534 22876 3946
rect 22940 3738 22968 4218
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23020 3664 23072 3670
rect 23124 3652 23152 4966
rect 23664 4820 23716 4826
rect 23768 4808 23796 5170
rect 23860 5098 23888 5306
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23716 4780 23796 4808
rect 23664 4762 23716 4768
rect 23952 4758 23980 6122
rect 24412 5846 24440 7346
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 4826 24256 5646
rect 24412 5370 24440 5782
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24412 4758 24440 5170
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23400 3942 23428 4558
rect 23952 4214 23980 4694
rect 24504 4604 24532 11494
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24596 10470 24624 11086
rect 24780 10674 24808 12378
rect 24872 12306 24900 12582
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24964 12102 24992 13262
rect 25148 12986 25176 13466
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24596 10266 24624 10406
rect 24780 10266 24808 10610
rect 24964 10538 24992 11290
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24872 9489 24900 10134
rect 24858 9480 24914 9489
rect 24858 9415 24914 9424
rect 24872 9382 24900 9415
rect 24860 9376 24912 9382
rect 24780 9336 24860 9364
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24596 5030 24624 7142
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24688 6118 24716 6802
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5914 24716 6054
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24596 4758 24624 4966
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24412 4576 24532 4604
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 24412 4078 24440 4576
rect 24596 4536 24624 4694
rect 24504 4508 24624 4536
rect 24504 4078 24532 4508
rect 24688 4468 24716 5306
rect 24596 4440 24716 4468
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 24412 3777 24440 4014
rect 24398 3768 24454 3777
rect 24398 3703 24454 3712
rect 24596 3670 24624 4440
rect 24780 4154 24808 9336
rect 24860 9318 24912 9324
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24964 8634 24992 8978
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25056 8022 25084 8910
rect 24952 8016 25004 8022
rect 24952 7958 25004 7964
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 24964 7546 24992 7958
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25056 7410 25084 7958
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24872 5846 24900 6258
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 25148 5098 25176 6054
rect 25136 5092 25188 5098
rect 25136 5034 25188 5040
rect 24688 4126 24808 4154
rect 23072 3624 23152 3652
rect 23020 3606 23072 3612
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22098 3088 22154 3097
rect 22098 3023 22154 3032
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22572 2582 22600 2926
rect 22848 2650 22876 3470
rect 23124 3194 23152 3624
rect 24584 3664 24636 3670
rect 24584 3606 24636 3612
rect 24688 3602 24716 4126
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24872 3602 24900 4014
rect 25136 4004 25188 4010
rect 25136 3946 25188 3952
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 2922 23152 3130
rect 24044 2990 24072 3334
rect 24412 3194 24440 3334
rect 24688 3194 24716 3538
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23112 2916 23164 2922
rect 23112 2858 23164 2864
rect 24768 2916 24820 2922
rect 24768 2858 24820 2864
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23400 2582 23428 2790
rect 24780 2582 24808 2858
rect 24872 2650 24900 3538
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24964 3058 24992 3470
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25056 2650 25084 2926
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 25148 2514 25176 3946
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 17774 82 17830 480
rect 17420 54 17830 82
rect 3514 0 3570 54
rect 10598 0 10654 54
rect 17774 0 17830 54
rect 24858 82 24914 480
rect 25240 82 25268 14554
rect 25332 12186 25360 21830
rect 25516 21554 25544 22170
rect 25608 22030 25636 22442
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 21690 25636 21966
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25608 21418 25636 21626
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25884 21010 25912 23446
rect 26068 23186 26096 25842
rect 26344 24313 26372 28018
rect 26436 27538 26464 28902
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26976 28620 27028 28626
rect 26976 28562 27028 28568
rect 26712 27878 26740 28562
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26700 27872 26752 27878
rect 26700 27814 26752 27820
rect 26516 27668 26568 27674
rect 26516 27610 26568 27616
rect 26424 27532 26476 27538
rect 26424 27474 26476 27480
rect 26436 27130 26464 27474
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26436 27033 26464 27066
rect 26422 27024 26478 27033
rect 26422 26959 26478 26968
rect 26528 25362 26556 27610
rect 26516 25356 26568 25362
rect 26516 25298 26568 25304
rect 26528 24954 26556 25298
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26330 24304 26386 24313
rect 26330 24239 26386 24248
rect 26344 24138 26372 24239
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 26344 23866 26372 24074
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26344 23662 26372 23802
rect 26332 23656 26384 23662
rect 26332 23598 26384 23604
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26056 23180 26108 23186
rect 26056 23122 26108 23128
rect 26344 22642 26372 23462
rect 26620 23254 26648 27814
rect 26988 26858 27016 28562
rect 26976 26852 27028 26858
rect 26976 26794 27028 26800
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 26884 25764 26936 25770
rect 26884 25706 26936 25712
rect 26700 25696 26752 25702
rect 26700 25638 26752 25644
rect 26712 24342 26740 25638
rect 26896 25498 26924 25706
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 26884 24608 26936 24614
rect 26884 24550 26936 24556
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26712 23866 26740 24278
rect 26896 23866 26924 24550
rect 26700 23860 26752 23866
rect 26700 23802 26752 23808
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26424 23248 26476 23254
rect 26424 23190 26476 23196
rect 26608 23248 26660 23254
rect 26608 23190 26660 23196
rect 26436 22778 26464 23190
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26988 22234 27016 22578
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 26608 22092 26660 22098
rect 26608 22034 26660 22040
rect 26620 21690 26648 22034
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 27080 21010 27108 26726
rect 27172 26450 27200 29158
rect 28276 28966 28304 29582
rect 28368 29306 28396 31622
rect 28460 31210 28488 32234
rect 28552 31958 28580 32846
rect 28644 32502 28672 32982
rect 29104 32842 29132 33866
rect 29092 32836 29144 32842
rect 29092 32778 29144 32784
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28644 32230 28672 32438
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28540 31952 28592 31958
rect 28540 31894 28592 31900
rect 28632 31884 28684 31890
rect 28632 31826 28684 31832
rect 28448 31204 28500 31210
rect 28448 31146 28500 31152
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28368 29034 28396 29242
rect 28460 29034 28488 31146
rect 28644 31142 28672 31826
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 28644 30977 28672 31078
rect 28630 30968 28686 30977
rect 28630 30903 28686 30912
rect 28644 30326 28672 30903
rect 28632 30320 28684 30326
rect 28632 30262 28684 30268
rect 28736 30054 28764 32166
rect 29104 30734 29132 32778
rect 29276 32360 29328 32366
rect 29276 32302 29328 32308
rect 29288 32026 29316 32302
rect 29276 32020 29328 32026
rect 29276 31962 29328 31968
rect 29368 31136 29420 31142
rect 29368 31078 29420 31084
rect 29184 30864 29236 30870
rect 29184 30806 29236 30812
rect 29092 30728 29144 30734
rect 29092 30670 29144 30676
rect 29196 30190 29224 30806
rect 29380 30258 29408 31078
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29184 30184 29236 30190
rect 29184 30126 29236 30132
rect 29092 30116 29144 30122
rect 29092 30058 29144 30064
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28736 29850 28764 29990
rect 28724 29844 28776 29850
rect 28724 29786 28776 29792
rect 28356 29028 28408 29034
rect 28356 28970 28408 28976
rect 28448 29028 28500 29034
rect 28448 28970 28500 28976
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28276 28762 28304 28902
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 28368 28626 28396 28970
rect 28736 28966 28764 29786
rect 28724 28960 28776 28966
rect 28724 28902 28776 28908
rect 28172 28620 28224 28626
rect 28172 28562 28224 28568
rect 28356 28620 28408 28626
rect 28356 28562 28408 28568
rect 28184 28218 28212 28562
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 28080 27872 28132 27878
rect 28080 27814 28132 27820
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 27172 25838 27200 26386
rect 27528 26240 27580 26246
rect 27528 26182 27580 26188
rect 27160 25832 27212 25838
rect 27160 25774 27212 25780
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27172 24410 27200 24618
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27172 22642 27200 24346
rect 27264 24342 27292 24754
rect 27448 24682 27476 25094
rect 27436 24676 27488 24682
rect 27436 24618 27488 24624
rect 27252 24336 27304 24342
rect 27252 24278 27304 24284
rect 27264 23254 27292 24278
rect 27342 23896 27398 23905
rect 27342 23831 27398 23840
rect 27356 23662 27384 23831
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27252 23248 27304 23254
rect 27356 23225 27384 23598
rect 27434 23352 27490 23361
rect 27434 23287 27490 23296
rect 27252 23190 27304 23196
rect 27342 23216 27398 23225
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27264 22098 27292 23190
rect 27342 23151 27398 23160
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27356 22234 27384 23054
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27448 22098 27476 23287
rect 27540 23254 27568 26182
rect 27908 25537 27936 26862
rect 28092 26382 28120 27814
rect 28276 26926 28304 28086
rect 28368 28082 28396 28562
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28736 27606 28764 28902
rect 29104 27996 29132 30058
rect 29196 29782 29224 30126
rect 29380 29850 29408 30194
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 29184 29776 29236 29782
rect 29184 29718 29236 29724
rect 29460 29504 29512 29510
rect 29460 29446 29512 29452
rect 29472 29034 29500 29446
rect 29368 29028 29420 29034
rect 29368 28970 29420 28976
rect 29460 29028 29512 29034
rect 29460 28970 29512 28976
rect 29380 28626 29408 28970
rect 29472 28762 29500 28970
rect 29460 28756 29512 28762
rect 29460 28698 29512 28704
rect 29368 28620 29420 28626
rect 29368 28562 29420 28568
rect 29184 28008 29236 28014
rect 29104 27968 29184 27996
rect 29184 27950 29236 27956
rect 28724 27600 28776 27606
rect 28724 27542 28776 27548
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 28264 26920 28316 26926
rect 28264 26862 28316 26868
rect 28276 26586 28304 26862
rect 28368 26858 28396 27406
rect 28736 27130 28764 27542
rect 29196 27402 29224 27950
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29288 27674 29316 27814
rect 29276 27668 29328 27674
rect 29276 27610 29328 27616
rect 29184 27396 29236 27402
rect 29184 27338 29236 27344
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 29104 27062 29132 27270
rect 29288 27062 29316 27610
rect 29092 27056 29144 27062
rect 29092 26998 29144 27004
rect 29276 27056 29328 27062
rect 29276 26998 29328 27004
rect 29104 26858 29132 26998
rect 28356 26852 28408 26858
rect 28356 26794 28408 26800
rect 29092 26852 29144 26858
rect 29092 26794 29144 26800
rect 28368 26586 28396 26794
rect 29104 26586 29132 26794
rect 28264 26580 28316 26586
rect 28264 26522 28316 26528
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 29092 26580 29144 26586
rect 29092 26522 29144 26528
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 28080 26376 28132 26382
rect 28080 26318 28132 26324
rect 28092 26042 28120 26318
rect 28080 26036 28132 26042
rect 28080 25978 28132 25984
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 27894 25528 27950 25537
rect 27894 25463 27950 25472
rect 27712 24268 27764 24274
rect 27712 24210 27764 24216
rect 27724 23594 27752 24210
rect 27712 23588 27764 23594
rect 27712 23530 27764 23536
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27252 22092 27304 22098
rect 27252 22034 27304 22040
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27448 21690 27476 22034
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27632 21146 27660 21422
rect 27724 21418 27752 22918
rect 28000 21962 28028 25774
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23730 28212 24142
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28184 23322 28212 23666
rect 28276 23662 28304 26522
rect 28908 26444 28960 26450
rect 28908 26386 28960 26392
rect 28920 25974 28948 26386
rect 29000 26240 29052 26246
rect 29000 26182 29052 26188
rect 29276 26240 29328 26246
rect 29276 26182 29328 26188
rect 28908 25968 28960 25974
rect 28722 25936 28778 25945
rect 28908 25910 28960 25916
rect 29012 25906 29040 26182
rect 28722 25871 28778 25880
rect 29000 25900 29052 25906
rect 28736 25838 28764 25871
rect 29000 25842 29052 25848
rect 28724 25832 28776 25838
rect 28724 25774 28776 25780
rect 28816 25764 28868 25770
rect 28816 25706 28868 25712
rect 28908 25764 28960 25770
rect 28908 25706 28960 25712
rect 28828 25294 28856 25706
rect 28920 25430 28948 25706
rect 28908 25424 28960 25430
rect 28908 25366 28960 25372
rect 28816 25288 28868 25294
rect 28816 25230 28868 25236
rect 28828 24410 28856 25230
rect 28920 24954 28948 25366
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28552 23866 28580 24346
rect 29288 24342 29316 26182
rect 29472 25770 29500 26522
rect 29564 26382 29592 34614
rect 29840 34542 29868 34682
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 29736 34128 29788 34134
rect 29656 34088 29736 34116
rect 29656 33590 29684 34088
rect 29736 34070 29788 34076
rect 29644 33584 29696 33590
rect 29644 33526 29696 33532
rect 29656 33114 29684 33526
rect 29736 33448 29788 33454
rect 29736 33390 29788 33396
rect 29748 33114 29776 33390
rect 30484 33386 30512 35702
rect 30748 35624 30800 35630
rect 30748 35566 30800 35572
rect 30760 35290 30788 35566
rect 30748 35284 30800 35290
rect 30748 35226 30800 35232
rect 30748 35148 30800 35154
rect 30748 35090 30800 35096
rect 30760 34746 30788 35090
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 29828 33380 29880 33386
rect 29828 33322 29880 33328
rect 30472 33380 30524 33386
rect 30472 33322 30524 33328
rect 29644 33108 29696 33114
rect 29644 33050 29696 33056
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 29840 32298 29868 33322
rect 30288 32972 30340 32978
rect 30288 32914 30340 32920
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 29828 32292 29880 32298
rect 29828 32234 29880 32240
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 29736 31680 29788 31686
rect 29736 31622 29788 31628
rect 29748 31278 29776 31622
rect 29736 31272 29788 31278
rect 29736 31214 29788 31220
rect 30024 30938 30052 31826
rect 30300 31686 30328 32914
rect 30576 32026 30604 32914
rect 30656 32224 30708 32230
rect 30656 32166 30708 32172
rect 30564 32020 30616 32026
rect 30564 31962 30616 31968
rect 30576 31890 30604 31962
rect 30564 31884 30616 31890
rect 30564 31826 30616 31832
rect 30288 31680 30340 31686
rect 30288 31622 30340 31628
rect 30196 31408 30248 31414
rect 30196 31350 30248 31356
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29736 30660 29788 30666
rect 29736 30602 29788 30608
rect 29656 29578 29684 30602
rect 29644 29572 29696 29578
rect 29644 29514 29696 29520
rect 29656 29170 29684 29514
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29748 28801 29776 30602
rect 30024 29306 30052 30874
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 29734 28792 29790 28801
rect 30024 28762 30052 29242
rect 29734 28727 29790 28736
rect 30012 28756 30064 28762
rect 30012 28698 30064 28704
rect 30104 28688 30156 28694
rect 30104 28630 30156 28636
rect 30116 28218 30144 28630
rect 30104 28212 30156 28218
rect 30104 28154 30156 28160
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 29460 25764 29512 25770
rect 29460 25706 29512 25712
rect 29748 25498 29776 25842
rect 29736 25492 29788 25498
rect 29736 25434 29788 25440
rect 29276 24336 29328 24342
rect 29276 24278 29328 24284
rect 29092 24064 29144 24070
rect 29092 24006 29144 24012
rect 29104 23866 29132 24006
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28276 22982 28304 23598
rect 28552 23474 28580 23802
rect 29104 23526 29132 23802
rect 29840 23730 29868 26930
rect 30012 26444 30064 26450
rect 30012 26386 30064 26392
rect 30024 25974 30052 26386
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 30208 25838 30236 31350
rect 30300 27849 30328 31622
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30484 29850 30512 31078
rect 30668 30734 30696 32166
rect 30748 31884 30800 31890
rect 30800 31844 30880 31872
rect 30748 31826 30800 31832
rect 30852 31142 30880 31844
rect 31036 31822 31064 36518
rect 31220 35154 31248 37420
rect 31300 37402 31352 37408
rect 31300 37120 31352 37126
rect 31300 37062 31352 37068
rect 31208 35148 31260 35154
rect 31208 35090 31260 35096
rect 31220 34610 31248 35090
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 31208 34400 31260 34406
rect 31208 34342 31260 34348
rect 31220 33998 31248 34342
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 31116 33856 31168 33862
rect 31116 33798 31168 33804
rect 31128 33522 31156 33798
rect 31312 33658 31340 37062
rect 31404 36106 31432 39510
rect 32048 39506 32076 43182
rect 32232 42906 32260 43250
rect 32220 42900 32272 42906
rect 32220 42842 32272 42848
rect 32232 42362 32260 42842
rect 32680 42696 32732 42702
rect 32680 42638 32732 42644
rect 32220 42356 32272 42362
rect 32220 42298 32272 42304
rect 32232 42158 32260 42298
rect 32692 42226 32720 42638
rect 32968 42634 32996 43823
rect 33048 43784 33100 43790
rect 33048 43726 33100 43732
rect 33060 43314 33088 43726
rect 33048 43308 33100 43314
rect 33048 43250 33100 43256
rect 33428 43110 33456 43930
rect 34704 43852 34756 43858
rect 34704 43794 34756 43800
rect 34244 43648 34296 43654
rect 34244 43590 34296 43596
rect 34256 43450 34284 43590
rect 34716 43450 34744 43794
rect 34244 43444 34296 43450
rect 34704 43444 34756 43450
rect 34244 43386 34296 43392
rect 34624 43404 34704 43432
rect 34256 43110 34284 43386
rect 33048 43104 33100 43110
rect 33048 43046 33100 43052
rect 33416 43104 33468 43110
rect 33416 43046 33468 43052
rect 34244 43104 34296 43110
rect 34244 43046 34296 43052
rect 33060 42906 33088 43046
rect 33048 42900 33100 42906
rect 33048 42842 33100 42848
rect 32956 42628 33008 42634
rect 32956 42570 33008 42576
rect 32680 42220 32732 42226
rect 32680 42162 32732 42168
rect 32220 42152 32272 42158
rect 32220 42094 32272 42100
rect 32232 40594 32260 42094
rect 33060 42022 33088 42842
rect 34624 42673 34652 43404
rect 34704 43386 34756 43392
rect 34808 43330 34836 44950
rect 35268 44810 35296 45290
rect 35256 44804 35308 44810
rect 35256 44746 35308 44752
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 35268 44266 35296 44746
rect 35348 44736 35400 44742
rect 35348 44678 35400 44684
rect 35360 44402 35388 44678
rect 35348 44396 35400 44402
rect 35348 44338 35400 44344
rect 35256 44260 35308 44266
rect 35256 44202 35308 44208
rect 35268 43926 35296 44202
rect 35360 43994 35388 44338
rect 35348 43988 35400 43994
rect 35348 43930 35400 43936
rect 35256 43920 35308 43926
rect 35256 43862 35308 43868
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34716 43302 34836 43330
rect 35348 43308 35400 43314
rect 34716 42702 34744 43302
rect 35348 43250 35400 43256
rect 34980 43172 35032 43178
rect 34980 43114 35032 43120
rect 34992 42838 35020 43114
rect 34796 42832 34848 42838
rect 34796 42774 34848 42780
rect 34980 42832 35032 42838
rect 34980 42774 35032 42780
rect 34704 42696 34756 42702
rect 34610 42664 34666 42673
rect 34704 42638 34756 42644
rect 34610 42599 34666 42608
rect 33508 42288 33560 42294
rect 33508 42230 33560 42236
rect 33048 42016 33100 42022
rect 33048 41958 33100 41964
rect 32312 41676 32364 41682
rect 32312 41618 32364 41624
rect 32324 41138 32352 41618
rect 32680 41472 32732 41478
rect 32680 41414 32732 41420
rect 32692 41138 32720 41414
rect 32312 41132 32364 41138
rect 32312 41074 32364 41080
rect 32680 41132 32732 41138
rect 32680 41074 32732 41080
rect 32324 41041 32352 41074
rect 32310 41032 32366 41041
rect 32310 40967 32366 40976
rect 32220 40588 32272 40594
rect 32220 40530 32272 40536
rect 32232 40186 32260 40530
rect 32220 40180 32272 40186
rect 32220 40122 32272 40128
rect 32220 39636 32272 39642
rect 32220 39578 32272 39584
rect 32036 39500 32088 39506
rect 32036 39442 32088 39448
rect 31852 39364 31904 39370
rect 31852 39306 31904 39312
rect 31484 38888 31536 38894
rect 31484 38830 31536 38836
rect 31496 38214 31524 38830
rect 31760 38752 31812 38758
rect 31760 38694 31812 38700
rect 31772 38486 31800 38694
rect 31864 38554 31892 39306
rect 32048 39098 32076 39442
rect 32036 39092 32088 39098
rect 32036 39034 32088 39040
rect 32128 38752 32180 38758
rect 32128 38694 32180 38700
rect 31852 38548 31904 38554
rect 31852 38490 31904 38496
rect 31760 38480 31812 38486
rect 31760 38422 31812 38428
rect 31576 38276 31628 38282
rect 31576 38218 31628 38224
rect 31484 38208 31536 38214
rect 31484 38150 31536 38156
rect 31496 37874 31524 38150
rect 31588 37874 31616 38218
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 31864 37806 31892 38490
rect 32140 38010 32168 38694
rect 32232 38418 32260 39578
rect 32324 39438 32352 40967
rect 32402 40624 32458 40633
rect 32402 40559 32458 40568
rect 32312 39432 32364 39438
rect 32312 39374 32364 39380
rect 32416 39284 32444 40559
rect 32692 40526 32720 41074
rect 33060 41002 33088 41958
rect 33048 40996 33100 41002
rect 33048 40938 33100 40944
rect 33324 40996 33376 41002
rect 33324 40938 33376 40944
rect 33336 40662 33364 40938
rect 33324 40656 33376 40662
rect 33324 40598 33376 40604
rect 32496 40520 32548 40526
rect 32496 40462 32548 40468
rect 32680 40520 32732 40526
rect 32680 40462 32732 40468
rect 32508 40118 32536 40462
rect 32864 40180 32916 40186
rect 32864 40122 32916 40128
rect 32496 40112 32548 40118
rect 32496 40054 32548 40060
rect 32324 39256 32444 39284
rect 32220 38412 32272 38418
rect 32220 38354 32272 38360
rect 32232 38010 32260 38354
rect 32128 38004 32180 38010
rect 32128 37946 32180 37952
rect 32220 38004 32272 38010
rect 32220 37946 32272 37952
rect 31852 37800 31904 37806
rect 31852 37742 31904 37748
rect 31760 36576 31812 36582
rect 31760 36518 31812 36524
rect 31392 36100 31444 36106
rect 31392 36042 31444 36048
rect 31772 34610 31800 36518
rect 32140 35766 32168 37946
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 32232 36922 32260 37198
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32324 36174 32352 39256
rect 32876 39098 32904 40122
rect 33232 39976 33284 39982
rect 33232 39918 33284 39924
rect 33244 39642 33272 39918
rect 33232 39636 33284 39642
rect 33232 39578 33284 39584
rect 33336 39574 33364 40598
rect 33416 39636 33468 39642
rect 33416 39578 33468 39584
rect 33324 39568 33376 39574
rect 33324 39510 33376 39516
rect 32864 39092 32916 39098
rect 32864 39034 32916 39040
rect 32876 38282 32904 39034
rect 33232 38888 33284 38894
rect 33232 38830 33284 38836
rect 33140 38820 33192 38826
rect 33140 38762 33192 38768
rect 33152 38654 33180 38762
rect 33060 38626 33180 38654
rect 33244 38654 33272 38830
rect 33336 38758 33364 39510
rect 33324 38752 33376 38758
rect 33324 38694 33376 38700
rect 33244 38626 33364 38654
rect 33060 38570 33088 38626
rect 33060 38542 33180 38570
rect 32864 38276 32916 38282
rect 32864 38218 32916 38224
rect 33152 38214 33180 38542
rect 33336 38486 33364 38626
rect 33324 38480 33376 38486
rect 33324 38422 33376 38428
rect 33428 38321 33456 39578
rect 33520 38350 33548 42230
rect 34060 42152 34112 42158
rect 34060 42094 34112 42100
rect 34150 42120 34206 42129
rect 33968 42016 34020 42022
rect 33968 41958 34020 41964
rect 33980 41750 34008 41958
rect 34072 41750 34100 42094
rect 34150 42055 34206 42064
rect 34164 42022 34192 42055
rect 34152 42016 34204 42022
rect 34152 41958 34204 41964
rect 33968 41744 34020 41750
rect 33968 41686 34020 41692
rect 34060 41744 34112 41750
rect 34060 41686 34112 41692
rect 33980 41274 34008 41686
rect 33968 41268 34020 41274
rect 33968 41210 34020 41216
rect 34072 41206 34100 41686
rect 34060 41200 34112 41206
rect 34060 41142 34112 41148
rect 34164 40769 34192 41958
rect 34716 41750 34744 42638
rect 34808 41818 34836 42774
rect 35360 42770 35388 43250
rect 35348 42764 35400 42770
rect 35348 42706 35400 42712
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 35636 42226 35664 45970
rect 36096 45966 36124 46582
rect 41524 46578 41552 46854
rect 41512 46572 41564 46578
rect 41512 46514 41564 46520
rect 36268 46504 36320 46510
rect 36268 46446 36320 46452
rect 36084 45960 36136 45966
rect 36084 45902 36136 45908
rect 36096 45286 36124 45902
rect 36280 45626 36308 46446
rect 41696 46436 41748 46442
rect 41696 46378 41748 46384
rect 42340 46436 42392 46442
rect 42340 46378 42392 46384
rect 36360 46368 36412 46374
rect 36360 46310 36412 46316
rect 36372 46170 36400 46310
rect 36360 46164 36412 46170
rect 36360 46106 36412 46112
rect 36268 45620 36320 45626
rect 36268 45562 36320 45568
rect 36280 45393 36308 45562
rect 36372 45490 36400 46106
rect 41604 46096 41656 46102
rect 41604 46038 41656 46044
rect 36544 46028 36596 46034
rect 36544 45970 36596 45976
rect 39856 46028 39908 46034
rect 39856 45970 39908 45976
rect 36452 45824 36504 45830
rect 36452 45766 36504 45772
rect 36360 45484 36412 45490
rect 36360 45426 36412 45432
rect 36266 45384 36322 45393
rect 36266 45319 36322 45328
rect 36464 45286 36492 45766
rect 36084 45280 36136 45286
rect 36084 45222 36136 45228
rect 36452 45280 36504 45286
rect 36452 45222 36504 45228
rect 36096 45082 36124 45222
rect 36084 45076 36136 45082
rect 36084 45018 36136 45024
rect 36464 45014 36492 45222
rect 36556 45014 36584 45970
rect 38108 45892 38160 45898
rect 38108 45834 38160 45840
rect 38120 45490 38148 45834
rect 39868 45626 39896 45970
rect 40592 45824 40644 45830
rect 40592 45766 40644 45772
rect 40684 45824 40736 45830
rect 40684 45766 40736 45772
rect 39856 45620 39908 45626
rect 39856 45562 39908 45568
rect 40604 45490 40632 45766
rect 36820 45484 36872 45490
rect 36820 45426 36872 45432
rect 38108 45484 38160 45490
rect 38108 45426 38160 45432
rect 38384 45484 38436 45490
rect 38384 45426 38436 45432
rect 40592 45484 40644 45490
rect 40592 45426 40644 45432
rect 36452 45008 36504 45014
rect 36452 44950 36504 44956
rect 36544 45008 36596 45014
rect 36544 44950 36596 44956
rect 36176 44872 36228 44878
rect 36176 44814 36228 44820
rect 35992 44396 36044 44402
rect 35992 44338 36044 44344
rect 35624 42220 35676 42226
rect 35544 42180 35624 42208
rect 34980 42084 35032 42090
rect 34980 42026 35032 42032
rect 34796 41812 34848 41818
rect 34796 41754 34848 41760
rect 34704 41744 34756 41750
rect 34704 41686 34756 41692
rect 34992 41546 35020 42026
rect 34980 41540 35032 41546
rect 34980 41482 35032 41488
rect 34612 41472 34664 41478
rect 34612 41414 34664 41420
rect 34796 41472 34848 41478
rect 34796 41414 34848 41420
rect 34624 41274 34652 41414
rect 34612 41268 34664 41274
rect 34612 41210 34664 41216
rect 34150 40760 34206 40769
rect 34808 40730 34836 41414
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 35164 40928 35216 40934
rect 35164 40870 35216 40876
rect 35176 40730 35204 40870
rect 34150 40695 34206 40704
rect 34796 40724 34848 40730
rect 34796 40666 34848 40672
rect 35164 40724 35216 40730
rect 35164 40666 35216 40672
rect 35256 40656 35308 40662
rect 35256 40598 35308 40604
rect 34244 40588 34296 40594
rect 34244 40530 34296 40536
rect 34256 40361 34284 40530
rect 34704 40520 34756 40526
rect 34704 40462 34756 40468
rect 34242 40352 34298 40361
rect 34242 40287 34298 40296
rect 34256 40186 34284 40287
rect 34244 40180 34296 40186
rect 34244 40122 34296 40128
rect 34716 40050 34744 40462
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 35268 40186 35296 40598
rect 35256 40180 35308 40186
rect 35256 40122 35308 40128
rect 35348 40180 35400 40186
rect 35348 40122 35400 40128
rect 34704 40044 34756 40050
rect 34704 39986 34756 39992
rect 34612 39500 34664 39506
rect 34612 39442 34664 39448
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 33704 38962 33732 39374
rect 34624 39098 34652 39442
rect 35360 39302 35388 40122
rect 35544 40050 35572 42180
rect 35624 42162 35676 42168
rect 35624 41744 35676 41750
rect 35624 41686 35676 41692
rect 35636 41206 35664 41686
rect 36004 41614 36032 44338
rect 36188 43994 36216 44814
rect 36464 44198 36492 44950
rect 36544 44260 36596 44266
rect 36544 44202 36596 44208
rect 36452 44192 36504 44198
rect 36452 44134 36504 44140
rect 36176 43988 36228 43994
rect 36176 43930 36228 43936
rect 36176 43852 36228 43858
rect 36176 43794 36228 43800
rect 36188 43450 36216 43794
rect 36176 43444 36228 43450
rect 36176 43386 36228 43392
rect 36084 42764 36136 42770
rect 36084 42706 36136 42712
rect 36176 42764 36228 42770
rect 36176 42706 36228 42712
rect 35992 41608 36044 41614
rect 35992 41550 36044 41556
rect 35624 41200 35676 41206
rect 35624 41142 35676 41148
rect 36004 41138 36032 41550
rect 36096 41138 36124 42706
rect 36188 42634 36216 42706
rect 36176 42628 36228 42634
rect 36176 42570 36228 42576
rect 36188 42362 36216 42570
rect 36176 42356 36228 42362
rect 36176 42298 36228 42304
rect 35992 41132 36044 41138
rect 35992 41074 36044 41080
rect 36084 41132 36136 41138
rect 36084 41074 36136 41080
rect 35900 40996 35952 41002
rect 35900 40938 35952 40944
rect 35912 40730 35940 40938
rect 36004 40730 36032 41074
rect 35900 40724 35952 40730
rect 35900 40666 35952 40672
rect 35992 40724 36044 40730
rect 35992 40666 36044 40672
rect 35532 40044 35584 40050
rect 35532 39986 35584 39992
rect 35544 39438 35572 39986
rect 35808 39976 35860 39982
rect 35808 39918 35860 39924
rect 35532 39432 35584 39438
rect 35532 39374 35584 39380
rect 35348 39296 35400 39302
rect 35348 39238 35400 39244
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34612 39092 34664 39098
rect 34612 39034 34664 39040
rect 33692 38956 33744 38962
rect 33692 38898 33744 38904
rect 35256 38888 35308 38894
rect 35256 38830 35308 38836
rect 33600 38752 33652 38758
rect 33600 38694 33652 38700
rect 33612 38418 33640 38694
rect 35268 38554 35296 38830
rect 35256 38548 35308 38554
rect 35256 38490 35308 38496
rect 33600 38412 33652 38418
rect 33600 38354 33652 38360
rect 33968 38412 34020 38418
rect 33968 38354 34020 38360
rect 35256 38412 35308 38418
rect 35256 38354 35308 38360
rect 33508 38344 33560 38350
rect 33414 38312 33470 38321
rect 33508 38286 33560 38292
rect 33414 38247 33470 38256
rect 33048 38208 33100 38214
rect 33048 38150 33100 38156
rect 33140 38208 33192 38214
rect 33140 38150 33192 38156
rect 33060 37738 33088 38150
rect 32680 37732 32732 37738
rect 32680 37674 32732 37680
rect 33048 37732 33100 37738
rect 33048 37674 33100 37680
rect 32692 37194 32720 37674
rect 33060 37466 33088 37674
rect 33048 37460 33100 37466
rect 33048 37402 33100 37408
rect 32680 37188 32732 37194
rect 32680 37130 32732 37136
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 32128 35760 32180 35766
rect 32128 35702 32180 35708
rect 32324 35494 32352 36110
rect 32128 35488 32180 35494
rect 32128 35430 32180 35436
rect 32312 35488 32364 35494
rect 32312 35430 32364 35436
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 31300 33652 31352 33658
rect 31300 33594 31352 33600
rect 31116 33516 31168 33522
rect 31116 33458 31168 33464
rect 31312 33134 31340 33594
rect 31392 33448 31444 33454
rect 31392 33390 31444 33396
rect 31128 33106 31340 33134
rect 31128 32842 31156 33106
rect 31116 32836 31168 32842
rect 31116 32778 31168 32784
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 30840 31136 30892 31142
rect 30840 31078 30892 31084
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30484 28014 30512 28494
rect 30852 28014 30880 31078
rect 31036 30394 31064 31758
rect 31404 30938 31432 33390
rect 31496 32201 31524 34478
rect 31760 33380 31812 33386
rect 31760 33322 31812 33328
rect 31668 32360 31720 32366
rect 31668 32302 31720 32308
rect 31482 32192 31538 32201
rect 31482 32127 31538 32136
rect 31392 30932 31444 30938
rect 31392 30874 31444 30880
rect 31116 30796 31168 30802
rect 31116 30738 31168 30744
rect 31024 30388 31076 30394
rect 31024 30330 31076 30336
rect 31128 30190 31156 30738
rect 31116 30184 31168 30190
rect 31116 30126 31168 30132
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 31036 29034 31064 29650
rect 31024 29028 31076 29034
rect 31024 28970 31076 28976
rect 31404 28626 31432 29990
rect 31496 29850 31524 32127
rect 31576 31204 31628 31210
rect 31680 31192 31708 32302
rect 31772 32026 31800 33322
rect 32140 33134 32168 35430
rect 32416 35290 32444 37062
rect 32692 36786 32720 37130
rect 32680 36780 32732 36786
rect 32680 36722 32732 36728
rect 32496 36644 32548 36650
rect 32496 36586 32548 36592
rect 32508 36378 32536 36586
rect 32496 36372 32548 36378
rect 32496 36314 32548 36320
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 32508 35834 32536 36314
rect 32864 36032 32916 36038
rect 32864 35974 32916 35980
rect 32496 35828 32548 35834
rect 32496 35770 32548 35776
rect 32876 35630 32904 35974
rect 32864 35624 32916 35630
rect 32864 35566 32916 35572
rect 32404 35284 32456 35290
rect 32404 35226 32456 35232
rect 32220 35148 32272 35154
rect 32220 35090 32272 35096
rect 32232 34066 32260 35090
rect 32416 34542 32444 35226
rect 32404 34536 32456 34542
rect 32404 34478 32456 34484
rect 32416 34202 32444 34478
rect 32404 34196 32456 34202
rect 32404 34138 32456 34144
rect 32876 34134 32904 35566
rect 32956 35080 33008 35086
rect 32956 35022 33008 35028
rect 32968 34610 32996 35022
rect 32956 34604 33008 34610
rect 32956 34546 33008 34552
rect 32864 34128 32916 34134
rect 32864 34070 32916 34076
rect 32220 34060 32272 34066
rect 32220 34002 32272 34008
rect 32232 33454 32260 34002
rect 32956 33924 33008 33930
rect 32956 33866 33008 33872
rect 32404 33856 32456 33862
rect 32404 33798 32456 33804
rect 32416 33658 32444 33798
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 32220 33448 32272 33454
rect 32220 33390 32272 33396
rect 32048 33106 32168 33134
rect 31852 32836 31904 32842
rect 31852 32778 31904 32784
rect 31864 32609 31892 32778
rect 31944 32768 31996 32774
rect 31944 32710 31996 32716
rect 31850 32600 31906 32609
rect 31850 32535 31906 32544
rect 31864 32502 31892 32535
rect 31852 32496 31904 32502
rect 31852 32438 31904 32444
rect 31760 32020 31812 32026
rect 31760 31962 31812 31968
rect 31864 31278 31892 32438
rect 31956 32366 31984 32710
rect 31944 32360 31996 32366
rect 31944 32302 31996 32308
rect 31956 31754 31984 32302
rect 32048 31890 32076 33106
rect 32324 32978 32352 33458
rect 32312 32972 32364 32978
rect 32312 32914 32364 32920
rect 32416 32774 32444 33594
rect 32968 33046 32996 33866
rect 32956 33040 33008 33046
rect 32586 33008 32642 33017
rect 32956 32982 33008 32988
rect 32586 32943 32642 32952
rect 32600 32910 32628 32943
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 32128 32496 32180 32502
rect 32416 32484 32444 32710
rect 32180 32456 32444 32484
rect 32128 32438 32180 32444
rect 32416 32230 32444 32456
rect 32404 32224 32456 32230
rect 32404 32166 32456 32172
rect 32128 31952 32180 31958
rect 32128 31894 32180 31900
rect 32312 31952 32364 31958
rect 32312 31894 32364 31900
rect 32036 31884 32088 31890
rect 32036 31826 32088 31832
rect 31944 31748 31996 31754
rect 31944 31690 31996 31696
rect 32036 31748 32088 31754
rect 32036 31690 32088 31696
rect 31956 31346 31984 31690
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 31628 31164 31708 31192
rect 31576 31146 31628 31152
rect 31680 30938 31708 31164
rect 31668 30932 31720 30938
rect 31668 30874 31720 30880
rect 31760 30932 31812 30938
rect 31760 30874 31812 30880
rect 31680 30122 31708 30874
rect 31772 30734 31800 30874
rect 31864 30802 31892 31214
rect 31852 30796 31904 30802
rect 31852 30738 31904 30744
rect 31956 30734 31984 31282
rect 31760 30728 31812 30734
rect 31944 30728 31996 30734
rect 31812 30676 31892 30682
rect 31760 30670 31892 30676
rect 31944 30670 31996 30676
rect 31772 30654 31892 30670
rect 31864 30258 31892 30654
rect 31944 30320 31996 30326
rect 31944 30262 31996 30268
rect 31852 30252 31904 30258
rect 31852 30194 31904 30200
rect 31668 30116 31720 30122
rect 31668 30058 31720 30064
rect 31680 29850 31708 30058
rect 31484 29844 31536 29850
rect 31484 29786 31536 29792
rect 31668 29844 31720 29850
rect 31668 29786 31720 29792
rect 31864 29782 31892 30194
rect 31852 29776 31904 29782
rect 31852 29718 31904 29724
rect 31668 29096 31720 29102
rect 31864 29073 31892 29718
rect 31668 29038 31720 29044
rect 31850 29064 31906 29073
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 31024 28620 31076 28626
rect 31024 28562 31076 28568
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31036 28218 31064 28562
rect 31024 28212 31076 28218
rect 31024 28154 31076 28160
rect 31496 28082 31524 28902
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30840 28008 30892 28014
rect 30840 27950 30892 27956
rect 30932 27940 30984 27946
rect 30932 27882 30984 27888
rect 30564 27872 30616 27878
rect 30286 27840 30342 27849
rect 30564 27814 30616 27820
rect 30286 27775 30342 27784
rect 30576 27606 30604 27814
rect 30564 27600 30616 27606
rect 30564 27542 30616 27548
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 30484 26586 30512 27406
rect 30576 27130 30604 27542
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30196 25832 30248 25838
rect 30196 25774 30248 25780
rect 30012 25764 30064 25770
rect 30012 25706 30064 25712
rect 30024 24886 30052 25706
rect 30576 25430 30604 27066
rect 30944 26994 30972 27882
rect 31496 27674 31524 28018
rect 31484 27668 31536 27674
rect 31484 27610 31536 27616
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 31036 27062 31064 27338
rect 31116 27328 31168 27334
rect 31116 27270 31168 27276
rect 31024 27056 31076 27062
rect 31024 26998 31076 27004
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 30944 26586 30972 26930
rect 31128 26858 31156 27270
rect 31588 27062 31616 28970
rect 31680 28558 31708 29038
rect 31850 28999 31906 29008
rect 31760 28960 31812 28966
rect 31760 28902 31812 28908
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 31680 27674 31708 28494
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31576 27056 31628 27062
rect 31576 26998 31628 27004
rect 31116 26852 31168 26858
rect 31116 26794 31168 26800
rect 30932 26580 30984 26586
rect 30932 26522 30984 26528
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30944 25702 30972 26386
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30564 25424 30616 25430
rect 30616 25384 30696 25412
rect 30564 25366 30616 25372
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30012 24880 30064 24886
rect 30012 24822 30064 24828
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 29368 23588 29420 23594
rect 29368 23530 29420 23536
rect 29092 23520 29144 23526
rect 28552 23446 28672 23474
rect 29092 23462 29144 23468
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28264 22976 28316 22982
rect 28552 22953 28580 23054
rect 28264 22918 28316 22924
rect 28538 22944 28594 22953
rect 28538 22879 28594 22888
rect 28552 22438 28580 22879
rect 28540 22432 28592 22438
rect 28540 22374 28592 22380
rect 28356 22024 28408 22030
rect 28552 22001 28580 22374
rect 28644 22166 28672 23446
rect 29380 22982 29408 23530
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29656 23254 29684 23462
rect 29552 23248 29604 23254
rect 29552 23190 29604 23196
rect 29644 23248 29696 23254
rect 29644 23190 29696 23196
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29196 22642 29224 22918
rect 29380 22778 29408 22918
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 28632 22160 28684 22166
rect 28632 22102 28684 22108
rect 28356 21966 28408 21972
rect 28538 21992 28594 22001
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 27712 21412 27764 21418
rect 27712 21354 27764 21360
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 25872 21004 25924 21010
rect 25872 20946 25924 20952
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 25884 20602 25912 20946
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 26528 20398 26556 20742
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19446 25452 19654
rect 25412 19440 25464 19446
rect 25412 19382 25464 19388
rect 25608 18426 25636 19790
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25700 19514 25728 19722
rect 26068 19514 26096 20266
rect 26528 20058 26556 20334
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26896 19854 26924 20402
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27264 19990 27292 20266
rect 27252 19984 27304 19990
rect 27252 19926 27304 19932
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26068 19174 26096 19450
rect 26896 19446 26924 19790
rect 27264 19514 27292 19926
rect 27632 19904 27660 21082
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27724 20398 27752 20810
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27724 20058 27752 20334
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27632 19876 27752 19904
rect 27724 19786 27752 19876
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27712 19780 27764 19786
rect 27712 19722 27764 19728
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26884 19440 26936 19446
rect 26884 19382 26936 19388
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26252 18630 26280 19178
rect 26700 18896 26752 18902
rect 26700 18838 26752 18844
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25608 18086 25636 18362
rect 26252 18154 26280 18566
rect 25780 18148 25832 18154
rect 25780 18090 25832 18096
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25516 16998 25544 17682
rect 25792 17542 25820 18090
rect 26620 17882 26648 18702
rect 26712 18426 26740 18838
rect 27632 18766 27660 19722
rect 28000 19417 28028 21898
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28184 21010 28212 21422
rect 28368 21418 28396 21966
rect 28538 21927 28594 21936
rect 28644 21690 28672 22102
rect 29564 22098 29592 23190
rect 29656 22506 29684 23190
rect 29644 22500 29696 22506
rect 29644 22442 29696 22448
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 28356 21412 28408 21418
rect 28356 21354 28408 21360
rect 28368 21146 28396 21354
rect 28356 21140 28408 21146
rect 28356 21082 28408 21088
rect 29288 21078 29316 21422
rect 29276 21072 29328 21078
rect 29276 21014 29328 21020
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28092 20534 28120 20946
rect 28184 20602 28212 20946
rect 29840 20942 29868 23666
rect 30024 23118 30052 24822
rect 30392 24818 30420 25230
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30104 24676 30156 24682
rect 30104 24618 30156 24624
rect 30116 23866 30144 24618
rect 30194 24440 30250 24449
rect 30194 24375 30250 24384
rect 30208 24274 30236 24375
rect 30196 24268 30248 24274
rect 30196 24210 30248 24216
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 30208 23730 30236 24210
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30024 21894 30052 23054
rect 30392 22710 30420 24754
rect 30576 24410 30604 25230
rect 30668 25158 30696 25384
rect 30838 25256 30894 25265
rect 30838 25191 30894 25200
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30668 24954 30696 25094
rect 30656 24948 30708 24954
rect 30656 24890 30708 24896
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30380 22704 30432 22710
rect 30380 22646 30432 22652
rect 30392 22012 30420 22646
rect 30748 22500 30800 22506
rect 30748 22442 30800 22448
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 30472 22024 30524 22030
rect 30392 21984 30472 22012
rect 30472 21966 30524 21972
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 30484 21622 30512 21966
rect 30576 21690 30604 22102
rect 30760 21865 30788 22442
rect 30746 21856 30802 21865
rect 30746 21791 30802 21800
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30748 21684 30800 21690
rect 30748 21626 30800 21632
rect 30472 21616 30524 21622
rect 30472 21558 30524 21564
rect 30760 21418 30788 21626
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30208 21078 30236 21286
rect 30196 21072 30248 21078
rect 30196 21014 30248 21020
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28080 20528 28132 20534
rect 28080 20470 28132 20476
rect 29000 20324 29052 20330
rect 29000 20266 29052 20272
rect 29012 19990 29040 20266
rect 29840 20058 29868 20878
rect 30208 20602 30236 21014
rect 30760 20602 30788 21354
rect 30196 20596 30248 20602
rect 30196 20538 30248 20544
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30116 20262 30144 20402
rect 30760 20330 30788 20538
rect 30196 20324 30248 20330
rect 30196 20266 30248 20272
rect 30748 20324 30800 20330
rect 30748 20266 30800 20272
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29828 20052 29880 20058
rect 29828 19994 29880 20000
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 27986 19408 28042 19417
rect 27986 19343 28042 19352
rect 27804 19236 27856 19242
rect 27804 19178 27856 19184
rect 27816 18902 27844 19178
rect 29012 18970 29040 19926
rect 29276 19916 29328 19922
rect 29276 19858 29328 19864
rect 29288 19310 29316 19858
rect 30116 19310 30144 20198
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 29288 18834 29316 19246
rect 29828 18896 29880 18902
rect 29828 18838 29880 18844
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 29276 18828 29328 18834
rect 29276 18770 29328 18776
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 26608 17876 26660 17882
rect 26528 17836 26608 17864
rect 25688 17536 25740 17542
rect 25688 17478 25740 17484
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25516 15094 25544 16934
rect 25700 16114 25728 17478
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25792 13938 25820 17478
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25976 16998 26004 17206
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25884 15638 25912 16934
rect 25976 16250 26004 16934
rect 26160 16250 26188 17002
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26528 16130 26556 17836
rect 26608 17818 26660 17824
rect 26712 17814 26740 18362
rect 27632 18290 27660 18702
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 27344 18148 27396 18154
rect 27344 18090 27396 18096
rect 26804 17814 26832 18090
rect 27356 17882 27384 18090
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 26700 17808 26752 17814
rect 26700 17750 26752 17756
rect 26792 17808 26844 17814
rect 26792 17750 26844 17756
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26620 17202 26648 17614
rect 26712 17338 26740 17750
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26620 16794 26648 17138
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 26792 16992 26844 16998
rect 27264 16946 27292 17002
rect 26844 16940 27292 16946
rect 26792 16934 27292 16940
rect 26804 16918 27292 16934
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26804 16726 26832 16918
rect 26792 16720 26844 16726
rect 26792 16662 26844 16668
rect 26884 16720 26936 16726
rect 26884 16662 26936 16668
rect 26528 16102 26740 16130
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25884 15162 25912 15574
rect 26160 15162 26188 15914
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26160 14890 26188 15098
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26436 14414 26464 15642
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25792 13462 25820 13874
rect 25780 13456 25832 13462
rect 25780 13398 25832 13404
rect 26528 12850 26556 14894
rect 26712 14550 26740 16102
rect 26804 14550 26832 16662
rect 26896 16250 26924 16662
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 27080 16114 27108 16526
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27080 15502 27108 16050
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 26700 14544 26752 14550
rect 26700 14486 26752 14492
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26712 13326 26740 14486
rect 26804 14074 26832 14486
rect 27356 14414 27384 17818
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27724 16998 27752 17206
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27724 16794 27752 16934
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27908 16522 27936 18566
rect 28368 18086 28396 18770
rect 29288 18426 29316 18770
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 28356 18080 28408 18086
rect 28356 18022 28408 18028
rect 28368 17882 28396 18022
rect 28356 17876 28408 17882
rect 28356 17818 28408 17824
rect 29196 17814 29224 18294
rect 29184 17808 29236 17814
rect 29184 17750 29236 17756
rect 28264 17740 28316 17746
rect 28264 17682 28316 17688
rect 27896 16516 27948 16522
rect 27896 16458 27948 16464
rect 28276 16454 28304 17682
rect 29196 17202 29224 17750
rect 29288 17746 29316 18362
rect 29564 18222 29592 18566
rect 29840 18290 29868 18838
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29276 17740 29328 17746
rect 29276 17682 29328 17688
rect 29288 17338 29316 17682
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28276 15162 28304 16390
rect 28368 15910 28396 16526
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28368 15706 28396 15846
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 28644 15638 28672 15846
rect 28632 15632 28684 15638
rect 28632 15574 28684 15580
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28736 15094 28764 15438
rect 28724 15088 28776 15094
rect 28724 15030 28776 15036
rect 28264 14952 28316 14958
rect 28264 14894 28316 14900
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27344 14408 27396 14414
rect 27344 14350 27396 14356
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26804 13462 26832 14010
rect 26988 13546 27016 14350
rect 27356 13938 27384 14350
rect 28276 14278 28304 14894
rect 28540 14816 28592 14822
rect 28592 14776 28672 14804
rect 28540 14758 28592 14764
rect 28264 14272 28316 14278
rect 28264 14214 28316 14220
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27080 13802 27108 13874
rect 27068 13796 27120 13802
rect 27068 13738 27120 13744
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 26988 13518 27108 13546
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 25688 12776 25740 12782
rect 26344 12753 26372 12786
rect 25688 12718 25740 12724
rect 26330 12744 26386 12753
rect 25332 12158 25452 12186
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11626 25360 12038
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 25332 10810 25360 11562
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25424 6866 25452 12158
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25516 10130 25544 10950
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25700 9722 25728 12718
rect 26056 12708 26108 12714
rect 26330 12679 26386 12688
rect 26056 12650 26108 12656
rect 26068 12442 26096 12650
rect 26620 12442 26648 13262
rect 26804 12986 26832 13398
rect 27080 13190 27108 13518
rect 27816 13258 27844 13670
rect 28276 13394 28304 14214
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28552 13462 28580 13670
rect 28540 13456 28592 13462
rect 28540 13398 28592 13404
rect 28264 13388 28316 13394
rect 28264 13330 28316 13336
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 27080 12918 27108 13126
rect 27068 12912 27120 12918
rect 27068 12854 27120 12860
rect 28092 12782 28120 13126
rect 28368 12850 28396 13262
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26792 12368 26844 12374
rect 26792 12310 26844 12316
rect 27804 12368 27856 12374
rect 27804 12310 27856 12316
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26252 11898 26280 12242
rect 26804 11898 26832 12310
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26792 11892 26844 11898
rect 26844 11852 27016 11880
rect 26792 11834 26844 11840
rect 26988 11626 27016 11852
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 26976 11620 27028 11626
rect 26976 11562 27028 11568
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 26712 11286 26740 11494
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26712 10810 26740 11222
rect 26804 11014 26832 11494
rect 27632 11286 27660 11630
rect 27816 11286 27844 12310
rect 27908 11665 27936 12718
rect 28368 12442 28396 12786
rect 28552 12646 28580 13398
rect 28644 12850 28672 14776
rect 29012 14770 29040 16934
rect 29092 16720 29144 16726
rect 29092 16662 29144 16668
rect 29104 15910 29132 16662
rect 29092 15904 29144 15910
rect 29092 15846 29144 15852
rect 29104 15094 29132 15846
rect 29380 15570 29408 18022
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 29472 16114 29500 17478
rect 29736 17264 29788 17270
rect 29736 17206 29788 17212
rect 29748 16114 29776 17206
rect 30116 17202 30144 17478
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30116 16114 30144 17138
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 29472 15706 29500 16050
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29184 15496 29236 15502
rect 29184 15438 29236 15444
rect 29092 15088 29144 15094
rect 29092 15030 29144 15036
rect 29012 14742 29132 14770
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28736 13802 28764 14418
rect 28724 13796 28776 13802
rect 28776 13756 28856 13784
rect 28724 13738 28776 13744
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28356 12436 28408 12442
rect 28356 12378 28408 12384
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28184 11898 28212 12174
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 27894 11656 27950 11665
rect 27894 11591 27950 11600
rect 28460 11558 28488 12242
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26804 10266 26832 10950
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 27080 10198 27108 10474
rect 27068 10192 27120 10198
rect 27068 10134 27120 10140
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 9178 25728 9454
rect 26252 9178 26280 10066
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 25700 8566 25728 9114
rect 26528 8974 26556 9386
rect 27080 9382 27108 10134
rect 27448 9926 27476 11086
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27540 10606 27568 10950
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27080 9110 27108 9318
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26528 8634 26556 8910
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 26700 8356 26752 8362
rect 26700 8298 26752 8304
rect 26068 7750 26096 8298
rect 26608 8016 26660 8022
rect 26712 8004 26740 8298
rect 27080 8294 27108 9046
rect 27448 8634 27476 9862
rect 27540 9382 27568 10542
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 28000 9178 28028 9454
rect 28184 9178 28212 10066
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 26660 7976 26740 8004
rect 26608 7958 26660 7964
rect 26712 7886 26740 7976
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 26068 7546 26096 7686
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25332 6322 25360 6598
rect 25424 6458 25452 6802
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 25332 5234 25360 5510
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 25424 4690 25452 6394
rect 25608 4690 25636 6598
rect 25976 4826 26004 7142
rect 26436 6186 26464 7142
rect 26712 7002 26740 7822
rect 26804 7206 26832 7958
rect 27632 7342 27660 8774
rect 28368 8430 28396 10406
rect 28460 10266 28488 11494
rect 28552 10538 28580 12582
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28644 10577 28672 11154
rect 28630 10568 28686 10577
rect 28540 10532 28592 10538
rect 28630 10503 28686 10512
rect 28540 10474 28592 10480
rect 28644 10470 28672 10503
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28644 9092 28672 10406
rect 28736 10130 28764 11290
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28644 9064 28764 9092
rect 28448 8560 28500 8566
rect 28448 8502 28500 8508
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 8090 28396 8366
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 28184 7546 28212 7958
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 26792 7200 26844 7206
rect 26792 7142 26844 7148
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 28184 6934 28212 7482
rect 28276 7274 28304 7822
rect 28264 7268 28316 7274
rect 28264 7210 28316 7216
rect 28172 6928 28224 6934
rect 28172 6870 28224 6876
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 27252 6724 27304 6730
rect 27252 6666 27304 6672
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27172 6322 27200 6598
rect 27264 6322 27292 6666
rect 28000 6390 28028 6734
rect 28184 6458 28212 6870
rect 28460 6458 28488 8502
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 26424 6180 26476 6186
rect 26424 6122 26476 6128
rect 27068 5840 27120 5846
rect 27068 5782 27120 5788
rect 26332 5636 26384 5642
rect 26332 5578 26384 5584
rect 26344 5370 26372 5578
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26896 5234 26924 5510
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25424 4282 25452 4626
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 26148 4208 26200 4214
rect 26148 4150 26200 4156
rect 26160 4010 26188 4150
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 26148 4004 26200 4010
rect 26148 3946 26200 3952
rect 26068 3398 26096 3946
rect 26436 3670 26464 4082
rect 26896 4010 26924 5170
rect 27080 5098 27108 5782
rect 27068 5092 27120 5098
rect 27068 5034 27120 5040
rect 27080 4826 27108 5034
rect 27068 4820 27120 4826
rect 27068 4762 27120 4768
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26988 4282 27016 4626
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 27172 4010 27200 6258
rect 27264 5681 27292 6258
rect 27356 5710 27384 6326
rect 28000 5914 28028 6326
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 28184 5846 28212 6394
rect 28460 6254 28488 6394
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28172 5840 28224 5846
rect 28172 5782 28224 5788
rect 28540 5840 28592 5846
rect 28540 5782 28592 5788
rect 27344 5704 27396 5710
rect 27250 5672 27306 5681
rect 27344 5646 27396 5652
rect 27250 5607 27306 5616
rect 28184 5370 28212 5782
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28460 5098 28488 5646
rect 28552 5370 28580 5782
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 28448 5092 28500 5098
rect 28448 5034 28500 5040
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 27160 4004 27212 4010
rect 27160 3946 27212 3952
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 26436 3194 26464 3606
rect 26896 3534 26924 3946
rect 28092 3942 28120 4558
rect 28276 4060 28304 4762
rect 28448 4752 28500 4758
rect 28448 4694 28500 4700
rect 28460 4146 28488 4694
rect 28552 4154 28580 5306
rect 28644 4282 28672 6598
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28448 4140 28500 4146
rect 28552 4126 28672 4154
rect 28448 4082 28500 4088
rect 28356 4072 28408 4078
rect 28276 4032 28356 4060
rect 28356 4014 28408 4020
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 26620 3194 26648 3470
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25884 2514 25912 2790
rect 26620 2650 26648 3130
rect 27632 2990 27660 3334
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 28184 2650 28212 3334
rect 28460 3126 28488 3878
rect 28644 3670 28672 4126
rect 28632 3664 28684 3670
rect 28632 3606 28684 3612
rect 28448 3120 28500 3126
rect 28448 3062 28500 3068
rect 28264 2984 28316 2990
rect 28264 2926 28316 2932
rect 28276 2650 28304 2926
rect 28356 2916 28408 2922
rect 28356 2858 28408 2864
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 28264 2644 28316 2650
rect 28264 2586 28316 2592
rect 28368 2514 28396 2858
rect 28644 2854 28672 3606
rect 28736 2922 28764 9064
rect 28828 9042 28856 13756
rect 29104 12714 29132 14742
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 28908 12640 28960 12646
rect 28908 12582 28960 12588
rect 28920 12374 28948 12582
rect 28908 12368 28960 12374
rect 28908 12310 28960 12316
rect 28920 11694 28948 12310
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 29104 11898 29132 12174
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 29000 10804 29052 10810
rect 29000 10746 29052 10752
rect 29012 9518 29040 10746
rect 29196 9722 29224 15438
rect 29380 15026 29408 15506
rect 29460 15088 29512 15094
rect 29460 15030 29512 15036
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29276 14952 29328 14958
rect 29276 14894 29328 14900
rect 29288 14550 29316 14894
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 29380 14482 29408 14962
rect 29472 14890 29500 15030
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29368 14476 29420 14482
rect 29368 14418 29420 14424
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29288 13190 29316 13942
rect 29380 13870 29408 14418
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29380 13530 29408 13806
rect 29472 13734 29500 14826
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 30104 13456 30156 13462
rect 30104 13398 30156 13404
rect 29276 13184 29328 13190
rect 29276 13126 29328 13132
rect 29288 11218 29316 13126
rect 30012 12912 30064 12918
rect 30012 12854 30064 12860
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29380 12442 29408 12786
rect 30024 12714 30052 12854
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 29368 12436 29420 12442
rect 29368 12378 29420 12384
rect 30024 11762 30052 12650
rect 30116 12646 30144 13398
rect 30104 12640 30156 12646
rect 30104 12582 30156 12588
rect 30012 11756 30064 11762
rect 30012 11698 30064 11704
rect 30116 11626 30144 12582
rect 29828 11620 29880 11626
rect 29828 11562 29880 11568
rect 30104 11620 30156 11626
rect 30104 11562 30156 11568
rect 29840 11354 29868 11562
rect 30116 11354 30144 11562
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 29276 11212 29328 11218
rect 29276 11154 29328 11160
rect 29288 10810 29316 11154
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29276 10804 29328 10810
rect 29276 10746 29328 10752
rect 30024 10266 30052 11086
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30012 10260 30064 10266
rect 30012 10202 30064 10208
rect 30024 10062 30052 10202
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 30116 9926 30144 10406
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29184 9716 29236 9722
rect 29184 9658 29236 9664
rect 29196 9518 29224 9658
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29288 9500 29316 9862
rect 30208 9518 30236 20266
rect 30852 19922 30880 25191
rect 30944 23474 30972 25638
rect 31128 24954 31156 26794
rect 31668 25696 31720 25702
rect 31668 25638 31720 25644
rect 31680 25498 31708 25638
rect 31668 25492 31720 25498
rect 31668 25434 31720 25440
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 31668 24812 31720 24818
rect 31668 24754 31720 24760
rect 31680 24410 31708 24754
rect 31668 24404 31720 24410
rect 31668 24346 31720 24352
rect 31300 24268 31352 24274
rect 31300 24210 31352 24216
rect 31312 23866 31340 24210
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31312 23474 31340 23802
rect 30944 23446 31064 23474
rect 31312 23446 31432 23474
rect 31036 22817 31064 23446
rect 31206 23216 31262 23225
rect 31206 23151 31262 23160
rect 31022 22808 31078 22817
rect 31022 22743 31078 22752
rect 31220 21622 31248 23151
rect 31404 22409 31432 23446
rect 31390 22400 31446 22409
rect 31390 22335 31446 22344
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31680 21554 31708 21830
rect 31668 21548 31720 21554
rect 31772 21536 31800 28902
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31864 27946 31892 28154
rect 31852 27940 31904 27946
rect 31852 27882 31904 27888
rect 31852 26036 31904 26042
rect 31852 25978 31904 25984
rect 31864 23662 31892 25978
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 31852 23248 31904 23254
rect 31852 23190 31904 23196
rect 31864 22778 31892 23190
rect 31852 22772 31904 22778
rect 31852 22714 31904 22720
rect 31772 21508 31892 21536
rect 31668 21490 31720 21496
rect 31760 21412 31812 21418
rect 31760 21354 31812 21360
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30944 19922 30972 20810
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 31036 20466 31064 20742
rect 31772 20602 31800 21354
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31024 20460 31076 20466
rect 31024 20402 31076 20408
rect 30840 19916 30892 19922
rect 30840 19858 30892 19864
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 30852 19514 30880 19858
rect 30944 19514 30972 19858
rect 31036 19854 31064 20402
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 31116 19780 31168 19786
rect 31116 19722 31168 19728
rect 31128 19514 31156 19722
rect 30840 19508 30892 19514
rect 30840 19450 30892 19456
rect 30932 19508 30984 19514
rect 30932 19450 30984 19456
rect 31116 19508 31168 19514
rect 31116 19450 31168 19456
rect 30748 19304 30800 19310
rect 30748 19246 30800 19252
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 30576 17814 30604 18838
rect 30760 18834 30788 19246
rect 31484 19168 31536 19174
rect 31298 19136 31354 19145
rect 31484 19110 31536 19116
rect 31298 19071 31354 19080
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30760 18426 30788 18770
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30852 18222 30880 18702
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30852 17746 30880 18158
rect 31116 18148 31168 18154
rect 31116 18090 31168 18096
rect 31208 18148 31260 18154
rect 31208 18090 31260 18096
rect 30656 17740 30708 17746
rect 30656 17682 30708 17688
rect 30840 17740 30892 17746
rect 30840 17682 30892 17688
rect 30668 17338 30696 17682
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30852 17066 30880 17682
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30840 17060 30892 17066
rect 30840 17002 30892 17008
rect 30380 16448 30432 16454
rect 30944 16425 30972 17478
rect 31128 16658 31156 18090
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 30380 16390 30432 16396
rect 30930 16416 30986 16425
rect 30392 16250 30420 16390
rect 30930 16351 30986 16360
rect 31128 16250 31156 16594
rect 31220 16561 31248 18090
rect 31312 17338 31340 19071
rect 31496 18698 31524 19110
rect 31864 18834 31892 21508
rect 31956 20040 31984 30262
rect 32048 28694 32076 31690
rect 32140 30870 32168 31894
rect 32324 31822 32352 31894
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32404 31816 32456 31822
rect 32508 31804 32536 32846
rect 32968 32502 32996 32982
rect 33152 32570 33180 36314
rect 33324 35556 33376 35562
rect 33324 35498 33376 35504
rect 33336 35290 33364 35498
rect 33324 35284 33376 35290
rect 33324 35226 33376 35232
rect 33336 34678 33364 35226
rect 33520 34746 33548 38286
rect 33980 38010 34008 38354
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 33968 38004 34020 38010
rect 33968 37946 34020 37952
rect 35268 37670 35296 38354
rect 35256 37664 35308 37670
rect 35256 37606 35308 37612
rect 33784 37392 33836 37398
rect 33784 37334 33836 37340
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33612 36650 33640 37198
rect 33600 36644 33652 36650
rect 33600 36586 33652 36592
rect 33796 36582 33824 37334
rect 35360 37330 35388 39238
rect 35532 38752 35584 38758
rect 35820 38729 35848 39918
rect 36096 39370 36124 41074
rect 36084 39364 36136 39370
rect 36084 39306 36136 39312
rect 36096 39030 36124 39306
rect 36084 39024 36136 39030
rect 36084 38966 36136 38972
rect 35532 38694 35584 38700
rect 35806 38720 35862 38729
rect 35440 38412 35492 38418
rect 35440 38354 35492 38360
rect 35452 38010 35480 38354
rect 35544 38010 35572 38694
rect 35806 38655 35862 38664
rect 35440 38004 35492 38010
rect 35440 37946 35492 37952
rect 35532 38004 35584 38010
rect 35532 37946 35584 37952
rect 35452 37330 35480 37946
rect 35544 37738 35572 37946
rect 35532 37732 35584 37738
rect 35532 37674 35584 37680
rect 35348 37324 35400 37330
rect 35348 37266 35400 37272
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 34336 37256 34388 37262
rect 34336 37198 34388 37204
rect 34152 36848 34204 36854
rect 34152 36790 34204 36796
rect 33784 36576 33836 36582
rect 33784 36518 33836 36524
rect 33692 36168 33744 36174
rect 33692 36110 33744 36116
rect 33704 35834 33732 36110
rect 33692 35828 33744 35834
rect 33692 35770 33744 35776
rect 33796 35737 33824 36518
rect 34060 36304 34112 36310
rect 34060 36246 34112 36252
rect 34072 35766 34100 36246
rect 34060 35760 34112 35766
rect 33782 35728 33838 35737
rect 34060 35702 34112 35708
rect 33782 35663 33838 35672
rect 33796 35630 33824 35663
rect 33784 35624 33836 35630
rect 33784 35566 33836 35572
rect 34072 35290 34100 35702
rect 34060 35284 34112 35290
rect 34060 35226 34112 35232
rect 34164 35154 34192 36790
rect 34348 36310 34376 37198
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35360 36854 35388 37266
rect 35452 36922 35480 37266
rect 35440 36916 35492 36922
rect 35440 36858 35492 36864
rect 35348 36848 35400 36854
rect 35348 36790 35400 36796
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 34336 36304 34388 36310
rect 34336 36246 34388 36252
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34152 35148 34204 35154
rect 34152 35090 34204 35096
rect 34796 35148 34848 35154
rect 34796 35090 34848 35096
rect 33416 34740 33468 34746
rect 33416 34682 33468 34688
rect 33508 34740 33560 34746
rect 33508 34682 33560 34688
rect 33324 34672 33376 34678
rect 33324 34614 33376 34620
rect 33428 34513 33456 34682
rect 33414 34504 33470 34513
rect 34808 34474 34836 35090
rect 35348 34944 35400 34950
rect 35348 34886 35400 34892
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 33414 34439 33470 34448
rect 34796 34468 34848 34474
rect 34796 34410 34848 34416
rect 35164 34468 35216 34474
rect 35164 34410 35216 34416
rect 34612 34060 34664 34066
rect 34612 34002 34664 34008
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33692 32836 33744 32842
rect 33692 32778 33744 32784
rect 33600 32768 33652 32774
rect 33600 32710 33652 32716
rect 33140 32564 33192 32570
rect 33140 32506 33192 32512
rect 32956 32496 33008 32502
rect 32956 32438 33008 32444
rect 33612 32366 33640 32710
rect 33600 32360 33652 32366
rect 33600 32302 33652 32308
rect 32456 31776 32536 31804
rect 32404 31758 32456 31764
rect 32220 31136 32272 31142
rect 32220 31078 32272 31084
rect 32128 30864 32180 30870
rect 32128 30806 32180 30812
rect 32140 29850 32168 30806
rect 32232 30297 32260 31078
rect 32416 30938 32444 31758
rect 33612 31754 33640 32302
rect 33704 31958 33732 32778
rect 33784 32768 33836 32774
rect 33784 32710 33836 32716
rect 33796 32026 33824 32710
rect 33888 32434 33916 33934
rect 34152 33856 34204 33862
rect 34152 33798 34204 33804
rect 33968 33380 34020 33386
rect 33968 33322 34020 33328
rect 33980 32842 34008 33322
rect 33968 32836 34020 32842
rect 33968 32778 34020 32784
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 33692 31952 33744 31958
rect 33692 31894 33744 31900
rect 33600 31748 33652 31754
rect 33600 31690 33652 31696
rect 34060 31748 34112 31754
rect 34060 31690 34112 31696
rect 32496 31680 32548 31686
rect 32548 31640 32628 31668
rect 32496 31622 32548 31628
rect 32600 31414 32628 31640
rect 32588 31408 32640 31414
rect 32588 31350 32640 31356
rect 32600 31142 32628 31350
rect 32588 31136 32640 31142
rect 32588 31078 32640 31084
rect 32404 30932 32456 30938
rect 32404 30874 32456 30880
rect 32496 30592 32548 30598
rect 32600 30580 32628 31078
rect 34072 30938 34100 31690
rect 34164 31278 34192 33798
rect 34336 33448 34388 33454
rect 34624 33425 34652 34002
rect 35176 33998 35204 34410
rect 35256 34400 35308 34406
rect 35256 34342 35308 34348
rect 35164 33992 35216 33998
rect 35164 33934 35216 33940
rect 35268 33930 35296 34342
rect 35360 34134 35388 34886
rect 35348 34128 35400 34134
rect 35348 34070 35400 34076
rect 34704 33924 34756 33930
rect 34704 33866 34756 33872
rect 35256 33924 35308 33930
rect 35256 33866 35308 33872
rect 34336 33390 34388 33396
rect 34610 33416 34666 33425
rect 34244 32972 34296 32978
rect 34244 32914 34296 32920
rect 34256 32570 34284 32914
rect 34244 32564 34296 32570
rect 34244 32506 34296 32512
rect 34348 31482 34376 33390
rect 34716 33386 34744 33866
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35268 33658 35296 33866
rect 35544 33658 35572 36518
rect 35624 35216 35676 35222
rect 35622 35184 35624 35193
rect 35676 35184 35678 35193
rect 35622 35119 35678 35128
rect 35636 34542 35664 35119
rect 35820 35018 35848 38655
rect 35992 38208 36044 38214
rect 35992 38150 36044 38156
rect 36004 37874 36032 38150
rect 36464 38010 36492 44134
rect 36556 43858 36584 44202
rect 36544 43852 36596 43858
rect 36544 43794 36596 43800
rect 36636 43648 36688 43654
rect 36636 43590 36688 43596
rect 36648 43178 36676 43590
rect 36832 43314 36860 45426
rect 38396 45082 38424 45426
rect 39580 45280 39632 45286
rect 39580 45222 39632 45228
rect 38384 45076 38436 45082
rect 38384 45018 38436 45024
rect 37740 44940 37792 44946
rect 37792 44900 37872 44928
rect 37740 44882 37792 44888
rect 37844 44402 37872 44900
rect 39304 44872 39356 44878
rect 39304 44814 39356 44820
rect 38568 44736 38620 44742
rect 38568 44678 38620 44684
rect 37832 44396 37884 44402
rect 37832 44338 37884 44344
rect 37844 44305 37872 44338
rect 38580 44334 38608 44678
rect 38568 44328 38620 44334
rect 37830 44296 37886 44305
rect 38568 44270 38620 44276
rect 37830 44231 37886 44240
rect 37832 44192 37884 44198
rect 37832 44134 37884 44140
rect 37464 43376 37516 43382
rect 37464 43318 37516 43324
rect 36820 43308 36872 43314
rect 36820 43250 36872 43256
rect 36544 43172 36596 43178
rect 36544 43114 36596 43120
rect 36636 43172 36688 43178
rect 36636 43114 36688 43120
rect 36556 42906 36584 43114
rect 36544 42900 36596 42906
rect 36544 42842 36596 42848
rect 36544 42560 36596 42566
rect 36544 42502 36596 42508
rect 36556 42226 36584 42502
rect 36544 42220 36596 42226
rect 36544 42162 36596 42168
rect 36648 42090 36676 43114
rect 36728 42832 36780 42838
rect 36832 42820 36860 43250
rect 36780 42792 36860 42820
rect 36728 42774 36780 42780
rect 36820 42696 36872 42702
rect 36820 42638 36872 42644
rect 36832 42226 36860 42638
rect 36820 42220 36872 42226
rect 36820 42162 36872 42168
rect 36636 42084 36688 42090
rect 36636 42026 36688 42032
rect 36648 41818 36676 42026
rect 36636 41812 36688 41818
rect 36636 41754 36688 41760
rect 36648 41002 36676 41754
rect 37372 41472 37424 41478
rect 37372 41414 37424 41420
rect 37384 41138 37412 41414
rect 37372 41132 37424 41138
rect 37372 41074 37424 41080
rect 36636 40996 36688 41002
rect 36636 40938 36688 40944
rect 37188 40996 37240 41002
rect 37188 40938 37240 40944
rect 36544 40588 36596 40594
rect 36544 40530 36596 40536
rect 36556 40118 36584 40530
rect 36544 40112 36596 40118
rect 36544 40054 36596 40060
rect 36648 39914 36676 40938
rect 37200 40662 37228 40938
rect 37384 40730 37412 41074
rect 37372 40724 37424 40730
rect 37372 40666 37424 40672
rect 37188 40656 37240 40662
rect 37188 40598 37240 40604
rect 36912 40044 36964 40050
rect 36912 39986 36964 39992
rect 36636 39908 36688 39914
rect 36636 39850 36688 39856
rect 36648 39642 36676 39850
rect 36820 39840 36872 39846
rect 36820 39782 36872 39788
rect 36832 39642 36860 39782
rect 36636 39636 36688 39642
rect 36636 39578 36688 39584
rect 36820 39636 36872 39642
rect 36820 39578 36872 39584
rect 36648 39098 36676 39578
rect 36924 39098 36952 39986
rect 36636 39092 36688 39098
rect 36636 39034 36688 39040
rect 36912 39092 36964 39098
rect 36912 39034 36964 39040
rect 37372 38752 37424 38758
rect 37372 38694 37424 38700
rect 36912 38412 36964 38418
rect 36912 38354 36964 38360
rect 36452 38004 36504 38010
rect 36452 37946 36504 37952
rect 35992 37868 36044 37874
rect 35992 37810 36044 37816
rect 36004 37398 36032 37810
rect 36636 37732 36688 37738
rect 36636 37674 36688 37680
rect 36544 37664 36596 37670
rect 36544 37606 36596 37612
rect 35992 37392 36044 37398
rect 35992 37334 36044 37340
rect 36268 37324 36320 37330
rect 36268 37266 36320 37272
rect 36280 36582 36308 37266
rect 36268 36576 36320 36582
rect 36268 36518 36320 36524
rect 36084 35148 36136 35154
rect 36084 35090 36136 35096
rect 35808 35012 35860 35018
rect 35808 34954 35860 34960
rect 36096 34746 36124 35090
rect 36176 35080 36228 35086
rect 36176 35022 36228 35028
rect 36084 34740 36136 34746
rect 36084 34682 36136 34688
rect 35624 34536 35676 34542
rect 35624 34478 35676 34484
rect 35636 34202 35664 34478
rect 35624 34196 35676 34202
rect 35624 34138 35676 34144
rect 35808 33992 35860 33998
rect 35808 33934 35860 33940
rect 35624 33856 35676 33862
rect 35624 33798 35676 33804
rect 35256 33652 35308 33658
rect 35532 33652 35584 33658
rect 35308 33612 35480 33640
rect 35256 33594 35308 33600
rect 34610 33351 34612 33360
rect 34664 33351 34666 33360
rect 34704 33380 34756 33386
rect 34612 33322 34664 33328
rect 34704 33322 34756 33328
rect 35256 33380 35308 33386
rect 35256 33322 35308 33328
rect 34624 32502 34652 33322
rect 35268 32978 35296 33322
rect 35346 33144 35402 33153
rect 35452 33114 35480 33612
rect 35532 33594 35584 33600
rect 35636 33590 35664 33798
rect 35624 33584 35676 33590
rect 35624 33526 35676 33532
rect 35820 33522 35848 33934
rect 35808 33516 35860 33522
rect 35808 33458 35860 33464
rect 35820 33134 35848 33458
rect 35346 33079 35402 33088
rect 35440 33108 35492 33114
rect 35256 32972 35308 32978
rect 35256 32914 35308 32920
rect 34704 32768 34756 32774
rect 34704 32710 34756 32716
rect 34716 32570 34744 32710
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34794 32600 34850 32609
rect 34704 32564 34756 32570
rect 34940 32592 35236 32612
rect 34794 32535 34850 32544
rect 34704 32506 34756 32512
rect 34612 32496 34664 32502
rect 34612 32438 34664 32444
rect 34336 31476 34388 31482
rect 34336 31418 34388 31424
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 33232 30728 33284 30734
rect 33284 30688 33364 30716
rect 33232 30670 33284 30676
rect 33140 30660 33192 30666
rect 33140 30602 33192 30608
rect 32548 30552 32628 30580
rect 32496 30534 32548 30540
rect 32600 30394 32628 30552
rect 32588 30388 32640 30394
rect 32588 30330 32640 30336
rect 32218 30288 32274 30297
rect 32218 30223 32274 30232
rect 32496 30184 32548 30190
rect 32496 30126 32548 30132
rect 32128 29844 32180 29850
rect 32128 29786 32180 29792
rect 32220 28756 32272 28762
rect 32220 28698 32272 28704
rect 32036 28688 32088 28694
rect 32036 28630 32088 28636
rect 32036 27940 32088 27946
rect 32036 27882 32088 27888
rect 32048 26450 32076 27882
rect 32232 27538 32260 28698
rect 32508 28626 32536 30126
rect 32600 30054 32628 30330
rect 32956 30116 33008 30122
rect 32956 30058 33008 30064
rect 32588 30048 32640 30054
rect 32588 29990 32640 29996
rect 32600 29306 32628 29990
rect 32588 29300 32640 29306
rect 32588 29242 32640 29248
rect 32968 29034 32996 30058
rect 33048 29572 33100 29578
rect 33048 29514 33100 29520
rect 32956 29028 33008 29034
rect 32956 28970 33008 28976
rect 32862 28656 32918 28665
rect 32496 28620 32548 28626
rect 32496 28562 32548 28568
rect 32680 28620 32732 28626
rect 32862 28591 32918 28600
rect 32680 28562 32732 28568
rect 32404 28212 32456 28218
rect 32404 28154 32456 28160
rect 32416 27656 32444 28154
rect 32508 27878 32536 28562
rect 32692 28218 32720 28562
rect 32680 28212 32732 28218
rect 32680 28154 32732 28160
rect 32496 27872 32548 27878
rect 32496 27814 32548 27820
rect 32496 27668 32548 27674
rect 32416 27628 32496 27656
rect 32496 27610 32548 27616
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32232 26586 32260 27474
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 32220 26580 32272 26586
rect 32220 26522 32272 26528
rect 32036 26444 32088 26450
rect 32036 26386 32088 26392
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32140 26042 32168 26386
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32036 25832 32088 25838
rect 32036 25774 32088 25780
rect 32048 23361 32076 25774
rect 32128 25696 32180 25702
rect 32128 25638 32180 25644
rect 32140 24818 32168 25638
rect 32312 25424 32364 25430
rect 32312 25366 32364 25372
rect 32324 25158 32352 25366
rect 32312 25152 32364 25158
rect 32312 25094 32364 25100
rect 32324 24954 32352 25094
rect 32312 24948 32364 24954
rect 32312 24890 32364 24896
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32312 24676 32364 24682
rect 32312 24618 32364 24624
rect 32324 24342 32352 24618
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32312 24336 32364 24342
rect 32312 24278 32364 24284
rect 32232 23866 32260 24278
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 32324 23730 32352 24278
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32034 23352 32090 23361
rect 32034 23287 32090 23296
rect 32220 23112 32272 23118
rect 32220 23054 32272 23060
rect 32232 22778 32260 23054
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32140 21146 32168 21966
rect 32312 21412 32364 21418
rect 32312 21354 32364 21360
rect 32128 21140 32180 21146
rect 32128 21082 32180 21088
rect 32324 21078 32352 21354
rect 32312 21072 32364 21078
rect 32312 21014 32364 21020
rect 32324 20233 32352 21014
rect 32310 20224 32366 20233
rect 32310 20159 32366 20168
rect 32416 20058 32444 26998
rect 32508 26790 32536 27610
rect 32496 26784 32548 26790
rect 32496 26726 32548 26732
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32508 24886 32536 25230
rect 32692 24886 32720 25774
rect 32496 24880 32548 24886
rect 32496 24822 32548 24828
rect 32680 24880 32732 24886
rect 32680 24822 32732 24828
rect 32876 23633 32904 28591
rect 33060 28014 33088 29514
rect 33048 28008 33100 28014
rect 33048 27950 33100 27956
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32968 26926 32996 27814
rect 33060 27674 33088 27950
rect 33048 27668 33100 27674
rect 33048 27610 33100 27616
rect 32956 26920 33008 26926
rect 32956 26862 33008 26868
rect 32586 23624 32642 23633
rect 32586 23559 32642 23568
rect 32862 23624 32918 23633
rect 32862 23559 32918 23568
rect 32496 23248 32548 23254
rect 32496 23190 32548 23196
rect 32508 22642 32536 23190
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32496 22228 32548 22234
rect 32496 22170 32548 22176
rect 32508 21690 32536 22170
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32600 21146 32628 23559
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32692 22098 32720 22578
rect 32680 22092 32732 22098
rect 32680 22034 32732 22040
rect 32692 21418 32720 22034
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32600 20602 32628 21082
rect 32680 21004 32732 21010
rect 32680 20946 32732 20952
rect 32692 20602 32720 20946
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32680 20596 32732 20602
rect 32680 20538 32732 20544
rect 32404 20052 32456 20058
rect 31956 20012 32076 20040
rect 31944 19916 31996 19922
rect 31944 19858 31996 19864
rect 31956 19174 31984 19858
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31852 18828 31904 18834
rect 31852 18770 31904 18776
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 31864 18426 31892 18770
rect 31852 18420 31904 18426
rect 31852 18362 31904 18368
rect 31864 18290 31892 18362
rect 31852 18284 31904 18290
rect 31852 18226 31904 18232
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31496 17814 31524 18022
rect 31484 17808 31536 17814
rect 31484 17750 31536 17756
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 31300 17332 31352 17338
rect 31300 17274 31352 17280
rect 31588 17134 31616 17546
rect 31668 17264 31720 17270
rect 31668 17206 31720 17212
rect 31576 17128 31628 17134
rect 31576 17070 31628 17076
rect 31680 16590 31708 17206
rect 31668 16584 31720 16590
rect 31206 16552 31262 16561
rect 31668 16526 31720 16532
rect 31206 16487 31262 16496
rect 31220 16454 31248 16487
rect 31208 16448 31260 16454
rect 31208 16390 31260 16396
rect 31576 16448 31628 16454
rect 31576 16390 31628 16396
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30392 16046 30420 16186
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30300 13326 30328 14758
rect 30392 13462 30420 15846
rect 31588 15570 31616 16390
rect 31680 16250 31708 16526
rect 31668 16244 31720 16250
rect 31668 16186 31720 16192
rect 31680 15706 31708 16186
rect 31668 15700 31720 15706
rect 31668 15642 31720 15648
rect 31576 15564 31628 15570
rect 31576 15506 31628 15512
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30576 13938 30604 14554
rect 31496 14074 31524 14894
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31772 14074 31800 14418
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30576 13530 30604 13874
rect 31956 13870 31984 19110
rect 32048 18970 32076 20012
rect 32404 19994 32456 20000
rect 32692 19990 32720 20538
rect 32680 19984 32732 19990
rect 32680 19926 32732 19932
rect 32404 19304 32456 19310
rect 32404 19246 32456 19252
rect 32416 19174 32444 19246
rect 32404 19168 32456 19174
rect 32784 19145 32812 21558
rect 32968 20602 32996 26862
rect 33048 26376 33100 26382
rect 33048 26318 33100 26324
rect 33060 25838 33088 26318
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 33048 22432 33100 22438
rect 33048 22374 33100 22380
rect 33060 22234 33088 22374
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 32956 20596 33008 20602
rect 32956 20538 33008 20544
rect 33048 20528 33100 20534
rect 33048 20470 33100 20476
rect 32956 19848 33008 19854
rect 32956 19790 33008 19796
rect 32404 19110 32456 19116
rect 32770 19136 32826 19145
rect 32416 18970 32444 19110
rect 32770 19071 32826 19080
rect 32036 18964 32088 18970
rect 32036 18906 32088 18912
rect 32404 18964 32456 18970
rect 32404 18906 32456 18912
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32232 17338 32260 17682
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 32036 17128 32088 17134
rect 32036 17070 32088 17076
rect 32048 16454 32076 17070
rect 32232 16658 32260 17274
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32036 16448 32088 16454
rect 32036 16390 32088 16396
rect 32128 16040 32180 16046
rect 32232 16028 32260 16594
rect 32180 16000 32260 16028
rect 32128 15982 32180 15988
rect 32232 15910 32260 16000
rect 32036 15904 32088 15910
rect 32036 15846 32088 15852
rect 32220 15904 32272 15910
rect 32220 15846 32272 15852
rect 32048 15638 32076 15846
rect 32232 15706 32260 15846
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32036 15632 32088 15638
rect 32036 15574 32088 15580
rect 32048 15162 32076 15574
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 32034 15056 32090 15065
rect 32034 14991 32090 15000
rect 31944 13864 31996 13870
rect 31944 13806 31996 13812
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30668 12986 30696 13262
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30392 12238 30420 12582
rect 30760 12374 30788 13194
rect 31300 12640 31352 12646
rect 31300 12582 31352 12588
rect 30748 12368 30800 12374
rect 30748 12310 30800 12316
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30484 10742 30512 11154
rect 30472 10736 30524 10742
rect 30472 10678 30524 10684
rect 30484 10606 30512 10678
rect 30380 10600 30432 10606
rect 30380 10542 30432 10548
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30392 10266 30420 10542
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30392 9722 30420 10066
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30668 9722 30696 9998
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30656 9716 30708 9722
rect 30656 9658 30708 9664
rect 29368 9512 29420 9518
rect 29288 9472 29368 9500
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 28828 8634 28856 8978
rect 28816 8628 28868 8634
rect 28816 8570 28868 8576
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 29012 6934 29040 8366
rect 29196 6934 29224 9454
rect 29288 9042 29316 9472
rect 29368 9454 29420 9460
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30392 9450 30420 9658
rect 30012 9444 30064 9450
rect 30012 9386 30064 9392
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29276 9036 29328 9042
rect 29276 8978 29328 8984
rect 29288 8566 29316 8978
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29276 8560 29328 8566
rect 29276 8502 29328 8508
rect 29564 8498 29592 8910
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29656 7954 29684 9318
rect 29644 7948 29696 7954
rect 29644 7890 29696 7896
rect 29656 7002 29684 7890
rect 29644 6996 29696 7002
rect 29644 6938 29696 6944
rect 29000 6928 29052 6934
rect 29000 6870 29052 6876
rect 29184 6928 29236 6934
rect 29184 6870 29236 6876
rect 28816 6724 28868 6730
rect 28816 6666 28868 6672
rect 28828 6390 28856 6666
rect 29012 6458 29040 6870
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28816 6384 28868 6390
rect 28816 6326 28868 6332
rect 29012 4282 29040 6394
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29644 5636 29696 5642
rect 29644 5578 29696 5584
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 29472 4826 29500 5510
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29656 4622 29684 5578
rect 29840 5166 29868 6054
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 29840 4826 29868 5102
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29644 4616 29696 4622
rect 29644 4558 29696 4564
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 29472 4010 29500 4218
rect 29656 4146 29684 4558
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29368 4004 29420 4010
rect 29368 3946 29420 3952
rect 29460 4004 29512 4010
rect 29460 3946 29512 3952
rect 29380 3602 29408 3946
rect 30024 3670 30052 9386
rect 30852 9178 30880 11494
rect 30932 11144 30984 11150
rect 30932 11086 30984 11092
rect 30944 10674 30972 11086
rect 31312 10810 31340 12582
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31588 11354 31616 11562
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31300 10804 31352 10810
rect 31300 10746 31352 10752
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30840 9036 30892 9042
rect 30840 8978 30892 8984
rect 30852 8634 30880 8978
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 31576 8560 31628 8566
rect 31576 8502 31628 8508
rect 31392 8492 31444 8498
rect 31312 8452 31392 8480
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30300 8022 30328 8298
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 30288 8016 30340 8022
rect 30288 7958 30340 7964
rect 30300 7478 30328 7958
rect 30484 7546 30512 8230
rect 31312 7750 31340 8452
rect 31392 8434 31444 8440
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30288 7472 30340 7478
rect 30288 7414 30340 7420
rect 30104 6928 30156 6934
rect 30104 6870 30156 6876
rect 30116 6118 30144 6870
rect 30300 6458 30328 7414
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6934 30604 7142
rect 30564 6928 30616 6934
rect 30564 6870 30616 6876
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30300 6186 30328 6394
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30288 6180 30340 6186
rect 30288 6122 30340 6128
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30116 4758 30144 6054
rect 30300 5846 30328 6122
rect 30288 5840 30340 5846
rect 30288 5782 30340 5788
rect 30484 5778 30512 6258
rect 30564 6248 30616 6254
rect 30564 6190 30616 6196
rect 30576 5914 30604 6190
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 30484 5370 30512 5714
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30104 4752 30156 4758
rect 30104 4694 30156 4700
rect 30668 4690 30696 7686
rect 30852 7410 30880 7686
rect 30840 7404 30892 7410
rect 30840 7346 30892 7352
rect 30932 7268 30984 7274
rect 30932 7210 30984 7216
rect 30944 6934 30972 7210
rect 30932 6928 30984 6934
rect 30932 6870 30984 6876
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 30840 5772 30892 5778
rect 30840 5714 30892 5720
rect 30852 5166 30880 5714
rect 31036 5234 31064 5850
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 30840 5160 30892 5166
rect 30840 5102 30892 5108
rect 30656 4684 30708 4690
rect 30656 4626 30708 4632
rect 30852 4622 30880 5102
rect 31024 5092 31076 5098
rect 31024 5034 31076 5040
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 30012 3664 30064 3670
rect 30012 3606 30064 3612
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 3194 29132 3334
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29104 2990 29132 3130
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 28724 2916 28776 2922
rect 28724 2858 28776 2864
rect 28632 2848 28684 2854
rect 28632 2790 28684 2796
rect 30024 2514 30052 3606
rect 30852 3602 30880 4558
rect 31036 4214 31064 5034
rect 31312 4826 31340 7686
rect 31496 7410 31524 8434
rect 31588 8362 31616 8502
rect 31576 8356 31628 8362
rect 31576 8298 31628 8304
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 31496 7206 31524 7346
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31772 6458 31800 6734
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31484 6112 31536 6118
rect 31484 6054 31536 6060
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31496 4690 31524 6054
rect 31772 4826 31800 6394
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31484 4684 31536 4690
rect 31484 4626 31536 4632
rect 31300 4276 31352 4282
rect 31300 4218 31352 4224
rect 31024 4208 31076 4214
rect 31024 4150 31076 4156
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30840 3596 30892 3602
rect 30840 3538 30892 3544
rect 30196 3188 30248 3194
rect 30196 3130 30248 3136
rect 30208 2514 30236 3130
rect 30300 2854 30328 3538
rect 30852 3194 30880 3538
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 30944 3058 30972 3470
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 30300 2310 30328 2790
rect 30944 2650 30972 2994
rect 31036 2922 31064 4150
rect 31312 4010 31340 4218
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31300 4004 31352 4010
rect 31300 3946 31352 3952
rect 31024 2916 31076 2922
rect 31024 2858 31076 2864
rect 31220 2650 31248 3946
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31208 2644 31260 2650
rect 31208 2586 31260 2592
rect 31956 2514 31984 4966
rect 32048 4154 32076 14991
rect 32324 10826 32352 18566
rect 32416 18222 32444 18906
rect 32968 18873 32996 19790
rect 33060 19334 33088 20470
rect 33152 20466 33180 30602
rect 33232 29844 33284 29850
rect 33232 29786 33284 29792
rect 33244 29510 33272 29786
rect 33336 29646 33364 30688
rect 33416 30592 33468 30598
rect 33416 30534 33468 30540
rect 33428 30190 33456 30534
rect 33784 30388 33836 30394
rect 33784 30330 33836 30336
rect 33416 30184 33468 30190
rect 33416 30126 33468 30132
rect 33692 29708 33744 29714
rect 33692 29650 33744 29656
rect 33324 29640 33376 29646
rect 33324 29582 33376 29588
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33336 28150 33364 29582
rect 33508 29232 33560 29238
rect 33508 29174 33560 29180
rect 33520 28762 33548 29174
rect 33704 29102 33732 29650
rect 33796 29170 33824 30330
rect 34072 30258 34100 30874
rect 34520 30796 34572 30802
rect 34520 30738 34572 30744
rect 34532 30258 34560 30738
rect 34624 30666 34652 32438
rect 34808 32366 34836 32535
rect 35360 32434 35388 33079
rect 35440 33050 35492 33056
rect 35728 33106 35848 33134
rect 35440 32972 35492 32978
rect 35492 32932 35572 32960
rect 35440 32914 35492 32920
rect 35440 32564 35492 32570
rect 35440 32506 35492 32512
rect 35348 32428 35400 32434
rect 35348 32370 35400 32376
rect 34796 32360 34848 32366
rect 34796 32302 34848 32308
rect 34888 32292 34940 32298
rect 34888 32234 34940 32240
rect 34900 32026 34928 32234
rect 34888 32020 34940 32026
rect 34808 31980 34888 32008
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34716 31482 34744 31758
rect 34808 31482 34836 31980
rect 34888 31962 34940 31968
rect 35070 31920 35126 31929
rect 35070 31855 35126 31864
rect 35084 31822 35112 31855
rect 35072 31816 35124 31822
rect 35072 31758 35124 31764
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35360 31482 35388 32370
rect 35452 32230 35480 32506
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 35452 31754 35480 32166
rect 35440 31748 35492 31754
rect 35440 31690 35492 31696
rect 35544 31686 35572 32932
rect 35728 32910 35756 33106
rect 36096 32978 36124 34682
rect 36084 32972 36136 32978
rect 36084 32914 36136 32920
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35728 32502 35756 32846
rect 35808 32836 35860 32842
rect 35808 32778 35860 32784
rect 35716 32496 35768 32502
rect 35716 32438 35768 32444
rect 35820 32026 35848 32778
rect 35900 32768 35952 32774
rect 35900 32710 35952 32716
rect 35808 32020 35860 32026
rect 35808 31962 35860 31968
rect 35912 31890 35940 32710
rect 35992 32360 36044 32366
rect 35992 32302 36044 32308
rect 36004 32026 36032 32302
rect 35992 32020 36044 32026
rect 35992 31962 36044 31968
rect 35900 31884 35952 31890
rect 35900 31826 35952 31832
rect 35532 31680 35584 31686
rect 35532 31622 35584 31628
rect 34704 31476 34756 31482
rect 34704 31418 34756 31424
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34716 31362 34744 31418
rect 34716 31334 34928 31362
rect 34704 31272 34756 31278
rect 34704 31214 34756 31220
rect 34716 31142 34744 31214
rect 34704 31136 34756 31142
rect 34704 31078 34756 31084
rect 34716 30938 34744 31078
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34612 30660 34664 30666
rect 34612 30602 34664 30608
rect 34624 30326 34652 30602
rect 34612 30320 34664 30326
rect 34612 30262 34664 30268
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 34520 30252 34572 30258
rect 34520 30194 34572 30200
rect 33968 29572 34020 29578
rect 33968 29514 34020 29520
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 33692 29096 33744 29102
rect 33692 29038 33744 29044
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 33704 28694 33732 29038
rect 33692 28688 33744 28694
rect 33692 28630 33744 28636
rect 33324 28144 33376 28150
rect 33324 28086 33376 28092
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 33612 26897 33640 26930
rect 33876 26920 33928 26926
rect 33598 26888 33654 26897
rect 33876 26862 33928 26868
rect 33598 26823 33654 26832
rect 33888 26586 33916 26862
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 33980 26450 34008 29514
rect 34072 28558 34100 30194
rect 34532 29850 34560 30194
rect 34520 29844 34572 29850
rect 34440 29804 34520 29832
rect 34336 29776 34388 29782
rect 34336 29718 34388 29724
rect 34348 29510 34376 29718
rect 34336 29504 34388 29510
rect 34336 29446 34388 29452
rect 34348 29034 34376 29446
rect 34336 29028 34388 29034
rect 34336 28970 34388 28976
rect 34244 28960 34296 28966
rect 34244 28902 34296 28908
rect 34256 28665 34284 28902
rect 34242 28656 34298 28665
rect 34242 28591 34298 28600
rect 34336 28620 34388 28626
rect 34440 28608 34468 29804
rect 34520 29786 34572 29792
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34532 29170 34560 29446
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 34532 28762 34560 28970
rect 34520 28756 34572 28762
rect 34520 28698 34572 28704
rect 34388 28580 34468 28608
rect 34336 28562 34388 28568
rect 34060 28552 34112 28558
rect 34060 28494 34112 28500
rect 34072 28218 34100 28494
rect 34060 28212 34112 28218
rect 34060 28154 34112 28160
rect 34440 27674 34468 28580
rect 34624 28490 34652 30262
rect 34716 30122 34744 30874
rect 34900 30734 34928 31334
rect 34888 30728 34940 30734
rect 34808 30688 34888 30716
rect 34808 30394 34836 30688
rect 34888 30670 34940 30676
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 34704 30116 34756 30122
rect 34704 30058 34756 30064
rect 34716 29714 34744 30058
rect 34704 29708 34756 29714
rect 34704 29650 34756 29656
rect 34716 29034 34744 29650
rect 35360 29646 35388 31418
rect 35544 30394 35572 31622
rect 35900 31204 35952 31210
rect 35900 31146 35952 31152
rect 35912 30938 35940 31146
rect 35900 30932 35952 30938
rect 35900 30874 35952 30880
rect 35624 30592 35676 30598
rect 35624 30534 35676 30540
rect 35532 30388 35584 30394
rect 35532 30330 35584 30336
rect 35636 30122 35664 30534
rect 35912 30394 35940 30874
rect 36188 30802 36216 35022
rect 36280 32570 36308 36518
rect 36556 36242 36584 37606
rect 36648 36922 36676 37674
rect 36924 37670 36952 38354
rect 36912 37664 36964 37670
rect 36912 37606 36964 37612
rect 36636 36916 36688 36922
rect 36636 36858 36688 36864
rect 36648 36650 36676 36858
rect 36636 36644 36688 36650
rect 36636 36586 36688 36592
rect 36544 36236 36596 36242
rect 36544 36178 36596 36184
rect 36556 35494 36584 36178
rect 36648 35834 36676 36586
rect 36728 36236 36780 36242
rect 36728 36178 36780 36184
rect 36636 35828 36688 35834
rect 36636 35770 36688 35776
rect 36648 35562 36676 35770
rect 36740 35630 36768 36178
rect 36728 35624 36780 35630
rect 36728 35566 36780 35572
rect 36636 35556 36688 35562
rect 36636 35498 36688 35504
rect 36544 35488 36596 35494
rect 36596 35436 36676 35442
rect 36544 35430 36676 35436
rect 36556 35414 36676 35430
rect 36452 34128 36504 34134
rect 36452 34070 36504 34076
rect 36360 33652 36412 33658
rect 36360 33594 36412 33600
rect 36372 32842 36400 33594
rect 36464 33386 36492 34070
rect 36452 33380 36504 33386
rect 36452 33322 36504 33328
rect 36464 33096 36492 33322
rect 36544 33108 36596 33114
rect 36464 33068 36544 33096
rect 36544 33050 36596 33056
rect 36360 32836 36412 32842
rect 36360 32778 36412 32784
rect 36268 32564 36320 32570
rect 36268 32506 36320 32512
rect 36556 32434 36584 33050
rect 36544 32428 36596 32434
rect 36544 32370 36596 32376
rect 36648 32366 36676 35414
rect 36740 35154 36768 35566
rect 36728 35148 36780 35154
rect 36728 35090 36780 35096
rect 36740 34406 36768 35090
rect 36818 34640 36874 34649
rect 36818 34575 36874 34584
rect 36728 34400 36780 34406
rect 36728 34342 36780 34348
rect 36740 34202 36768 34342
rect 36728 34196 36780 34202
rect 36728 34138 36780 34144
rect 36728 33924 36780 33930
rect 36728 33866 36780 33872
rect 36740 33658 36768 33866
rect 36728 33652 36780 33658
rect 36728 33594 36780 33600
rect 36832 33522 36860 34575
rect 36924 33658 36952 37606
rect 37096 37120 37148 37126
rect 37096 37062 37148 37068
rect 37108 36786 37136 37062
rect 37096 36780 37148 36786
rect 37096 36722 37148 36728
rect 37108 36310 37136 36722
rect 37096 36304 37148 36310
rect 37096 36246 37148 36252
rect 37096 36032 37148 36038
rect 37096 35974 37148 35980
rect 37108 35698 37136 35974
rect 37188 35760 37240 35766
rect 37188 35702 37240 35708
rect 37096 35692 37148 35698
rect 37096 35634 37148 35640
rect 37108 35222 37136 35634
rect 37096 35216 37148 35222
rect 37096 35158 37148 35164
rect 37200 34950 37228 35702
rect 37188 34944 37240 34950
rect 37188 34886 37240 34892
rect 37200 34542 37228 34886
rect 37004 34536 37056 34542
rect 37004 34478 37056 34484
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 36912 33652 36964 33658
rect 36912 33594 36964 33600
rect 36820 33516 36872 33522
rect 36820 33458 36872 33464
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 36912 32360 36964 32366
rect 36912 32302 36964 32308
rect 36268 32292 36320 32298
rect 36268 32234 36320 32240
rect 36280 32201 36308 32234
rect 36266 32192 36322 32201
rect 36266 32127 36322 32136
rect 36924 31958 36952 32302
rect 36912 31952 36964 31958
rect 36912 31894 36964 31900
rect 36268 31884 36320 31890
rect 36268 31826 36320 31832
rect 36280 31482 36308 31826
rect 36924 31754 36952 31894
rect 36912 31748 36964 31754
rect 36912 31690 36964 31696
rect 36268 31476 36320 31482
rect 36268 31418 36320 31424
rect 36924 30802 36952 31690
rect 36176 30796 36228 30802
rect 36176 30738 36228 30744
rect 36912 30796 36964 30802
rect 36912 30738 36964 30744
rect 35900 30388 35952 30394
rect 35900 30330 35952 30336
rect 35624 30116 35676 30122
rect 35624 30058 35676 30064
rect 35636 29850 35664 30058
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 35624 29844 35676 29850
rect 35624 29786 35676 29792
rect 35348 29640 35400 29646
rect 35348 29582 35400 29588
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 35256 29164 35308 29170
rect 35256 29106 35308 29112
rect 34704 29028 34756 29034
rect 34704 28970 34756 28976
rect 35268 28626 35296 29106
rect 35360 28762 35388 29582
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35256 28620 35308 28626
rect 35256 28562 35308 28568
rect 34612 28484 34664 28490
rect 34612 28426 34664 28432
rect 34624 28218 34652 28426
rect 34704 28416 34756 28422
rect 34704 28358 34756 28364
rect 34612 28212 34664 28218
rect 34612 28154 34664 28160
rect 34428 27668 34480 27674
rect 34428 27610 34480 27616
rect 34152 27532 34204 27538
rect 34152 27474 34204 27480
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34164 27062 34192 27474
rect 34152 27056 34204 27062
rect 34152 26998 34204 27004
rect 34348 26926 34376 27474
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34336 26920 34388 26926
rect 34336 26862 34388 26868
rect 34440 26450 34468 27406
rect 34520 26580 34572 26586
rect 34520 26522 34572 26528
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 34428 26444 34480 26450
rect 34428 26386 34480 26392
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 33244 24818 33272 26182
rect 33336 26042 33364 26386
rect 34152 26308 34204 26314
rect 34152 26250 34204 26256
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33692 25968 33744 25974
rect 33598 25936 33654 25945
rect 33692 25910 33744 25916
rect 33598 25871 33654 25880
rect 33324 24948 33376 24954
rect 33324 24890 33376 24896
rect 33232 24812 33284 24818
rect 33232 24754 33284 24760
rect 33244 24410 33272 24754
rect 33336 24682 33364 24890
rect 33508 24812 33560 24818
rect 33508 24754 33560 24760
rect 33324 24676 33376 24682
rect 33324 24618 33376 24624
rect 33232 24404 33284 24410
rect 33232 24346 33284 24352
rect 33520 24342 33548 24754
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 33336 23118 33364 23598
rect 33520 23322 33548 24278
rect 33612 23594 33640 25871
rect 33704 25401 33732 25910
rect 33874 25528 33930 25537
rect 33874 25463 33930 25472
rect 33690 25392 33746 25401
rect 33690 25327 33746 25336
rect 33600 23588 33652 23594
rect 33600 23530 33652 23536
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 33888 23186 33916 25463
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 34072 23322 34100 24006
rect 34060 23316 34112 23322
rect 34060 23258 34112 23264
rect 34164 23186 34192 26250
rect 34440 25498 34468 26386
rect 34532 25702 34560 26522
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34428 25492 34480 25498
rect 34428 25434 34480 25440
rect 34244 25356 34296 25362
rect 34244 25298 34296 25304
rect 34256 24682 34284 25298
rect 34244 24676 34296 24682
rect 34244 24618 34296 24624
rect 34256 24585 34284 24618
rect 34242 24576 34298 24585
rect 34242 24511 34298 24520
rect 34256 23798 34284 24511
rect 34532 24342 34560 25638
rect 34612 25424 34664 25430
rect 34612 25366 34664 25372
rect 34624 24954 34652 25366
rect 34612 24948 34664 24954
rect 34612 24890 34664 24896
rect 34520 24336 34572 24342
rect 34520 24278 34572 24284
rect 34244 23792 34296 23798
rect 34244 23734 34296 23740
rect 34532 23526 34560 24278
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 33876 23180 33928 23186
rect 33876 23122 33928 23128
rect 34152 23180 34204 23186
rect 34152 23122 34204 23128
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33888 22778 33916 23122
rect 33876 22772 33928 22778
rect 33796 22732 33876 22760
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 33336 20806 33364 21422
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 33336 20534 33364 20742
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 33060 19306 33180 19334
rect 33152 19174 33180 19306
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 32954 18864 33010 18873
rect 32772 18828 32824 18834
rect 32954 18799 33010 18808
rect 32772 18770 32824 18776
rect 32784 18222 32812 18770
rect 33244 18290 33272 20334
rect 33428 19174 33456 20334
rect 33796 20058 33824 22732
rect 33876 22714 33928 22720
rect 34164 22438 34192 23122
rect 34152 22432 34204 22438
rect 34152 22374 34204 22380
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 33888 21554 33916 21966
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 34164 21486 34192 22374
rect 34532 22166 34560 23462
rect 34520 22160 34572 22166
rect 34520 22102 34572 22108
rect 34532 21690 34560 22102
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 34152 21480 34204 21486
rect 34152 21422 34204 21428
rect 34532 21350 34560 21626
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34152 21004 34204 21010
rect 34152 20946 34204 20952
rect 34164 20262 34192 20946
rect 34532 20602 34560 21286
rect 34520 20596 34572 20602
rect 34520 20538 34572 20544
rect 34532 20330 34560 20538
rect 34520 20324 34572 20330
rect 34520 20266 34572 20272
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 33784 20052 33836 20058
rect 33784 19994 33836 20000
rect 33876 19984 33928 19990
rect 33876 19926 33928 19932
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33416 19168 33468 19174
rect 33416 19110 33468 19116
rect 33520 18834 33548 19450
rect 33888 19174 33916 19926
rect 33600 19168 33652 19174
rect 33600 19110 33652 19116
rect 33876 19168 33928 19174
rect 33876 19110 33928 19116
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 33232 18284 33284 18290
rect 33232 18226 33284 18232
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32416 17542 32444 18158
rect 32772 17808 32824 17814
rect 32772 17750 32824 17756
rect 32496 17604 32548 17610
rect 32496 17546 32548 17552
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32416 17134 32444 17478
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32416 16046 32444 17070
rect 32508 16998 32536 17546
rect 32784 16998 32812 17750
rect 32496 16992 32548 16998
rect 32496 16934 32548 16940
rect 32772 16992 32824 16998
rect 32772 16934 32824 16940
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 32416 15706 32444 15982
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32404 14816 32456 14822
rect 32404 14758 32456 14764
rect 32416 13870 32444 14758
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32404 13728 32456 13734
rect 32404 13670 32456 13676
rect 32416 12918 32444 13670
rect 32404 12912 32456 12918
rect 32404 12854 32456 12860
rect 32508 12374 32536 16934
rect 32784 15570 32812 16934
rect 32772 15564 32824 15570
rect 32772 15506 32824 15512
rect 32784 14958 32812 15506
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32876 14550 32904 18226
rect 33324 18148 33376 18154
rect 33324 18090 33376 18096
rect 33336 17882 33364 18090
rect 33612 18086 33640 19110
rect 33600 18080 33652 18086
rect 33600 18022 33652 18028
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33428 16590 33456 16934
rect 33508 16652 33560 16658
rect 33508 16594 33560 16600
rect 33416 16584 33468 16590
rect 33416 16526 33468 16532
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33140 15428 33192 15434
rect 33140 15370 33192 15376
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 32876 14074 32904 14486
rect 33152 14414 33180 15370
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33244 15026 33272 15302
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 32784 13394 32812 13806
rect 32876 13462 32904 14010
rect 32864 13456 32916 13462
rect 32864 13398 32916 13404
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 32588 13320 32640 13326
rect 32588 13262 32640 13268
rect 32600 12646 32628 13262
rect 32876 12918 32904 13398
rect 32864 12912 32916 12918
rect 32864 12854 32916 12860
rect 33336 12782 33364 16050
rect 33520 15978 33548 16594
rect 33508 15972 33560 15978
rect 33508 15914 33560 15920
rect 33520 15638 33548 15914
rect 33508 15632 33560 15638
rect 33508 15574 33560 15580
rect 33520 15094 33548 15574
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33428 13870 33456 14350
rect 33416 13864 33468 13870
rect 33416 13806 33468 13812
rect 33428 13530 33456 13806
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33520 13190 33548 14486
rect 33508 13184 33560 13190
rect 33508 13126 33560 13132
rect 33520 12782 33548 13126
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 32956 12708 33008 12714
rect 32956 12650 33008 12656
rect 32588 12640 32640 12646
rect 32588 12582 32640 12588
rect 32496 12368 32548 12374
rect 32496 12310 32548 12316
rect 32508 11354 32536 12310
rect 32600 12306 32628 12582
rect 32588 12300 32640 12306
rect 32588 12242 32640 12248
rect 32600 11694 32628 12242
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32680 11620 32732 11626
rect 32680 11562 32732 11568
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 32324 10798 32444 10826
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32140 9042 32168 10406
rect 32324 10266 32352 10610
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 32416 9722 32444 10798
rect 32692 9722 32720 11562
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32416 9518 32444 9658
rect 32692 9518 32720 9658
rect 32404 9512 32456 9518
rect 32404 9454 32456 9460
rect 32680 9512 32732 9518
rect 32680 9454 32732 9460
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32600 9042 32628 9318
rect 32968 9042 32996 12650
rect 33336 12442 33364 12718
rect 33324 12436 33376 12442
rect 33324 12378 33376 12384
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 33060 10130 33088 11630
rect 33336 11626 33364 12378
rect 33324 11620 33376 11626
rect 33324 11562 33376 11568
rect 33508 11620 33560 11626
rect 33508 11562 33560 11568
rect 33520 10606 33548 11562
rect 33612 11354 33640 18022
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 33704 12374 33732 16526
rect 33888 16114 33916 19110
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 34072 17882 34100 18634
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34164 17270 34192 20198
rect 34532 20058 34560 20266
rect 34520 20052 34572 20058
rect 34520 19994 34572 20000
rect 34532 19310 34560 19994
rect 34612 19712 34664 19718
rect 34612 19654 34664 19660
rect 34716 19666 34744 28358
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 28218 35296 28562
rect 35256 28212 35308 28218
rect 35256 28154 35308 28160
rect 35624 27872 35676 27878
rect 35624 27814 35676 27820
rect 35256 27328 35308 27334
rect 35256 27270 35308 27276
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35268 26994 35296 27270
rect 35256 26988 35308 26994
rect 35256 26930 35308 26936
rect 35636 26518 35664 27814
rect 35716 27464 35768 27470
rect 35716 27406 35768 27412
rect 35624 26512 35676 26518
rect 35624 26454 35676 26460
rect 35624 26240 35676 26246
rect 35728 26228 35756 27406
rect 35676 26200 35756 26228
rect 35624 26182 35676 26188
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35636 26042 35664 26182
rect 35624 26036 35676 26042
rect 35624 25978 35676 25984
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 34808 25809 34836 25842
rect 34794 25800 34850 25809
rect 34794 25735 34850 25744
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 34808 25498 34836 25638
rect 34796 25492 34848 25498
rect 34796 25434 34848 25440
rect 34808 24818 34836 25434
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34796 24812 34848 24818
rect 34796 24754 34848 24760
rect 35360 24449 35388 25638
rect 35532 25288 35584 25294
rect 35532 25230 35584 25236
rect 35440 25220 35492 25226
rect 35440 25162 35492 25168
rect 35452 24818 35480 25162
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 35346 24440 35402 24449
rect 35346 24375 35402 24384
rect 35256 24132 35308 24138
rect 35256 24074 35308 24080
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 35268 23594 35296 24074
rect 35348 23724 35400 23730
rect 35452 23712 35480 24754
rect 35544 24410 35572 25230
rect 35532 24404 35584 24410
rect 35532 24346 35584 24352
rect 35400 23684 35480 23712
rect 35348 23666 35400 23672
rect 35256 23588 35308 23594
rect 35256 23530 35308 23536
rect 35268 23322 35296 23530
rect 35256 23316 35308 23322
rect 35256 23258 35308 23264
rect 35256 22976 35308 22982
rect 35256 22918 35308 22924
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35268 22710 35296 22918
rect 35360 22710 35388 23666
rect 35820 23474 35848 29990
rect 35912 29850 35940 30330
rect 36188 30326 36216 30738
rect 36268 30592 36320 30598
rect 36268 30534 36320 30540
rect 36176 30320 36228 30326
rect 36176 30262 36228 30268
rect 36188 29850 36216 30262
rect 36280 30190 36308 30534
rect 36360 30252 36412 30258
rect 36360 30194 36412 30200
rect 36268 30184 36320 30190
rect 36268 30126 36320 30132
rect 36280 29850 36308 30126
rect 35900 29844 35952 29850
rect 35900 29786 35952 29792
rect 36176 29844 36228 29850
rect 36176 29786 36228 29792
rect 36268 29844 36320 29850
rect 36268 29786 36320 29792
rect 35912 29306 35940 29786
rect 35900 29300 35952 29306
rect 35900 29242 35952 29248
rect 36280 29170 36308 29786
rect 36372 29510 36400 30194
rect 37016 29850 37044 34478
rect 37280 33448 37332 33454
rect 37280 33390 37332 33396
rect 37292 31822 37320 33390
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 37188 31272 37240 31278
rect 37188 31214 37240 31220
rect 37096 30048 37148 30054
rect 37096 29990 37148 29996
rect 37004 29844 37056 29850
rect 37004 29786 37056 29792
rect 36636 29708 36688 29714
rect 36636 29650 36688 29656
rect 36360 29504 36412 29510
rect 36360 29446 36412 29452
rect 36372 29170 36400 29446
rect 36648 29170 36676 29650
rect 37016 29306 37044 29786
rect 37004 29300 37056 29306
rect 37004 29242 37056 29248
rect 36268 29164 36320 29170
rect 36268 29106 36320 29112
rect 36360 29164 36412 29170
rect 36360 29106 36412 29112
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 37004 29164 37056 29170
rect 37004 29106 37056 29112
rect 36372 29073 36400 29106
rect 36358 29064 36414 29073
rect 36084 29028 36136 29034
rect 36358 28999 36414 29008
rect 36084 28970 36136 28976
rect 36096 28626 36124 28970
rect 36084 28620 36136 28626
rect 36084 28562 36136 28568
rect 36096 28529 36124 28562
rect 36082 28520 36138 28529
rect 36082 28455 36138 28464
rect 36372 28218 36400 28999
rect 36360 28212 36412 28218
rect 36360 28154 36412 28160
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 35900 27600 35952 27606
rect 35900 27542 35952 27548
rect 35912 26790 35940 27542
rect 35992 26852 36044 26858
rect 35992 26794 36044 26800
rect 35900 26784 35952 26790
rect 35900 26726 35952 26732
rect 35912 25430 35940 26726
rect 36004 26586 36032 26794
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 36004 26314 36032 26522
rect 36084 26512 36136 26518
rect 36084 26454 36136 26460
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36004 25702 36032 26250
rect 35992 25696 36044 25702
rect 35992 25638 36044 25644
rect 35900 25424 35952 25430
rect 35900 25366 35952 25372
rect 35912 24342 35940 25366
rect 36004 24682 36032 25638
rect 36096 25498 36124 26454
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 36188 24993 36216 27814
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 36372 26382 36400 27406
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36740 26994 36768 27270
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 36360 26376 36412 26382
rect 36360 26318 36412 26324
rect 36268 25356 36320 25362
rect 36268 25298 36320 25304
rect 36174 24984 36230 24993
rect 36174 24919 36230 24928
rect 36280 24886 36308 25298
rect 36268 24880 36320 24886
rect 36268 24822 36320 24828
rect 35992 24676 36044 24682
rect 35992 24618 36044 24624
rect 35900 24336 35952 24342
rect 35952 24296 36032 24324
rect 35900 24278 35952 24284
rect 35900 24064 35952 24070
rect 35900 24006 35952 24012
rect 35912 23798 35940 24006
rect 36004 23798 36032 24296
rect 36176 24200 36228 24206
rect 36176 24142 36228 24148
rect 35900 23792 35952 23798
rect 35900 23734 35952 23740
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 35636 23446 35848 23474
rect 35256 22704 35308 22710
rect 35256 22646 35308 22652
rect 35348 22704 35400 22710
rect 35348 22646 35400 22652
rect 34796 22500 34848 22506
rect 34796 22442 34848 22448
rect 34808 22234 34836 22442
rect 35268 22234 35296 22646
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 35256 22228 35308 22234
rect 35256 22170 35308 22176
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35256 21004 35308 21010
rect 35256 20946 35308 20952
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 34808 20466 34836 20878
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35268 20466 35296 20946
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 35256 20460 35308 20466
rect 35256 20402 35308 20408
rect 35256 19712 35308 19718
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34520 19168 34572 19174
rect 34520 19110 34572 19116
rect 34532 18873 34560 19110
rect 34624 18970 34652 19654
rect 34716 19638 34836 19666
rect 35256 19654 35308 19660
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 34612 18964 34664 18970
rect 34612 18906 34664 18912
rect 34716 18902 34744 19314
rect 34808 18970 34836 19638
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35268 19378 35296 19654
rect 35256 19372 35308 19378
rect 35256 19314 35308 19320
rect 35360 18970 35388 22646
rect 35636 19922 35664 23446
rect 36188 23322 36216 24142
rect 36176 23316 36228 23322
rect 36176 23258 36228 23264
rect 35992 23180 36044 23186
rect 35992 23122 36044 23128
rect 35808 22500 35860 22506
rect 35808 22442 35860 22448
rect 35820 22166 35848 22442
rect 36004 22438 36032 23122
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 35808 22160 35860 22166
rect 35808 22102 35860 22108
rect 35716 22024 35768 22030
rect 35716 21966 35768 21972
rect 35728 21690 35756 21966
rect 35820 21690 35848 22102
rect 36004 22001 36032 22374
rect 36372 22166 36400 26318
rect 36740 26042 36768 26930
rect 36728 26036 36780 26042
rect 36728 25978 36780 25984
rect 36912 25152 36964 25158
rect 36912 25094 36964 25100
rect 36924 24682 36952 25094
rect 36636 24676 36688 24682
rect 36636 24618 36688 24624
rect 36912 24676 36964 24682
rect 36912 24618 36964 24624
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36360 22160 36412 22166
rect 36360 22102 36412 22108
rect 35990 21992 36046 22001
rect 35990 21927 36046 21936
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 35900 21072 35952 21078
rect 35820 21032 35900 21060
rect 35820 20262 35848 21032
rect 35900 21014 35952 21020
rect 36372 20942 36400 22102
rect 36360 20936 36412 20942
rect 36360 20878 36412 20884
rect 35808 20256 35860 20262
rect 35808 20198 35860 20204
rect 35820 20058 35848 20198
rect 36372 20058 36400 20878
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 36360 20052 36412 20058
rect 36360 19994 36412 20000
rect 35624 19916 35676 19922
rect 35624 19858 35676 19864
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 35636 19514 35664 19858
rect 35624 19508 35676 19514
rect 35624 19450 35676 19456
rect 36188 19417 36216 19858
rect 36464 19446 36492 24278
rect 36648 24206 36676 24618
rect 36636 24200 36688 24206
rect 36636 24142 36688 24148
rect 36648 23866 36676 24142
rect 36924 24070 36952 24618
rect 37016 24274 37044 29106
rect 37108 28801 37136 29990
rect 37094 28792 37150 28801
rect 37094 28727 37150 28736
rect 37096 28620 37148 28626
rect 37096 28562 37148 28568
rect 37108 27878 37136 28562
rect 37200 28218 37228 31214
rect 37280 30116 37332 30122
rect 37280 30058 37332 30064
rect 37292 29238 37320 30058
rect 37280 29232 37332 29238
rect 37280 29174 37332 29180
rect 37188 28212 37240 28218
rect 37188 28154 37240 28160
rect 37188 28008 37240 28014
rect 37188 27950 37240 27956
rect 37096 27872 37148 27878
rect 37096 27814 37148 27820
rect 37004 24268 37056 24274
rect 37004 24210 37056 24216
rect 36912 24064 36964 24070
rect 36912 24006 36964 24012
rect 36924 23866 36952 24006
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 36912 23860 36964 23866
rect 36964 23820 37044 23848
rect 36912 23802 36964 23808
rect 37016 23594 37044 23820
rect 36912 23588 36964 23594
rect 36912 23530 36964 23536
rect 37004 23588 37056 23594
rect 37004 23530 37056 23536
rect 36924 23322 36952 23530
rect 37108 23322 37136 27814
rect 37200 25430 37228 27950
rect 37280 25696 37332 25702
rect 37280 25638 37332 25644
rect 37188 25424 37240 25430
rect 37188 25366 37240 25372
rect 37292 24721 37320 25638
rect 37278 24712 37334 24721
rect 37278 24647 37334 24656
rect 37280 24132 37332 24138
rect 37280 24074 37332 24080
rect 37292 23730 37320 24074
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 36912 23316 36964 23322
rect 36912 23258 36964 23264
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 36636 23180 36688 23186
rect 36636 23122 36688 23128
rect 36648 22778 36676 23122
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 36636 22772 36688 22778
rect 36636 22714 36688 22720
rect 37200 22642 37228 22918
rect 37292 22642 37320 23666
rect 37188 22636 37240 22642
rect 37188 22578 37240 22584
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37200 22234 37228 22578
rect 37188 22228 37240 22234
rect 37188 22170 37240 22176
rect 36728 21888 36780 21894
rect 36728 21830 36780 21836
rect 36740 21486 36768 21830
rect 36728 21480 36780 21486
rect 36728 21422 36780 21428
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36648 19446 36676 20334
rect 36740 20262 36768 21422
rect 37292 20942 37320 22578
rect 37280 20936 37332 20942
rect 37280 20878 37332 20884
rect 36820 20392 36872 20398
rect 36820 20334 36872 20340
rect 36728 20256 36780 20262
rect 36728 20198 36780 20204
rect 36452 19440 36504 19446
rect 36174 19408 36230 19417
rect 36174 19343 36230 19352
rect 36358 19408 36414 19417
rect 36452 19382 36504 19388
rect 36636 19440 36688 19446
rect 36636 19382 36688 19388
rect 36358 19343 36414 19352
rect 36188 19310 36216 19343
rect 36176 19304 36228 19310
rect 36176 19246 36228 19252
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 34796 18964 34848 18970
rect 34796 18906 34848 18912
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34704 18896 34756 18902
rect 34518 18864 34574 18873
rect 34336 18828 34388 18834
rect 34704 18838 34756 18844
rect 34518 18799 34574 18808
rect 34336 18770 34388 18776
rect 34348 18086 34376 18770
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 34336 18080 34388 18086
rect 34336 18022 34388 18028
rect 34256 17678 34284 18022
rect 34532 17746 34560 18799
rect 34808 18358 34836 18906
rect 35360 18766 35388 18906
rect 35636 18902 35664 19110
rect 35624 18896 35676 18902
rect 35624 18838 35676 18844
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34796 18352 34848 18358
rect 34796 18294 34848 18300
rect 34808 18222 34836 18294
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 35256 18080 35308 18086
rect 35256 18022 35308 18028
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34244 17672 34296 17678
rect 34244 17614 34296 17620
rect 34532 17338 34560 17682
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34152 17264 34204 17270
rect 34152 17206 34204 17212
rect 34612 17196 34664 17202
rect 34612 17138 34664 17144
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34348 16794 34376 17070
rect 34336 16788 34388 16794
rect 34388 16748 34560 16776
rect 34336 16730 34388 16736
rect 34152 16652 34204 16658
rect 34152 16594 34204 16600
rect 34164 16250 34192 16594
rect 34532 16454 34560 16748
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34152 16244 34204 16250
rect 34152 16186 34204 16192
rect 34244 16176 34296 16182
rect 34244 16118 34296 16124
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33796 15502 33824 15846
rect 33968 15564 34020 15570
rect 33968 15506 34020 15512
rect 33784 15496 33836 15502
rect 33784 15438 33836 15444
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33796 14618 33824 15098
rect 33980 14890 34008 15506
rect 34256 15502 34284 16118
rect 34336 15700 34388 15706
rect 34336 15642 34388 15648
rect 34428 15700 34480 15706
rect 34428 15642 34480 15648
rect 34348 15570 34376 15642
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34244 15496 34296 15502
rect 34244 15438 34296 15444
rect 34256 15162 34284 15438
rect 34348 15366 34376 15506
rect 34336 15360 34388 15366
rect 34336 15302 34388 15308
rect 34244 15156 34296 15162
rect 34244 15098 34296 15104
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33980 14618 34008 14826
rect 34348 14804 34376 15302
rect 34440 15162 34468 15642
rect 34532 15434 34560 16390
rect 34520 15428 34572 15434
rect 34520 15370 34572 15376
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34440 14958 34468 15098
rect 34532 15094 34560 15370
rect 34520 15088 34572 15094
rect 34520 15030 34572 15036
rect 34624 14958 34652 17138
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 34716 15910 34744 15982
rect 34704 15904 34756 15910
rect 34704 15846 34756 15852
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 34612 14952 34664 14958
rect 34612 14894 34664 14900
rect 34348 14776 34560 14804
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 34336 14340 34388 14346
rect 34336 14282 34388 14288
rect 33874 13832 33930 13841
rect 33874 13767 33930 13776
rect 33888 13734 33916 13767
rect 33876 13728 33928 13734
rect 33876 13670 33928 13676
rect 33888 12753 33916 13670
rect 33874 12744 33930 12753
rect 33874 12679 33930 12688
rect 33692 12368 33744 12374
rect 33692 12310 33744 12316
rect 33704 11898 33732 12310
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 33612 10810 33640 11290
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 33508 10600 33560 10606
rect 33508 10542 33560 10548
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 33060 9722 33088 10066
rect 33048 9716 33100 9722
rect 33048 9658 33100 9664
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32588 9036 32640 9042
rect 32588 8978 32640 8984
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32600 8634 32628 8978
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32232 7546 32260 7890
rect 32600 7546 32628 8570
rect 32968 8090 32996 8978
rect 33060 8634 33088 9318
rect 33428 9042 33456 10542
rect 33704 10198 33732 11834
rect 33888 11354 33916 12174
rect 33876 11348 33928 11354
rect 33876 11290 33928 11296
rect 33888 11218 33916 11290
rect 33876 11212 33928 11218
rect 33876 11154 33928 11160
rect 33888 10810 33916 11154
rect 33876 10804 33928 10810
rect 33876 10746 33928 10752
rect 33692 10192 33744 10198
rect 33692 10134 33744 10140
rect 33704 9722 33732 10134
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33416 9036 33468 9042
rect 33416 8978 33468 8984
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 33060 8430 33088 8570
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32220 7540 32272 7546
rect 32220 7482 32272 7488
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32600 7342 32628 7482
rect 32588 7336 32640 7342
rect 32588 7278 32640 7284
rect 32772 7336 32824 7342
rect 32772 7278 32824 7284
rect 32600 6866 32628 7278
rect 32784 7002 32812 7278
rect 32772 6996 32824 7002
rect 32772 6938 32824 6944
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32956 6860 33008 6866
rect 32956 6802 33008 6808
rect 32968 6458 32996 6802
rect 32956 6452 33008 6458
rect 32956 6394 33008 6400
rect 33060 5846 33088 8366
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33336 7410 33364 7822
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 33428 6984 33456 8978
rect 33692 8832 33744 8838
rect 33692 8774 33744 8780
rect 33704 8498 33732 8774
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 34348 8430 34376 14282
rect 34532 13802 34560 14776
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 34624 14074 34652 14350
rect 34716 14074 34744 15846
rect 34612 14068 34664 14074
rect 34612 14010 34664 14016
rect 34704 14068 34756 14074
rect 34704 14010 34756 14016
rect 34808 13814 34836 16934
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 16182 35296 18022
rect 35636 17882 35664 18838
rect 35806 18320 35862 18329
rect 35806 18255 35862 18264
rect 35820 18222 35848 18255
rect 35808 18216 35860 18222
rect 35808 18158 35860 18164
rect 35624 17876 35676 17882
rect 35624 17818 35676 17824
rect 35348 17740 35400 17746
rect 35348 17682 35400 17688
rect 35360 16998 35388 17682
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 35440 17264 35492 17270
rect 35440 17206 35492 17212
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35360 16794 35388 16934
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 35256 16176 35308 16182
rect 35256 16118 35308 16124
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 15144 35296 15302
rect 35176 15116 35296 15144
rect 34980 15088 35032 15094
rect 34980 15030 35032 15036
rect 34992 14260 35020 15030
rect 35176 14890 35204 15116
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 35164 14884 35216 14890
rect 35164 14826 35216 14832
rect 35176 14414 35204 14826
rect 35268 14550 35296 14962
rect 35256 14544 35308 14550
rect 35256 14486 35308 14492
rect 35164 14408 35216 14414
rect 35164 14350 35216 14356
rect 34992 14232 35296 14260
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 35268 13938 35296 14232
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 34520 13796 34572 13802
rect 34520 13738 34572 13744
rect 34716 13786 34836 13814
rect 34532 13530 34560 13738
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34716 13394 34744 13786
rect 35268 13530 35296 13874
rect 35256 13524 35308 13530
rect 35256 13466 35308 13472
rect 34704 13388 34756 13394
rect 34704 13330 34756 13336
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34716 12442 34744 13330
rect 34808 12714 34836 13330
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 35360 12850 35388 15982
rect 35452 15706 35480 17206
rect 35544 17134 35572 17614
rect 36372 17270 36400 19343
rect 36464 18426 36492 19382
rect 36832 18630 36860 20334
rect 36820 18624 36872 18630
rect 36820 18566 36872 18572
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36464 18222 36492 18362
rect 36832 18222 36860 18566
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36820 18216 36872 18222
rect 36820 18158 36872 18164
rect 36912 18216 36964 18222
rect 36912 18158 36964 18164
rect 36464 17882 36492 18158
rect 36452 17876 36504 17882
rect 36452 17818 36504 17824
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36556 17270 36584 17478
rect 36924 17338 36952 18158
rect 37384 17921 37412 38694
rect 37476 34066 37504 43318
rect 37740 38412 37792 38418
rect 37740 38354 37792 38360
rect 37752 37738 37780 38354
rect 37740 37732 37792 37738
rect 37740 37674 37792 37680
rect 37844 37330 37872 44134
rect 38384 43716 38436 43722
rect 38384 43658 38436 43664
rect 38108 43104 38160 43110
rect 38108 43046 38160 43052
rect 38120 42770 38148 43046
rect 38200 42900 38252 42906
rect 38200 42842 38252 42848
rect 38212 42794 38240 42842
rect 38016 42764 38068 42770
rect 38016 42706 38068 42712
rect 38108 42764 38160 42770
rect 38212 42766 38332 42794
rect 38108 42706 38160 42712
rect 37924 42288 37976 42294
rect 37924 42230 37976 42236
rect 37936 41682 37964 42230
rect 38028 42226 38056 42706
rect 38016 42220 38068 42226
rect 38016 42162 38068 42168
rect 38120 41682 38148 42706
rect 38200 42152 38252 42158
rect 38200 42094 38252 42100
rect 38212 41818 38240 42094
rect 38304 42090 38332 42766
rect 38396 42548 38424 43658
rect 38476 43104 38528 43110
rect 38476 43046 38528 43052
rect 38488 42702 38516 43046
rect 38476 42696 38528 42702
rect 38476 42638 38528 42644
rect 38476 42560 38528 42566
rect 38396 42520 38476 42548
rect 38476 42502 38528 42508
rect 38292 42084 38344 42090
rect 38292 42026 38344 42032
rect 38200 41812 38252 41818
rect 38200 41754 38252 41760
rect 37924 41676 37976 41682
rect 37924 41618 37976 41624
rect 38108 41676 38160 41682
rect 38108 41618 38160 41624
rect 37936 41206 37964 41618
rect 38120 41274 38148 41618
rect 38108 41268 38160 41274
rect 38108 41210 38160 41216
rect 37924 41200 37976 41206
rect 37924 41142 37976 41148
rect 38120 41138 38148 41210
rect 38108 41132 38160 41138
rect 38108 41074 38160 41080
rect 38016 40384 38068 40390
rect 38016 40326 38068 40332
rect 37924 40180 37976 40186
rect 37924 40122 37976 40128
rect 37936 39982 37964 40122
rect 38028 39982 38056 40326
rect 37924 39976 37976 39982
rect 37924 39918 37976 39924
rect 38016 39976 38068 39982
rect 38016 39918 38068 39924
rect 38028 39506 38056 39918
rect 38120 39642 38148 41074
rect 38384 40928 38436 40934
rect 38384 40870 38436 40876
rect 38396 40458 38424 40870
rect 38384 40452 38436 40458
rect 38384 40394 38436 40400
rect 38108 39636 38160 39642
rect 38108 39578 38160 39584
rect 38016 39500 38068 39506
rect 38016 39442 38068 39448
rect 38028 38758 38056 39442
rect 38120 39098 38148 39578
rect 38108 39092 38160 39098
rect 38108 39034 38160 39040
rect 38016 38752 38068 38758
rect 38016 38694 38068 38700
rect 38028 38554 38056 38694
rect 38016 38548 38068 38554
rect 38016 38490 38068 38496
rect 38028 38418 38056 38490
rect 38016 38412 38068 38418
rect 38016 38354 38068 38360
rect 38292 37800 38344 37806
rect 38396 37788 38424 40394
rect 38488 37890 38516 42502
rect 38580 40050 38608 44270
rect 39316 43926 39344 44814
rect 39592 44538 39620 45222
rect 40604 45082 40632 45426
rect 40696 45354 40724 45766
rect 40684 45348 40736 45354
rect 40684 45290 40736 45296
rect 41512 45348 41564 45354
rect 41512 45290 41564 45296
rect 40592 45076 40644 45082
rect 40592 45018 40644 45024
rect 39948 45008 40000 45014
rect 39948 44950 40000 44956
rect 40224 45008 40276 45014
rect 40224 44950 40276 44956
rect 39580 44532 39632 44538
rect 39580 44474 39632 44480
rect 39960 44470 39988 44950
rect 40236 44742 40264 44950
rect 41524 44878 41552 45290
rect 41616 45286 41644 46038
rect 41708 45830 41736 46378
rect 41788 45960 41840 45966
rect 41788 45902 41840 45908
rect 41696 45824 41748 45830
rect 41696 45766 41748 45772
rect 41800 45558 41828 45902
rect 42352 45898 42380 46378
rect 43732 46170 43760 49558
rect 49514 48512 49570 48521
rect 49514 48447 49570 48456
rect 43720 46164 43772 46170
rect 43720 46106 43772 46112
rect 42340 45892 42392 45898
rect 42340 45834 42392 45840
rect 42156 45824 42208 45830
rect 42156 45766 42208 45772
rect 42168 45626 42196 45766
rect 42156 45620 42208 45626
rect 42156 45562 42208 45568
rect 41788 45552 41840 45558
rect 41788 45494 41840 45500
rect 41604 45280 41656 45286
rect 41604 45222 41656 45228
rect 41616 45014 41644 45222
rect 41604 45008 41656 45014
rect 41604 44950 41656 44956
rect 41512 44872 41564 44878
rect 41512 44814 41564 44820
rect 41328 44804 41380 44810
rect 41328 44746 41380 44752
rect 40224 44736 40276 44742
rect 40224 44678 40276 44684
rect 40236 44538 40264 44678
rect 40224 44532 40276 44538
rect 40224 44474 40276 44480
rect 39948 44464 40000 44470
rect 39948 44406 40000 44412
rect 39304 43920 39356 43926
rect 39304 43862 39356 43868
rect 38936 43852 38988 43858
rect 38936 43794 38988 43800
rect 38948 43246 38976 43794
rect 39764 43308 39816 43314
rect 39764 43250 39816 43256
rect 38936 43240 38988 43246
rect 38856 43200 38936 43228
rect 38856 42770 38884 43200
rect 38936 43182 38988 43188
rect 39488 43104 39540 43110
rect 39488 43046 39540 43052
rect 38844 42764 38896 42770
rect 38844 42706 38896 42712
rect 39212 42696 39264 42702
rect 39212 42638 39264 42644
rect 39224 41818 39252 42638
rect 39500 42226 39528 43046
rect 39488 42220 39540 42226
rect 39488 42162 39540 42168
rect 39212 41812 39264 41818
rect 39212 41754 39264 41760
rect 38936 41132 38988 41138
rect 38936 41074 38988 41080
rect 38948 40730 38976 41074
rect 39120 40928 39172 40934
rect 39120 40870 39172 40876
rect 38936 40724 38988 40730
rect 38936 40666 38988 40672
rect 38936 40588 38988 40594
rect 38936 40530 38988 40536
rect 38568 40044 38620 40050
rect 38568 39986 38620 39992
rect 38948 39846 38976 40530
rect 39132 40050 39160 40870
rect 39500 40633 39528 42162
rect 39776 42129 39804 43250
rect 39762 42120 39818 42129
rect 39762 42055 39818 42064
rect 39580 42016 39632 42022
rect 39580 41958 39632 41964
rect 39592 41274 39620 41958
rect 39580 41268 39632 41274
rect 39580 41210 39632 41216
rect 39672 41064 39724 41070
rect 39672 41006 39724 41012
rect 39486 40624 39542 40633
rect 39486 40559 39542 40568
rect 39580 40588 39632 40594
rect 39120 40044 39172 40050
rect 39120 39986 39172 39992
rect 38936 39840 38988 39846
rect 38936 39782 38988 39788
rect 38948 39574 38976 39782
rect 39132 39642 39160 39986
rect 39120 39636 39172 39642
rect 39120 39578 39172 39584
rect 38660 39568 38712 39574
rect 38660 39510 38712 39516
rect 38936 39568 38988 39574
rect 38936 39510 38988 39516
rect 38488 37862 38608 37890
rect 38344 37760 38424 37788
rect 38476 37800 38528 37806
rect 38292 37742 38344 37748
rect 38476 37742 38528 37748
rect 37832 37324 37884 37330
rect 37832 37266 37884 37272
rect 37844 36854 37872 37266
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 37832 36848 37884 36854
rect 37832 36790 37884 36796
rect 38212 36786 38240 37062
rect 38200 36780 38252 36786
rect 38200 36722 38252 36728
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 37648 35828 37700 35834
rect 37648 35770 37700 35776
rect 37464 34060 37516 34066
rect 37464 34002 37516 34008
rect 37464 32972 37516 32978
rect 37464 32914 37516 32920
rect 37476 32570 37504 32914
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37464 31272 37516 31278
rect 37464 31214 37516 31220
rect 37476 30666 37504 31214
rect 37556 31204 37608 31210
rect 37556 31146 37608 31152
rect 37464 30660 37516 30666
rect 37464 30602 37516 30608
rect 37476 30394 37504 30602
rect 37464 30388 37516 30394
rect 37464 30330 37516 30336
rect 37568 30297 37596 31146
rect 37554 30288 37610 30297
rect 37554 30223 37610 30232
rect 37556 30184 37608 30190
rect 37556 30126 37608 30132
rect 37568 29782 37596 30126
rect 37556 29776 37608 29782
rect 37556 29718 37608 29724
rect 37462 29608 37518 29617
rect 37462 29543 37518 29552
rect 37476 29510 37504 29543
rect 37464 29504 37516 29510
rect 37464 29446 37516 29452
rect 37660 28762 37688 35770
rect 37844 34513 37872 36518
rect 38108 35624 38160 35630
rect 38108 35566 38160 35572
rect 38016 35556 38068 35562
rect 38016 35498 38068 35504
rect 38028 35222 38056 35498
rect 38016 35216 38068 35222
rect 37936 35176 38016 35204
rect 37936 34746 37964 35176
rect 38016 35158 38068 35164
rect 38016 35080 38068 35086
rect 38016 35022 38068 35028
rect 37924 34740 37976 34746
rect 37924 34682 37976 34688
rect 38028 34610 38056 35022
rect 38016 34604 38068 34610
rect 38016 34546 38068 34552
rect 37830 34504 37886 34513
rect 37830 34439 37886 34448
rect 37740 31680 37792 31686
rect 37740 31622 37792 31628
rect 37752 30394 37780 31622
rect 37844 31346 37872 34439
rect 38028 34202 38056 34546
rect 38016 34196 38068 34202
rect 38016 34138 38068 34144
rect 38120 33114 38148 35566
rect 38200 35488 38252 35494
rect 38200 35430 38252 35436
rect 38212 34202 38240 35430
rect 38200 34196 38252 34202
rect 38200 34138 38252 34144
rect 38200 33312 38252 33318
rect 38200 33254 38252 33260
rect 38212 33153 38240 33254
rect 38198 33144 38254 33153
rect 38108 33108 38160 33114
rect 38198 33079 38254 33088
rect 38108 33050 38160 33056
rect 38200 32972 38252 32978
rect 38200 32914 38252 32920
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38016 32768 38068 32774
rect 38016 32710 38068 32716
rect 38028 32434 38056 32710
rect 38016 32428 38068 32434
rect 38016 32370 38068 32376
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 37832 31340 37884 31346
rect 37832 31282 37884 31288
rect 37740 30388 37792 30394
rect 37740 30330 37792 30336
rect 37752 29578 37780 30330
rect 37740 29572 37792 29578
rect 37740 29514 37792 29520
rect 37648 28756 37700 28762
rect 37648 28698 37700 28704
rect 37740 28620 37792 28626
rect 37740 28562 37792 28568
rect 37556 28008 37608 28014
rect 37556 27950 37608 27956
rect 37464 27056 37516 27062
rect 37464 26998 37516 27004
rect 37476 24818 37504 26998
rect 37464 24812 37516 24818
rect 37464 24754 37516 24760
rect 37568 22438 37596 27950
rect 37752 27878 37780 28562
rect 37740 27872 37792 27878
rect 37740 27814 37792 27820
rect 37936 26432 37964 32166
rect 38120 31890 38148 32846
rect 38212 32570 38240 32914
rect 38200 32564 38252 32570
rect 38200 32506 38252 32512
rect 38212 32366 38240 32506
rect 38200 32360 38252 32366
rect 38200 32302 38252 32308
rect 38108 31884 38160 31890
rect 38108 31826 38160 31832
rect 38120 31482 38148 31826
rect 38108 31476 38160 31482
rect 38108 31418 38160 31424
rect 38304 31278 38332 37742
rect 38488 37126 38516 37742
rect 38476 37120 38528 37126
rect 38476 37062 38528 37068
rect 38580 36718 38608 37862
rect 38568 36712 38620 36718
rect 38568 36654 38620 36660
rect 38568 36032 38620 36038
rect 38568 35974 38620 35980
rect 38580 35494 38608 35974
rect 38672 35766 38700 39510
rect 38752 39432 38804 39438
rect 38752 39374 38804 39380
rect 38764 38486 38792 39374
rect 38844 38888 38896 38894
rect 38844 38830 38896 38836
rect 38856 38554 38884 38830
rect 39132 38826 39160 39578
rect 39120 38820 39172 38826
rect 39120 38762 39172 38768
rect 38844 38548 38896 38554
rect 38844 38490 38896 38496
rect 38752 38480 38804 38486
rect 38752 38422 38804 38428
rect 38856 36242 38884 38490
rect 39028 38412 39080 38418
rect 39028 38354 39080 38360
rect 39040 38010 39068 38354
rect 39028 38004 39080 38010
rect 39028 37946 39080 37952
rect 38936 37732 38988 37738
rect 38936 37674 38988 37680
rect 38948 37262 38976 37674
rect 39132 37466 39160 38762
rect 39120 37460 39172 37466
rect 39120 37402 39172 37408
rect 38936 37256 38988 37262
rect 38936 37198 38988 37204
rect 38948 36378 38976 37198
rect 39028 37120 39080 37126
rect 39028 37062 39080 37068
rect 39040 36718 39068 37062
rect 39132 36854 39160 37402
rect 39120 36848 39172 36854
rect 39120 36790 39172 36796
rect 39028 36712 39080 36718
rect 39028 36654 39080 36660
rect 38936 36372 38988 36378
rect 38936 36314 38988 36320
rect 38844 36236 38896 36242
rect 38844 36178 38896 36184
rect 38856 35834 38884 36178
rect 39040 36174 39068 36654
rect 39028 36168 39080 36174
rect 39028 36110 39080 36116
rect 38844 35828 38896 35834
rect 38844 35770 38896 35776
rect 39500 35766 39528 40559
rect 39580 40530 39632 40536
rect 39592 40186 39620 40530
rect 39684 40526 39712 41006
rect 39672 40520 39724 40526
rect 39672 40462 39724 40468
rect 39580 40180 39632 40186
rect 39580 40122 39632 40128
rect 39580 39976 39632 39982
rect 39580 39918 39632 39924
rect 39592 38962 39620 39918
rect 39580 38956 39632 38962
rect 39580 38898 39632 38904
rect 39672 38344 39724 38350
rect 39776 38332 39804 42055
rect 39960 42022 39988 44406
rect 41340 44198 41368 44746
rect 41328 44192 41380 44198
rect 41328 44134 41380 44140
rect 41340 43994 41368 44134
rect 41328 43988 41380 43994
rect 41328 43930 41380 43936
rect 41052 43852 41104 43858
rect 41052 43794 41104 43800
rect 41064 43314 41092 43794
rect 41052 43308 41104 43314
rect 41052 43250 41104 43256
rect 40868 43104 40920 43110
rect 40868 43046 40920 43052
rect 40776 42900 40828 42906
rect 40776 42842 40828 42848
rect 40316 42628 40368 42634
rect 40316 42570 40368 42576
rect 40132 42560 40184 42566
rect 40132 42502 40184 42508
rect 40144 42362 40172 42502
rect 40132 42356 40184 42362
rect 40132 42298 40184 42304
rect 40144 42090 40172 42298
rect 40132 42084 40184 42090
rect 40132 42026 40184 42032
rect 39948 42016 40000 42022
rect 39948 41958 40000 41964
rect 39960 41750 39988 41958
rect 39948 41744 40000 41750
rect 39948 41686 40000 41692
rect 39856 41608 39908 41614
rect 39856 41550 39908 41556
rect 39868 41138 39896 41550
rect 39856 41132 39908 41138
rect 39856 41074 39908 41080
rect 39960 40934 39988 41686
rect 39948 40928 40000 40934
rect 39948 40870 40000 40876
rect 39856 40520 39908 40526
rect 39856 40462 39908 40468
rect 39868 39506 39896 40462
rect 39856 39500 39908 39506
rect 39856 39442 39908 39448
rect 40224 39500 40276 39506
rect 40224 39442 40276 39448
rect 40236 39098 40264 39442
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 40328 38418 40356 42570
rect 40788 42226 40816 42842
rect 40880 42838 40908 43046
rect 41524 42906 41552 44814
rect 41800 44538 41828 45494
rect 42168 44538 42196 45562
rect 41788 44532 41840 44538
rect 41788 44474 41840 44480
rect 42156 44532 42208 44538
rect 42156 44474 42208 44480
rect 42156 44192 42208 44198
rect 42156 44134 42208 44140
rect 41878 43888 41934 43897
rect 41878 43823 41934 43832
rect 41892 43790 41920 43823
rect 41880 43784 41932 43790
rect 41880 43726 41932 43732
rect 42168 43722 42196 44134
rect 42156 43716 42208 43722
rect 42156 43658 42208 43664
rect 41788 43648 41840 43654
rect 41788 43590 41840 43596
rect 41800 43314 41828 43590
rect 42168 43450 42196 43658
rect 42156 43444 42208 43450
rect 42156 43386 42208 43392
rect 41788 43308 41840 43314
rect 41788 43250 41840 43256
rect 42064 43172 42116 43178
rect 42064 43114 42116 43120
rect 41788 43104 41840 43110
rect 41788 43046 41840 43052
rect 41512 42900 41564 42906
rect 41512 42842 41564 42848
rect 40868 42832 40920 42838
rect 40868 42774 40920 42780
rect 41144 42832 41196 42838
rect 41144 42774 41196 42780
rect 40776 42220 40828 42226
rect 40776 42162 40828 42168
rect 40880 41818 40908 42774
rect 41156 42004 41184 42774
rect 41800 42634 41828 43046
rect 41788 42628 41840 42634
rect 41788 42570 41840 42576
rect 41328 42016 41380 42022
rect 41156 41976 41328 42004
rect 41328 41958 41380 41964
rect 40868 41812 40920 41818
rect 40868 41754 40920 41760
rect 40776 41744 40828 41750
rect 40776 41686 40828 41692
rect 40788 41274 40816 41686
rect 40776 41268 40828 41274
rect 40776 41210 40828 41216
rect 40500 40384 40552 40390
rect 40500 40326 40552 40332
rect 40512 39982 40540 40326
rect 40500 39976 40552 39982
rect 40500 39918 40552 39924
rect 40776 39908 40828 39914
rect 40776 39850 40828 39856
rect 40788 39574 40816 39850
rect 41340 39846 41368 41958
rect 41800 41614 41828 42570
rect 41972 42084 42024 42090
rect 41972 42026 42024 42032
rect 41984 41750 42012 42026
rect 42076 42022 42104 43114
rect 42352 43110 42380 45834
rect 42524 45620 42576 45626
rect 42524 45562 42576 45568
rect 42432 45484 42484 45490
rect 42432 45426 42484 45432
rect 42444 45082 42472 45426
rect 42536 45354 42564 45562
rect 42524 45348 42576 45354
rect 42524 45290 42576 45296
rect 43720 45348 43772 45354
rect 43720 45290 43772 45296
rect 42432 45076 42484 45082
rect 42432 45018 42484 45024
rect 43732 44878 43760 45290
rect 43812 45280 43864 45286
rect 43812 45222 43864 45228
rect 44824 45280 44876 45286
rect 44824 45222 44876 45228
rect 43824 45014 43852 45222
rect 43812 45008 43864 45014
rect 43812 44950 43864 44956
rect 43444 44872 43496 44878
rect 43720 44872 43772 44878
rect 43444 44814 43496 44820
rect 43548 44832 43720 44860
rect 42708 44396 42760 44402
rect 42708 44338 42760 44344
rect 42720 43994 42748 44338
rect 43456 44266 43484 44814
rect 43444 44260 43496 44266
rect 43444 44202 43496 44208
rect 42708 43988 42760 43994
rect 42708 43930 42760 43936
rect 43456 43926 43484 44202
rect 43444 43920 43496 43926
rect 43444 43862 43496 43868
rect 42524 43852 42576 43858
rect 42524 43794 42576 43800
rect 42536 43178 42564 43794
rect 42708 43716 42760 43722
rect 42708 43658 42760 43664
rect 42616 43240 42668 43246
rect 42616 43182 42668 43188
rect 42524 43172 42576 43178
rect 42524 43114 42576 43120
rect 42340 43104 42392 43110
rect 42340 43046 42392 43052
rect 42628 42702 42656 43182
rect 42616 42696 42668 42702
rect 42616 42638 42668 42644
rect 42340 42560 42392 42566
rect 42340 42502 42392 42508
rect 42352 42090 42380 42502
rect 42340 42084 42392 42090
rect 42340 42026 42392 42032
rect 42064 42016 42116 42022
rect 42064 41958 42116 41964
rect 41972 41744 42024 41750
rect 41972 41686 42024 41692
rect 41604 41608 41656 41614
rect 41604 41550 41656 41556
rect 41788 41608 41840 41614
rect 41788 41550 41840 41556
rect 41420 41064 41472 41070
rect 41420 41006 41472 41012
rect 41328 39840 41380 39846
rect 41328 39782 41380 39788
rect 41340 39642 41368 39782
rect 41328 39636 41380 39642
rect 41328 39578 41380 39584
rect 40776 39568 40828 39574
rect 40776 39510 40828 39516
rect 40788 39098 40816 39510
rect 41432 39098 41460 41006
rect 41616 40730 41644 41550
rect 42076 41546 42104 41958
rect 42064 41540 42116 41546
rect 42064 41482 42116 41488
rect 42352 41274 42380 42026
rect 42616 41744 42668 41750
rect 42616 41686 42668 41692
rect 42340 41268 42392 41274
rect 42340 41210 42392 41216
rect 42628 41206 42656 41686
rect 42616 41200 42668 41206
rect 42616 41142 42668 41148
rect 42522 41032 42578 41041
rect 42522 40967 42578 40976
rect 41696 40928 41748 40934
rect 41696 40870 41748 40876
rect 41604 40724 41656 40730
rect 41604 40666 41656 40672
rect 41708 40186 41736 40870
rect 41880 40656 41932 40662
rect 41880 40598 41932 40604
rect 42432 40656 42484 40662
rect 42432 40598 42484 40604
rect 41788 40520 41840 40526
rect 41788 40462 41840 40468
rect 41800 40186 41828 40462
rect 41696 40180 41748 40186
rect 41696 40122 41748 40128
rect 41788 40180 41840 40186
rect 41788 40122 41840 40128
rect 41892 40050 41920 40598
rect 42248 40112 42300 40118
rect 42248 40054 42300 40060
rect 41880 40044 41932 40050
rect 41880 39986 41932 39992
rect 41892 39642 41920 39986
rect 41880 39636 41932 39642
rect 41880 39578 41932 39584
rect 41788 39568 41840 39574
rect 41788 39510 41840 39516
rect 40776 39092 40828 39098
rect 40776 39034 40828 39040
rect 41420 39092 41472 39098
rect 41420 39034 41472 39040
rect 41432 38894 41460 39034
rect 41800 38894 41828 39510
rect 42260 39506 42288 40054
rect 42444 39574 42472 40598
rect 42432 39568 42484 39574
rect 42432 39510 42484 39516
rect 42248 39500 42300 39506
rect 42300 39460 42380 39488
rect 42248 39442 42300 39448
rect 41236 38888 41288 38894
rect 41236 38830 41288 38836
rect 41420 38888 41472 38894
rect 41420 38830 41472 38836
rect 41788 38888 41840 38894
rect 41788 38830 41840 38836
rect 40960 38752 41012 38758
rect 40960 38694 41012 38700
rect 40972 38486 41000 38694
rect 40960 38480 41012 38486
rect 40960 38422 41012 38428
rect 40316 38412 40368 38418
rect 40316 38354 40368 38360
rect 39724 38304 39804 38332
rect 39672 38286 39724 38292
rect 39684 37670 39712 38286
rect 40328 38010 40356 38354
rect 40592 38208 40644 38214
rect 40592 38150 40644 38156
rect 40868 38208 40920 38214
rect 40868 38150 40920 38156
rect 41052 38208 41104 38214
rect 41052 38150 41104 38156
rect 40316 38004 40368 38010
rect 40316 37946 40368 37952
rect 40604 37874 40632 38150
rect 40592 37868 40644 37874
rect 40592 37810 40644 37816
rect 39764 37732 39816 37738
rect 39764 37674 39816 37680
rect 39672 37664 39724 37670
rect 39672 37606 39724 37612
rect 38660 35760 38712 35766
rect 38660 35702 38712 35708
rect 39488 35760 39540 35766
rect 39488 35702 39540 35708
rect 38568 35488 38620 35494
rect 38568 35430 38620 35436
rect 38580 35290 38608 35430
rect 38568 35284 38620 35290
rect 38568 35226 38620 35232
rect 38580 34474 38608 35226
rect 38660 34536 38712 34542
rect 38660 34478 38712 34484
rect 38568 34468 38620 34474
rect 38568 34410 38620 34416
rect 38580 34066 38608 34410
rect 38672 34134 38700 34478
rect 38660 34128 38712 34134
rect 38660 34070 38712 34076
rect 38476 34060 38528 34066
rect 38476 34002 38528 34008
rect 38568 34060 38620 34066
rect 38568 34002 38620 34008
rect 38488 33658 38516 34002
rect 38476 33652 38528 33658
rect 38476 33594 38528 33600
rect 38292 31272 38344 31278
rect 38292 31214 38344 31220
rect 38016 30796 38068 30802
rect 38016 30738 38068 30744
rect 38028 30394 38056 30738
rect 38304 30598 38332 31214
rect 38292 30592 38344 30598
rect 38292 30534 38344 30540
rect 38016 30388 38068 30394
rect 38016 30330 38068 30336
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 38028 29170 38056 29446
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 38304 28762 38332 30534
rect 38488 30394 38516 33594
rect 38580 33590 38608 34002
rect 38568 33584 38620 33590
rect 38568 33526 38620 33532
rect 39396 33584 39448 33590
rect 39396 33526 39448 33532
rect 39212 33516 39264 33522
rect 39212 33458 39264 33464
rect 38936 33108 38988 33114
rect 38936 33050 38988 33056
rect 38660 32292 38712 32298
rect 38660 32234 38712 32240
rect 38672 31958 38700 32234
rect 38660 31952 38712 31958
rect 38660 31894 38712 31900
rect 38672 31142 38700 31894
rect 38844 31272 38896 31278
rect 38844 31214 38896 31220
rect 38660 31136 38712 31142
rect 38660 31078 38712 31084
rect 38476 30388 38528 30394
rect 38476 30330 38528 30336
rect 38488 30190 38516 30330
rect 38476 30184 38528 30190
rect 38476 30126 38528 30132
rect 38672 29850 38700 31078
rect 38856 30734 38884 31214
rect 38948 30802 38976 33050
rect 38936 30796 38988 30802
rect 38936 30738 38988 30744
rect 38844 30728 38896 30734
rect 38844 30670 38896 30676
rect 38660 29844 38712 29850
rect 38660 29786 38712 29792
rect 38384 29640 38436 29646
rect 38384 29582 38436 29588
rect 38396 29102 38424 29582
rect 38384 29096 38436 29102
rect 38384 29038 38436 29044
rect 38396 28762 38424 29038
rect 38672 28966 38700 29786
rect 39028 29232 39080 29238
rect 39028 29174 39080 29180
rect 38660 28960 38712 28966
rect 38660 28902 38712 28908
rect 38936 28960 38988 28966
rect 38936 28902 38988 28908
rect 38948 28762 38976 28902
rect 38292 28756 38344 28762
rect 38292 28698 38344 28704
rect 38384 28756 38436 28762
rect 38384 28698 38436 28704
rect 38936 28756 38988 28762
rect 38936 28698 38988 28704
rect 38476 28416 38528 28422
rect 38476 28358 38528 28364
rect 38488 28014 38516 28358
rect 38476 28008 38528 28014
rect 38476 27950 38528 27956
rect 38752 28008 38804 28014
rect 38752 27950 38804 27956
rect 38488 27674 38516 27950
rect 38764 27674 38792 27950
rect 38844 27872 38896 27878
rect 38844 27814 38896 27820
rect 38476 27668 38528 27674
rect 38476 27610 38528 27616
rect 38752 27668 38804 27674
rect 38752 27610 38804 27616
rect 38108 27532 38160 27538
rect 38108 27474 38160 27480
rect 38120 27130 38148 27474
rect 38108 27124 38160 27130
rect 38108 27066 38160 27072
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38016 26444 38068 26450
rect 37936 26404 38016 26432
rect 38016 26386 38068 26392
rect 38028 25702 38056 26386
rect 38396 26246 38424 26930
rect 38474 26888 38530 26897
rect 38474 26823 38530 26832
rect 38384 26240 38436 26246
rect 38384 26182 38436 26188
rect 38016 25696 38068 25702
rect 38016 25638 38068 25644
rect 37830 25392 37886 25401
rect 37830 25327 37832 25336
rect 37884 25327 37886 25336
rect 37832 25298 37884 25304
rect 37844 24954 37872 25298
rect 37832 24948 37884 24954
rect 37832 24890 37884 24896
rect 37648 24812 37700 24818
rect 37648 24754 37700 24760
rect 37556 22432 37608 22438
rect 37556 22374 37608 22380
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37476 20058 37504 21830
rect 37568 21554 37596 22374
rect 37660 22234 37688 24754
rect 37924 24268 37976 24274
rect 37924 24210 37976 24216
rect 37936 23866 37964 24210
rect 37924 23860 37976 23866
rect 37924 23802 37976 23808
rect 38028 23474 38056 25638
rect 38396 25498 38424 26182
rect 38488 25838 38516 26823
rect 38764 25838 38792 27610
rect 38856 26450 38884 27814
rect 38948 27674 38976 28698
rect 39040 28082 39068 29174
rect 39028 28076 39080 28082
rect 39028 28018 39080 28024
rect 38936 27668 38988 27674
rect 38936 27610 38988 27616
rect 38844 26444 38896 26450
rect 38844 26386 38896 26392
rect 38476 25832 38528 25838
rect 38476 25774 38528 25780
rect 38752 25832 38804 25838
rect 38752 25774 38804 25780
rect 38384 25492 38436 25498
rect 38384 25434 38436 25440
rect 38292 25424 38344 25430
rect 38292 25366 38344 25372
rect 38108 25288 38160 25294
rect 38108 25230 38160 25236
rect 37936 23446 38056 23474
rect 37740 23180 37792 23186
rect 37740 23122 37792 23128
rect 37752 22710 37780 23122
rect 37936 23118 37964 23446
rect 37924 23112 37976 23118
rect 37924 23054 37976 23060
rect 37740 22704 37792 22710
rect 37740 22646 37792 22652
rect 37648 22228 37700 22234
rect 37648 22170 37700 22176
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37568 21078 37596 21286
rect 37556 21072 37608 21078
rect 37556 21014 37608 21020
rect 37568 20602 37596 21014
rect 37556 20596 37608 20602
rect 37556 20538 37608 20544
rect 37464 20052 37516 20058
rect 37464 19994 37516 20000
rect 37660 19378 37688 22170
rect 37752 21321 37780 22646
rect 37832 22500 37884 22506
rect 37832 22442 37884 22448
rect 37844 22166 37872 22442
rect 37832 22160 37884 22166
rect 37832 22102 37884 22108
rect 37844 21690 37872 22102
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 37738 21312 37794 21321
rect 37738 21247 37794 21256
rect 37844 21146 37872 21626
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37936 19378 37964 23054
rect 38120 21690 38148 25230
rect 38200 23044 38252 23050
rect 38200 22986 38252 22992
rect 38212 22778 38240 22986
rect 38200 22772 38252 22778
rect 38200 22714 38252 22720
rect 38108 21684 38160 21690
rect 38108 21626 38160 21632
rect 38016 21412 38068 21418
rect 38016 21354 38068 21360
rect 38028 20262 38056 21354
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 38120 20602 38148 20878
rect 38108 20596 38160 20602
rect 38108 20538 38160 20544
rect 38016 20256 38068 20262
rect 38016 20198 38068 20204
rect 37648 19372 37700 19378
rect 37648 19314 37700 19320
rect 37924 19372 37976 19378
rect 37924 19314 37976 19320
rect 37464 19236 37516 19242
rect 37464 19178 37516 19184
rect 37556 19236 37608 19242
rect 37556 19178 37608 19184
rect 37476 18272 37504 19178
rect 37568 18970 37596 19178
rect 37556 18964 37608 18970
rect 37556 18906 37608 18912
rect 37660 18902 37688 19314
rect 38028 18902 38056 20198
rect 38212 19242 38240 20878
rect 38200 19236 38252 19242
rect 38200 19178 38252 19184
rect 37648 18896 37700 18902
rect 37648 18838 37700 18844
rect 38016 18896 38068 18902
rect 38016 18838 38068 18844
rect 37740 18760 37792 18766
rect 37740 18702 37792 18708
rect 37752 18426 37780 18702
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 38028 18358 38056 18838
rect 38212 18834 38240 19178
rect 38200 18828 38252 18834
rect 38200 18770 38252 18776
rect 38016 18352 38068 18358
rect 38016 18294 38068 18300
rect 37556 18284 37608 18290
rect 37476 18244 37556 18272
rect 37556 18226 37608 18232
rect 38028 18154 38056 18294
rect 37648 18148 37700 18154
rect 37648 18090 37700 18096
rect 38016 18148 38068 18154
rect 38016 18090 38068 18096
rect 37370 17912 37426 17921
rect 37370 17847 37426 17856
rect 37660 17746 37688 18090
rect 37648 17740 37700 17746
rect 37648 17682 37700 17688
rect 37660 17338 37688 17682
rect 37924 17536 37976 17542
rect 37924 17478 37976 17484
rect 36912 17332 36964 17338
rect 36912 17274 36964 17280
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 36360 17264 36412 17270
rect 36360 17206 36412 17212
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36372 17134 36400 17206
rect 35532 17128 35584 17134
rect 35532 17070 35584 17076
rect 36360 17128 36412 17134
rect 36360 17070 36412 17076
rect 35544 16454 35572 17070
rect 36360 16992 36412 16998
rect 35806 16960 35862 16969
rect 36360 16934 36412 16940
rect 35806 16895 35862 16904
rect 35820 16658 35848 16895
rect 35808 16652 35860 16658
rect 35808 16594 35860 16600
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35440 15700 35492 15706
rect 35440 15642 35492 15648
rect 35452 15570 35480 15642
rect 35544 15638 35572 16390
rect 35820 16250 35848 16594
rect 36372 16250 36400 16934
rect 36556 16726 36584 17206
rect 37936 16794 37964 17478
rect 36912 16788 36964 16794
rect 36912 16730 36964 16736
rect 37924 16788 37976 16794
rect 37924 16730 37976 16736
rect 36544 16720 36596 16726
rect 36544 16662 36596 16668
rect 35808 16244 35860 16250
rect 35808 16186 35860 16192
rect 36360 16244 36412 16250
rect 36360 16186 36412 16192
rect 35532 15632 35584 15638
rect 35532 15574 35584 15580
rect 35440 15564 35492 15570
rect 35440 15506 35492 15512
rect 35544 15162 35572 15574
rect 36452 15564 36504 15570
rect 36452 15506 36504 15512
rect 35532 15156 35584 15162
rect 35532 15098 35584 15104
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35452 14006 35480 14894
rect 35544 14618 35572 15098
rect 35624 14884 35676 14890
rect 35624 14826 35676 14832
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35636 14482 35664 14826
rect 36464 14618 36492 15506
rect 36556 15502 36584 16662
rect 36924 16046 36952 16730
rect 38028 16726 38056 18090
rect 38304 18086 38332 25366
rect 38488 25294 38516 25774
rect 38856 25702 38884 26386
rect 38844 25696 38896 25702
rect 38844 25638 38896 25644
rect 38476 25288 38528 25294
rect 38476 25230 38528 25236
rect 38384 25220 38436 25226
rect 38384 25162 38436 25168
rect 38396 24818 38424 25162
rect 38384 24812 38436 24818
rect 38384 24754 38436 24760
rect 38476 24812 38528 24818
rect 38476 24754 38528 24760
rect 38384 24268 38436 24274
rect 38384 24210 38436 24216
rect 38396 23866 38424 24210
rect 38384 23860 38436 23866
rect 38384 23802 38436 23808
rect 38488 23730 38516 24754
rect 38476 23724 38528 23730
rect 38476 23666 38528 23672
rect 38660 23656 38712 23662
rect 38658 23624 38660 23633
rect 38712 23624 38714 23633
rect 38658 23559 38714 23568
rect 38672 23526 38700 23559
rect 38660 23520 38712 23526
rect 38660 23462 38712 23468
rect 38856 23254 38884 25638
rect 38844 23248 38896 23254
rect 38844 23190 38896 23196
rect 38384 21344 38436 21350
rect 38384 21286 38436 21292
rect 38396 19786 38424 21286
rect 38856 20602 38884 23190
rect 38936 23112 38988 23118
rect 38936 23054 38988 23060
rect 38948 22778 38976 23054
rect 38936 22772 38988 22778
rect 38936 22714 38988 22720
rect 39040 21010 39068 28018
rect 39224 26382 39252 33458
rect 39408 30938 39436 33526
rect 39684 33134 39712 37606
rect 39776 37466 39804 37674
rect 39764 37460 39816 37466
rect 39764 37402 39816 37408
rect 40684 37392 40736 37398
rect 40684 37334 40736 37340
rect 40592 37256 40644 37262
rect 40592 37198 40644 37204
rect 40604 36650 40632 37198
rect 40696 36718 40724 37334
rect 40684 36712 40736 36718
rect 40684 36654 40736 36660
rect 40592 36644 40644 36650
rect 40592 36586 40644 36592
rect 40040 36576 40092 36582
rect 40040 36518 40092 36524
rect 39856 36168 39908 36174
rect 39856 36110 39908 36116
rect 39868 35154 39896 36110
rect 39948 35624 40000 35630
rect 39948 35566 40000 35572
rect 39856 35148 39908 35154
rect 39856 35090 39908 35096
rect 39868 34746 39896 35090
rect 39856 34740 39908 34746
rect 39856 34682 39908 34688
rect 39856 34060 39908 34066
rect 39960 34048 39988 35566
rect 39908 34020 39988 34048
rect 39856 34002 39908 34008
rect 39868 33522 39896 34002
rect 40052 33658 40080 36518
rect 40604 36378 40632 36586
rect 40592 36372 40644 36378
rect 40592 36314 40644 36320
rect 40408 35556 40460 35562
rect 40408 35498 40460 35504
rect 40420 34610 40448 35498
rect 40696 35222 40724 36654
rect 40880 36310 40908 38150
rect 41064 37738 41092 38150
rect 41052 37732 41104 37738
rect 41052 37674 41104 37680
rect 41052 37188 41104 37194
rect 41052 37130 41104 37136
rect 41064 36854 41092 37130
rect 41144 36916 41196 36922
rect 41144 36858 41196 36864
rect 41052 36848 41104 36854
rect 41052 36790 41104 36796
rect 41064 36650 41092 36790
rect 41052 36644 41104 36650
rect 41052 36586 41104 36592
rect 41156 36310 41184 36858
rect 40868 36304 40920 36310
rect 40868 36246 40920 36252
rect 41144 36304 41196 36310
rect 41144 36246 41196 36252
rect 40880 35834 40908 36246
rect 41156 35834 41184 36246
rect 40868 35828 40920 35834
rect 40868 35770 40920 35776
rect 41144 35828 41196 35834
rect 41144 35770 41196 35776
rect 40868 35488 40920 35494
rect 40868 35430 40920 35436
rect 40684 35216 40736 35222
rect 40684 35158 40736 35164
rect 40696 34746 40724 35158
rect 40684 34740 40736 34746
rect 40684 34682 40736 34688
rect 40408 34604 40460 34610
rect 40408 34546 40460 34552
rect 40696 34474 40724 34682
rect 40684 34468 40736 34474
rect 40684 34410 40736 34416
rect 40696 34134 40724 34410
rect 40880 34134 40908 35430
rect 40408 34128 40460 34134
rect 40408 34070 40460 34076
rect 40684 34128 40736 34134
rect 40684 34070 40736 34076
rect 40868 34128 40920 34134
rect 40868 34070 40920 34076
rect 40040 33652 40092 33658
rect 40040 33594 40092 33600
rect 39856 33516 39908 33522
rect 39856 33458 39908 33464
rect 40052 33454 40080 33594
rect 40040 33448 40092 33454
rect 40040 33390 40092 33396
rect 39684 33106 39804 33134
rect 39776 32978 39804 33106
rect 39764 32972 39816 32978
rect 39764 32914 39816 32920
rect 39776 32230 39804 32914
rect 39764 32224 39816 32230
rect 39764 32166 39816 32172
rect 39764 31816 39816 31822
rect 39764 31758 39816 31764
rect 39776 31346 39804 31758
rect 39764 31340 39816 31346
rect 39764 31282 39816 31288
rect 39396 30932 39448 30938
rect 39396 30874 39448 30880
rect 39396 30796 39448 30802
rect 39580 30796 39632 30802
rect 39448 30756 39528 30784
rect 39396 30738 39448 30744
rect 39304 30252 39356 30258
rect 39304 30194 39356 30200
rect 39316 29850 39344 30194
rect 39500 30054 39528 30756
rect 39580 30738 39632 30744
rect 39592 30190 39620 30738
rect 39672 30728 39724 30734
rect 39672 30670 39724 30676
rect 39580 30184 39632 30190
rect 39580 30126 39632 30132
rect 39488 30048 39540 30054
rect 39488 29990 39540 29996
rect 39304 29844 39356 29850
rect 39304 29786 39356 29792
rect 39396 28960 39448 28966
rect 39396 28902 39448 28908
rect 39304 28620 39356 28626
rect 39304 28562 39356 28568
rect 39316 28218 39344 28562
rect 39304 28212 39356 28218
rect 39304 28154 39356 28160
rect 39408 28014 39436 28902
rect 39500 28150 39528 29990
rect 39592 29510 39620 30126
rect 39684 29850 39712 30670
rect 39764 30184 39816 30190
rect 39764 30126 39816 30132
rect 39672 29844 39724 29850
rect 39672 29786 39724 29792
rect 39580 29504 39632 29510
rect 39580 29446 39632 29452
rect 39592 29170 39620 29446
rect 39580 29164 39632 29170
rect 39580 29106 39632 29112
rect 39592 28626 39620 29106
rect 39776 28694 39804 30126
rect 39764 28688 39816 28694
rect 39764 28630 39816 28636
rect 39580 28620 39632 28626
rect 39580 28562 39632 28568
rect 39592 28218 39620 28562
rect 39580 28212 39632 28218
rect 39580 28154 39632 28160
rect 39488 28144 39540 28150
rect 39488 28086 39540 28092
rect 39396 28008 39448 28014
rect 39396 27950 39448 27956
rect 40052 27878 40080 33390
rect 40316 32904 40368 32910
rect 40316 32846 40368 32852
rect 40328 32570 40356 32846
rect 40316 32564 40368 32570
rect 40316 32506 40368 32512
rect 40420 31958 40448 34070
rect 40500 33856 40552 33862
rect 40500 33798 40552 33804
rect 40512 31958 40540 33798
rect 40880 33658 40908 34070
rect 40868 33652 40920 33658
rect 40868 33594 40920 33600
rect 41248 33590 41276 38830
rect 42352 38758 42380 39460
rect 41972 38752 42024 38758
rect 41972 38694 42024 38700
rect 42340 38752 42392 38758
rect 42340 38694 42392 38700
rect 41788 38480 41840 38486
rect 41788 38422 41840 38428
rect 41880 38480 41932 38486
rect 41880 38422 41932 38428
rect 41512 37732 41564 37738
rect 41512 37674 41564 37680
rect 41524 36854 41552 37674
rect 41800 37466 41828 38422
rect 41892 37670 41920 38422
rect 41880 37664 41932 37670
rect 41880 37606 41932 37612
rect 41788 37460 41840 37466
rect 41788 37402 41840 37408
rect 41512 36848 41564 36854
rect 41512 36790 41564 36796
rect 41524 36174 41552 36790
rect 41512 36168 41564 36174
rect 41512 36110 41564 36116
rect 41524 35698 41552 36110
rect 41512 35692 41564 35698
rect 41512 35634 41564 35640
rect 41420 34128 41472 34134
rect 41420 34070 41472 34076
rect 41432 33590 41460 34070
rect 41524 33998 41552 35634
rect 41788 35556 41840 35562
rect 41788 35498 41840 35504
rect 41800 35018 41828 35498
rect 41788 35012 41840 35018
rect 41788 34954 41840 34960
rect 41512 33992 41564 33998
rect 41512 33934 41564 33940
rect 41236 33584 41288 33590
rect 41236 33526 41288 33532
rect 41420 33584 41472 33590
rect 41420 33526 41472 33532
rect 40592 33380 40644 33386
rect 40592 33322 40644 33328
rect 40408 31952 40460 31958
rect 40408 31894 40460 31900
rect 40500 31952 40552 31958
rect 40500 31894 40552 31900
rect 40604 31346 40632 33322
rect 40960 33312 41012 33318
rect 40960 33254 41012 33260
rect 40972 32434 41000 33254
rect 41052 33040 41104 33046
rect 41052 32982 41104 32988
rect 41064 32570 41092 32982
rect 41880 32904 41932 32910
rect 41880 32846 41932 32852
rect 41052 32564 41104 32570
rect 41052 32506 41104 32512
rect 40960 32428 41012 32434
rect 40960 32370 41012 32376
rect 41064 32280 41092 32506
rect 41788 32360 41840 32366
rect 41788 32302 41840 32308
rect 41144 32292 41196 32298
rect 41064 32252 41144 32280
rect 41064 32026 41092 32252
rect 41144 32234 41196 32240
rect 41052 32020 41104 32026
rect 41052 31962 41104 31968
rect 41064 31482 41092 31962
rect 41604 31952 41656 31958
rect 41604 31894 41656 31900
rect 41696 31952 41748 31958
rect 41696 31894 41748 31900
rect 41052 31476 41104 31482
rect 41052 31418 41104 31424
rect 40592 31340 40644 31346
rect 40592 31282 40644 31288
rect 41064 31142 41092 31418
rect 41144 31340 41196 31346
rect 41144 31282 41196 31288
rect 41052 31136 41104 31142
rect 41052 31078 41104 31084
rect 40314 30968 40370 30977
rect 41156 30938 41184 31282
rect 41616 30938 41644 31894
rect 41708 31754 41736 31894
rect 41696 31748 41748 31754
rect 41696 31690 41748 31696
rect 41708 31482 41736 31690
rect 41696 31476 41748 31482
rect 41696 31418 41748 31424
rect 40314 30903 40370 30912
rect 40592 30932 40644 30938
rect 40224 30048 40276 30054
rect 40224 29990 40276 29996
rect 40132 29708 40184 29714
rect 40132 29650 40184 29656
rect 40144 29238 40172 29650
rect 40132 29232 40184 29238
rect 40132 29174 40184 29180
rect 40236 28966 40264 29990
rect 40328 29578 40356 30903
rect 40592 30874 40644 30880
rect 41144 30932 41196 30938
rect 41144 30874 41196 30880
rect 41604 30932 41656 30938
rect 41604 30874 41656 30880
rect 40500 30592 40552 30598
rect 40500 30534 40552 30540
rect 40512 30190 40540 30534
rect 40500 30184 40552 30190
rect 40500 30126 40552 30132
rect 40500 29844 40552 29850
rect 40500 29786 40552 29792
rect 40316 29572 40368 29578
rect 40316 29514 40368 29520
rect 40512 29170 40540 29786
rect 40500 29164 40552 29170
rect 40500 29106 40552 29112
rect 40224 28960 40276 28966
rect 40224 28902 40276 28908
rect 40236 28762 40264 28902
rect 40224 28756 40276 28762
rect 40224 28698 40276 28704
rect 40604 28626 40632 30874
rect 41512 30864 41564 30870
rect 41512 30806 41564 30812
rect 41524 30258 41552 30806
rect 41512 30252 41564 30258
rect 41512 30194 41564 30200
rect 40684 30116 40736 30122
rect 40684 30058 40736 30064
rect 40696 29714 40724 30058
rect 41420 30048 41472 30054
rect 41420 29990 41472 29996
rect 40684 29708 40736 29714
rect 40684 29650 40736 29656
rect 41432 28694 41460 29990
rect 41512 29708 41564 29714
rect 41512 29650 41564 29656
rect 41524 28762 41552 29650
rect 41512 28756 41564 28762
rect 41512 28698 41564 28704
rect 41420 28688 41472 28694
rect 41420 28630 41472 28636
rect 40592 28620 40644 28626
rect 40592 28562 40644 28568
rect 40604 28218 40632 28562
rect 41800 28558 41828 32302
rect 41892 31822 41920 32846
rect 41880 31816 41932 31822
rect 41880 31758 41932 31764
rect 41892 30734 41920 31758
rect 41880 30728 41932 30734
rect 41880 30670 41932 30676
rect 41892 30394 41920 30670
rect 41880 30388 41932 30394
rect 41880 30330 41932 30336
rect 41788 28552 41840 28558
rect 41788 28494 41840 28500
rect 40960 28416 41012 28422
rect 40960 28358 41012 28364
rect 41144 28416 41196 28422
rect 41144 28358 41196 28364
rect 40224 28212 40276 28218
rect 40224 28154 40276 28160
rect 40592 28212 40644 28218
rect 40592 28154 40644 28160
rect 40040 27872 40092 27878
rect 40040 27814 40092 27820
rect 39488 27668 39540 27674
rect 39488 27610 39540 27616
rect 39396 27328 39448 27334
rect 39396 27270 39448 27276
rect 39408 26450 39436 27270
rect 39500 26858 39528 27610
rect 39580 27464 39632 27470
rect 39580 27406 39632 27412
rect 39488 26852 39540 26858
rect 39488 26794 39540 26800
rect 39396 26444 39448 26450
rect 39396 26386 39448 26392
rect 39212 26376 39264 26382
rect 39212 26318 39264 26324
rect 39224 24886 39252 26318
rect 39408 26042 39436 26386
rect 39396 26036 39448 26042
rect 39396 25978 39448 25984
rect 39408 25362 39436 25978
rect 39304 25356 39356 25362
rect 39304 25298 39356 25304
rect 39396 25356 39448 25362
rect 39396 25298 39448 25304
rect 39316 24954 39344 25298
rect 39408 24954 39436 25298
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 39396 24948 39448 24954
rect 39396 24890 39448 24896
rect 39212 24880 39264 24886
rect 39212 24822 39264 24828
rect 39224 22098 39252 24822
rect 39408 24274 39436 24890
rect 39500 24342 39528 26794
rect 39592 26790 39620 27406
rect 39672 26920 39724 26926
rect 39672 26862 39724 26868
rect 39580 26784 39632 26790
rect 39580 26726 39632 26732
rect 39592 25906 39620 26726
rect 39684 26518 39712 26862
rect 39672 26512 39724 26518
rect 39672 26454 39724 26460
rect 39580 25900 39632 25906
rect 39580 25842 39632 25848
rect 39948 25288 40000 25294
rect 39948 25230 40000 25236
rect 39488 24336 39540 24342
rect 39488 24278 39540 24284
rect 39396 24268 39448 24274
rect 39396 24210 39448 24216
rect 39408 23662 39436 24210
rect 39488 24200 39540 24206
rect 39488 24142 39540 24148
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 39408 23186 39436 23598
rect 39500 23322 39528 24142
rect 39960 23730 39988 25230
rect 40052 23798 40080 27814
rect 40132 27328 40184 27334
rect 40132 27270 40184 27276
rect 40144 25770 40172 27270
rect 40132 25764 40184 25770
rect 40132 25706 40184 25712
rect 40040 23792 40092 23798
rect 40040 23734 40092 23740
rect 39948 23724 40000 23730
rect 39948 23666 40000 23672
rect 39488 23316 39540 23322
rect 39488 23258 39540 23264
rect 39304 23180 39356 23186
rect 39304 23122 39356 23128
rect 39396 23180 39448 23186
rect 39396 23122 39448 23128
rect 39316 22438 39344 23122
rect 40052 22778 40080 23734
rect 40236 23050 40264 28154
rect 40972 27606 41000 28358
rect 41156 27946 41184 28358
rect 41800 28132 41828 28494
rect 41880 28144 41932 28150
rect 41800 28104 41880 28132
rect 41880 28086 41932 28092
rect 41984 28098 42012 38694
rect 42352 36786 42380 38694
rect 42432 37732 42484 37738
rect 42432 37674 42484 37680
rect 42444 37466 42472 37674
rect 42432 37460 42484 37466
rect 42432 37402 42484 37408
rect 42444 36922 42472 37402
rect 42432 36916 42484 36922
rect 42432 36858 42484 36864
rect 42340 36780 42392 36786
rect 42340 36722 42392 36728
rect 42536 36718 42564 40967
rect 42628 40662 42656 41142
rect 42616 40656 42668 40662
rect 42616 40598 42668 40604
rect 42720 39522 42748 43658
rect 43548 43330 43576 44832
rect 43720 44814 43772 44820
rect 43824 44402 43852 44950
rect 43812 44396 43864 44402
rect 43812 44338 43864 44344
rect 43720 44328 43772 44334
rect 43720 44270 43772 44276
rect 43628 44192 43680 44198
rect 43628 44134 43680 44140
rect 43640 43790 43668 44134
rect 43732 43790 43760 44270
rect 43824 43926 43852 44338
rect 44272 44328 44324 44334
rect 44836 44305 44864 45222
rect 44914 44840 44970 44849
rect 44914 44775 44970 44784
rect 44272 44270 44324 44276
rect 44822 44296 44878 44305
rect 43812 43920 43864 43926
rect 43812 43862 43864 43868
rect 44088 43920 44140 43926
rect 44088 43862 44140 43868
rect 43628 43784 43680 43790
rect 43628 43726 43680 43732
rect 43720 43784 43772 43790
rect 43772 43744 43852 43772
rect 43720 43726 43772 43732
rect 43640 43450 43668 43726
rect 43628 43444 43680 43450
rect 43628 43386 43680 43392
rect 43548 43302 43760 43330
rect 43536 43104 43588 43110
rect 43456 43064 43536 43092
rect 43456 42702 43484 43064
rect 43536 43046 43588 43052
rect 43536 42832 43588 42838
rect 43536 42774 43588 42780
rect 43444 42696 43496 42702
rect 43444 42638 43496 42644
rect 43076 42288 43128 42294
rect 43076 42230 43128 42236
rect 43088 41274 43116 42230
rect 43456 42226 43484 42638
rect 43548 42362 43576 42774
rect 43536 42356 43588 42362
rect 43536 42298 43588 42304
rect 43732 42294 43760 43302
rect 43824 42294 43852 43744
rect 44100 43450 44128 43862
rect 44088 43444 44140 43450
rect 44088 43386 44140 43392
rect 43996 43172 44048 43178
rect 44048 43132 44128 43160
rect 43996 43114 44048 43120
rect 43720 42288 43772 42294
rect 43720 42230 43772 42236
rect 43812 42288 43864 42294
rect 43812 42230 43864 42236
rect 43444 42220 43496 42226
rect 43444 42162 43496 42168
rect 43904 42084 43956 42090
rect 43904 42026 43956 42032
rect 43996 42084 44048 42090
rect 43996 42026 44048 42032
rect 43916 41818 43944 42026
rect 43904 41812 43956 41818
rect 43904 41754 43956 41760
rect 43352 41676 43404 41682
rect 43352 41618 43404 41624
rect 43076 41268 43128 41274
rect 43076 41210 43128 41216
rect 42800 40384 42852 40390
rect 42800 40326 42852 40332
rect 42812 40050 42840 40326
rect 43088 40050 43116 41210
rect 43364 41138 43392 41618
rect 44008 41614 44036 42026
rect 43996 41608 44048 41614
rect 43996 41550 44048 41556
rect 43352 41132 43404 41138
rect 43352 41074 43404 41080
rect 43364 41041 43392 41074
rect 43350 41032 43406 41041
rect 43350 40967 43406 40976
rect 43812 40588 43864 40594
rect 43812 40530 43864 40536
rect 42800 40044 42852 40050
rect 42800 39986 42852 39992
rect 43076 40044 43128 40050
rect 43076 39986 43128 39992
rect 42812 39642 42840 39986
rect 43824 39846 43852 40530
rect 43352 39840 43404 39846
rect 43352 39782 43404 39788
rect 43812 39840 43864 39846
rect 43812 39782 43864 39788
rect 42800 39636 42852 39642
rect 42800 39578 42852 39584
rect 43364 39556 43392 39782
rect 43444 39568 43496 39574
rect 43364 39528 43444 39556
rect 42628 39494 42748 39522
rect 43444 39510 43496 39516
rect 42524 36712 42576 36718
rect 42524 36654 42576 36660
rect 42628 35630 42656 39494
rect 42708 39432 42760 39438
rect 42708 39374 42760 39380
rect 42720 39098 42748 39374
rect 43456 39098 43484 39510
rect 42708 39092 42760 39098
rect 42708 39034 42760 39040
rect 43444 39092 43496 39098
rect 43444 39034 43496 39040
rect 43824 38729 43852 39782
rect 43810 38720 43866 38729
rect 43810 38655 43866 38664
rect 43628 38276 43680 38282
rect 43628 38218 43680 38224
rect 42616 35624 42668 35630
rect 42616 35566 42668 35572
rect 43260 35624 43312 35630
rect 43260 35566 43312 35572
rect 42800 35556 42852 35562
rect 42800 35498 42852 35504
rect 42812 35018 42840 35498
rect 43168 35080 43220 35086
rect 43168 35022 43220 35028
rect 42800 35012 42852 35018
rect 42800 34954 42852 34960
rect 42812 34610 42840 34954
rect 42800 34604 42852 34610
rect 42800 34546 42852 34552
rect 42524 34468 42576 34474
rect 42524 34410 42576 34416
rect 42536 34202 42564 34410
rect 42524 34196 42576 34202
rect 42524 34138 42576 34144
rect 43180 34134 43208 35022
rect 43168 34128 43220 34134
rect 43168 34070 43220 34076
rect 43180 33930 43208 34070
rect 43168 33924 43220 33930
rect 43168 33866 43220 33872
rect 42984 33448 43036 33454
rect 42984 33390 43036 33396
rect 42156 33312 42208 33318
rect 42156 33254 42208 33260
rect 42168 32434 42196 33254
rect 42156 32428 42208 32434
rect 42156 32370 42208 32376
rect 42892 32428 42944 32434
rect 42892 32370 42944 32376
rect 42904 32298 42932 32370
rect 42892 32292 42944 32298
rect 42892 32234 42944 32240
rect 42616 32224 42668 32230
rect 42616 32166 42668 32172
rect 42628 31958 42656 32166
rect 42904 32026 42932 32234
rect 42892 32020 42944 32026
rect 42892 31962 42944 31968
rect 42616 31952 42668 31958
rect 42616 31894 42668 31900
rect 42628 31414 42656 31894
rect 42616 31408 42668 31414
rect 42616 31350 42668 31356
rect 42064 31204 42116 31210
rect 42064 31146 42116 31152
rect 42076 31113 42104 31146
rect 42062 31104 42118 31113
rect 42062 31039 42118 31048
rect 42076 29152 42104 31039
rect 42800 30252 42852 30258
rect 42800 30194 42852 30200
rect 42432 30048 42484 30054
rect 42432 29990 42484 29996
rect 42444 29850 42472 29990
rect 42432 29844 42484 29850
rect 42432 29786 42484 29792
rect 42524 29776 42576 29782
rect 42524 29718 42576 29724
rect 42536 29238 42564 29718
rect 42812 29714 42840 30194
rect 42800 29708 42852 29714
rect 42800 29650 42852 29656
rect 42524 29232 42576 29238
rect 42524 29174 42576 29180
rect 42156 29164 42208 29170
rect 42076 29124 42156 29152
rect 42156 29106 42208 29112
rect 42340 29164 42392 29170
rect 42340 29106 42392 29112
rect 42352 28762 42380 29106
rect 42536 28966 42564 29174
rect 42996 28994 43024 33390
rect 43168 33312 43220 33318
rect 43168 33254 43220 33260
rect 43180 31822 43208 33254
rect 43168 31816 43220 31822
rect 43168 31758 43220 31764
rect 43180 31482 43208 31758
rect 43168 31476 43220 31482
rect 43168 31418 43220 31424
rect 43076 31204 43128 31210
rect 43076 31146 43128 31152
rect 43088 30938 43116 31146
rect 43076 30932 43128 30938
rect 43076 30874 43128 30880
rect 43272 30802 43300 35566
rect 43444 35488 43496 35494
rect 43444 35430 43496 35436
rect 43456 34610 43484 35430
rect 43536 35216 43588 35222
rect 43536 35158 43588 35164
rect 43548 34746 43576 35158
rect 43640 35086 43668 38218
rect 43720 36236 43772 36242
rect 43824 36224 43852 38655
rect 43996 38344 44048 38350
rect 43996 38286 44048 38292
rect 43904 38004 43956 38010
rect 43904 37946 43956 37952
rect 43916 37126 43944 37946
rect 44008 37670 44036 38286
rect 44100 38010 44128 43132
rect 44180 42288 44232 42294
rect 44180 42230 44232 42236
rect 44192 40186 44220 42230
rect 44180 40180 44232 40186
rect 44180 40122 44232 40128
rect 44192 39574 44220 40122
rect 44180 39568 44232 39574
rect 44180 39510 44232 39516
rect 44284 38894 44312 44270
rect 44822 44231 44878 44240
rect 44272 38888 44324 38894
rect 44272 38830 44324 38836
rect 44180 38752 44232 38758
rect 44180 38694 44232 38700
rect 44456 38752 44508 38758
rect 44456 38694 44508 38700
rect 44088 38004 44140 38010
rect 44088 37946 44140 37952
rect 44192 37874 44220 38694
rect 44272 38480 44324 38486
rect 44272 38422 44324 38428
rect 44180 37868 44232 37874
rect 44180 37810 44232 37816
rect 44284 37738 44312 38422
rect 44272 37732 44324 37738
rect 44272 37674 44324 37680
rect 43996 37664 44048 37670
rect 43996 37606 44048 37612
rect 44008 37466 44036 37606
rect 43996 37460 44048 37466
rect 43996 37402 44048 37408
rect 44284 37194 44312 37674
rect 44364 37256 44416 37262
rect 44364 37198 44416 37204
rect 44272 37188 44324 37194
rect 44272 37130 44324 37136
rect 43904 37120 43956 37126
rect 43904 37062 43956 37068
rect 44284 36650 44312 37130
rect 44376 36922 44404 37198
rect 44364 36916 44416 36922
rect 44364 36858 44416 36864
rect 44272 36644 44324 36650
rect 44272 36586 44324 36592
rect 43904 36576 43956 36582
rect 43904 36518 43956 36524
rect 43772 36196 43852 36224
rect 43720 36178 43772 36184
rect 43732 35494 43760 36178
rect 43720 35488 43772 35494
rect 43720 35430 43772 35436
rect 43628 35080 43680 35086
rect 43628 35022 43680 35028
rect 43536 34740 43588 34746
rect 43536 34682 43588 34688
rect 43444 34604 43496 34610
rect 43444 34546 43496 34552
rect 43628 33856 43680 33862
rect 43628 33798 43680 33804
rect 43640 33386 43668 33798
rect 43628 33380 43680 33386
rect 43628 33322 43680 33328
rect 43260 30796 43312 30802
rect 43260 30738 43312 30744
rect 43076 30728 43128 30734
rect 43076 30670 43128 30676
rect 43088 30258 43116 30670
rect 43272 30394 43300 30738
rect 43260 30388 43312 30394
rect 43260 30330 43312 30336
rect 43076 30252 43128 30258
rect 43076 30194 43128 30200
rect 43088 29170 43116 30194
rect 43076 29164 43128 29170
rect 43076 29106 43128 29112
rect 42904 28966 43024 28994
rect 42524 28960 42576 28966
rect 42524 28902 42576 28908
rect 42340 28756 42392 28762
rect 42340 28698 42392 28704
rect 42064 28688 42116 28694
rect 42064 28630 42116 28636
rect 42076 28218 42104 28630
rect 42064 28212 42116 28218
rect 42064 28154 42116 28160
rect 41984 28070 42196 28098
rect 41144 27940 41196 27946
rect 41144 27882 41196 27888
rect 41236 27940 41288 27946
rect 41236 27882 41288 27888
rect 42064 27940 42116 27946
rect 42064 27882 42116 27888
rect 40960 27600 41012 27606
rect 40960 27542 41012 27548
rect 40500 27328 40552 27334
rect 40500 27270 40552 27276
rect 40512 26926 40540 27270
rect 40500 26920 40552 26926
rect 40500 26862 40552 26868
rect 41156 26586 41184 27882
rect 41248 27674 41276 27882
rect 41236 27668 41288 27674
rect 41236 27610 41288 27616
rect 41788 27600 41840 27606
rect 41788 27542 41840 27548
rect 41972 27600 42024 27606
rect 41972 27542 42024 27548
rect 41800 27130 41828 27542
rect 41788 27124 41840 27130
rect 41788 27066 41840 27072
rect 41984 26790 42012 27542
rect 41972 26784 42024 26790
rect 41972 26726 42024 26732
rect 41144 26580 41196 26586
rect 41144 26522 41196 26528
rect 41984 26518 42012 26726
rect 41972 26512 42024 26518
rect 41972 26454 42024 26460
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 40696 26042 40724 26318
rect 41052 26240 41104 26246
rect 41052 26182 41104 26188
rect 40684 26036 40736 26042
rect 40684 25978 40736 25984
rect 41064 25906 41092 26182
rect 41984 26042 42012 26454
rect 41972 26036 42024 26042
rect 41972 25978 42024 25984
rect 42076 25906 42104 27882
rect 41052 25900 41104 25906
rect 41052 25842 41104 25848
rect 41696 25900 41748 25906
rect 41696 25842 41748 25848
rect 42064 25900 42116 25906
rect 42064 25842 42116 25848
rect 41052 25764 41104 25770
rect 41052 25706 41104 25712
rect 41064 25498 41092 25706
rect 41052 25492 41104 25498
rect 41052 25434 41104 25440
rect 41708 25294 41736 25842
rect 41788 25424 41840 25430
rect 41788 25366 41840 25372
rect 41696 25288 41748 25294
rect 41696 25230 41748 25236
rect 40960 24676 41012 24682
rect 40880 24636 40960 24664
rect 40316 24336 40368 24342
rect 40316 24278 40368 24284
rect 40328 23526 40356 24278
rect 40880 24070 40908 24636
rect 40960 24618 41012 24624
rect 41800 24614 41828 25366
rect 41972 25288 42024 25294
rect 41972 25230 42024 25236
rect 41984 24818 42012 25230
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 41788 24608 41840 24614
rect 41788 24550 41840 24556
rect 42064 24608 42116 24614
rect 42064 24550 42116 24556
rect 41800 24410 41828 24550
rect 41788 24404 41840 24410
rect 41788 24346 41840 24352
rect 42076 24342 42104 24550
rect 42064 24336 42116 24342
rect 42064 24278 42116 24284
rect 41236 24200 41288 24206
rect 41236 24142 41288 24148
rect 40868 24064 40920 24070
rect 40868 24006 40920 24012
rect 40880 23798 40908 24006
rect 41248 23866 41276 24142
rect 41236 23860 41288 23866
rect 41236 23802 41288 23808
rect 40868 23792 40920 23798
rect 40868 23734 40920 23740
rect 40684 23724 40736 23730
rect 40684 23666 40736 23672
rect 40316 23520 40368 23526
rect 40316 23462 40368 23468
rect 40224 23044 40276 23050
rect 40224 22986 40276 22992
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40236 22574 40264 22986
rect 40224 22568 40276 22574
rect 40224 22510 40276 22516
rect 39672 22500 39724 22506
rect 39592 22460 39672 22488
rect 39304 22432 39356 22438
rect 39304 22374 39356 22380
rect 39212 22092 39264 22098
rect 39212 22034 39264 22040
rect 39028 21004 39080 21010
rect 39028 20946 39080 20952
rect 38936 20800 38988 20806
rect 38936 20742 38988 20748
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38856 20398 38884 20538
rect 38948 20398 38976 20742
rect 39040 20602 39068 20946
rect 39028 20596 39080 20602
rect 39028 20538 39080 20544
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38936 20392 38988 20398
rect 38936 20334 38988 20340
rect 38948 20058 38976 20334
rect 38936 20052 38988 20058
rect 38936 19994 38988 20000
rect 38384 19780 38436 19786
rect 38384 19722 38436 19728
rect 38396 19514 38424 19722
rect 38948 19514 38976 19994
rect 39316 19922 39344 22374
rect 39304 19916 39356 19922
rect 39304 19858 39356 19864
rect 38384 19508 38436 19514
rect 38384 19450 38436 19456
rect 38936 19508 38988 19514
rect 38936 19450 38988 19456
rect 38948 18426 38976 19450
rect 39316 19446 39344 19858
rect 39304 19440 39356 19446
rect 39304 19382 39356 19388
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 38948 18222 38976 18362
rect 39212 18284 39264 18290
rect 39212 18226 39264 18232
rect 38936 18216 38988 18222
rect 38936 18158 38988 18164
rect 38292 18080 38344 18086
rect 38292 18022 38344 18028
rect 38304 17338 38332 18022
rect 38660 17808 38712 17814
rect 38660 17750 38712 17756
rect 38672 17338 38700 17750
rect 38292 17332 38344 17338
rect 38292 17274 38344 17280
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 38304 17134 38332 17274
rect 38292 17128 38344 17134
rect 38292 17070 38344 17076
rect 38016 16720 38068 16726
rect 38016 16662 38068 16668
rect 37832 16584 37884 16590
rect 37832 16526 37884 16532
rect 36912 16040 36964 16046
rect 36912 15982 36964 15988
rect 36924 15706 36952 15982
rect 37844 15978 37872 16526
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37832 15972 37884 15978
rect 37832 15914 37884 15920
rect 37844 15706 37872 15914
rect 37936 15706 37964 15982
rect 38028 15910 38056 16662
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 36912 15700 36964 15706
rect 36912 15642 36964 15648
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 36544 15496 36596 15502
rect 36544 15438 36596 15444
rect 36556 15162 36584 15438
rect 36820 15360 36872 15366
rect 36820 15302 36872 15308
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36832 14822 36860 15302
rect 36912 14952 36964 14958
rect 36912 14894 36964 14900
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 36820 14816 36872 14822
rect 36820 14758 36872 14764
rect 36452 14612 36504 14618
rect 36452 14554 36504 14560
rect 35624 14476 35676 14482
rect 35624 14418 35676 14424
rect 36268 14476 36320 14482
rect 36268 14418 36320 14424
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 35440 14000 35492 14006
rect 35440 13942 35492 13948
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34796 12708 34848 12714
rect 34796 12650 34848 12656
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34808 12306 34836 12650
rect 35360 12442 35388 12786
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 34440 9518 34468 12174
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35544 11694 35572 12038
rect 35532 11688 35584 11694
rect 35820 11665 35848 14214
rect 36280 14074 36308 14418
rect 36360 14272 36412 14278
rect 36360 14214 36412 14220
rect 36268 14068 36320 14074
rect 36268 14010 36320 14016
rect 36372 13841 36400 14214
rect 36358 13832 36414 13841
rect 36358 13767 36414 13776
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 36004 12918 36032 13330
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 35992 12912 36044 12918
rect 35992 12854 36044 12860
rect 36188 12782 36216 13262
rect 36176 12776 36228 12782
rect 36176 12718 36228 12724
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 36096 12306 36124 12378
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 36096 11898 36124 12242
rect 36084 11892 36136 11898
rect 36084 11834 36136 11840
rect 35532 11630 35584 11636
rect 35806 11656 35862 11665
rect 35544 11218 35572 11630
rect 35716 11620 35768 11626
rect 35806 11591 35862 11600
rect 35716 11562 35768 11568
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 35532 11212 35584 11218
rect 35532 11154 35584 11160
rect 34624 10674 34652 11154
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 34624 10577 34652 10610
rect 34610 10568 34666 10577
rect 34610 10503 34666 10512
rect 35544 10470 35572 11154
rect 35728 10674 35756 11562
rect 35716 10668 35768 10674
rect 35716 10610 35768 10616
rect 35716 10532 35768 10538
rect 35716 10474 35768 10480
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35544 10130 35572 10406
rect 35532 10124 35584 10130
rect 35532 10066 35584 10072
rect 35256 9988 35308 9994
rect 35256 9930 35308 9936
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35268 9654 35296 9930
rect 35544 9722 35572 10066
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35532 9716 35584 9722
rect 35532 9658 35584 9664
rect 35256 9648 35308 9654
rect 35256 9590 35308 9596
rect 34428 9512 34480 9518
rect 34428 9454 34480 9460
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 34440 8634 34468 8978
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34336 8424 34388 8430
rect 34336 8366 34388 8372
rect 33784 8016 33836 8022
rect 33784 7958 33836 7964
rect 33796 7546 33824 7958
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33336 6956 33456 6984
rect 33336 6322 33364 6956
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 33428 6662 33456 6802
rect 33416 6656 33468 6662
rect 33416 6598 33468 6604
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33428 6254 33456 6598
rect 33416 6248 33468 6254
rect 33416 6190 33468 6196
rect 33428 6118 33456 6190
rect 33968 6180 34020 6186
rect 33968 6122 34020 6128
rect 33416 6112 33468 6118
rect 33416 6054 33468 6060
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 32324 5370 32352 5714
rect 32312 5364 32364 5370
rect 32312 5306 32364 5312
rect 32692 4826 32720 5714
rect 33060 5098 33088 5782
rect 33428 5574 33456 6054
rect 33980 5778 34008 6122
rect 33968 5772 34020 5778
rect 33968 5714 34020 5720
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 33428 5234 33456 5510
rect 33980 5370 34008 5714
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33600 5228 33652 5234
rect 33600 5170 33652 5176
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 33060 4826 33088 5034
rect 33428 5030 33456 5170
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 32680 4820 32732 4826
rect 32680 4762 32732 4768
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 32588 4752 32640 4758
rect 32588 4694 32640 4700
rect 32128 4684 32180 4690
rect 32128 4626 32180 4632
rect 32140 4282 32168 4626
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 32048 4126 32168 4154
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 32048 3194 32076 3538
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 24858 54 25268 82
rect 32034 82 32090 480
rect 32140 82 32168 4126
rect 32600 3942 32628 4694
rect 32692 4622 32720 4762
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32772 4004 32824 4010
rect 32772 3946 32824 3952
rect 32588 3936 32640 3942
rect 32588 3878 32640 3884
rect 32784 3738 32812 3946
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 33428 3602 33456 4966
rect 33612 4622 33640 5170
rect 33692 5024 33744 5030
rect 33692 4966 33744 4972
rect 33704 4758 33732 4966
rect 33692 4752 33744 4758
rect 33692 4694 33744 4700
rect 33600 4616 33652 4622
rect 33600 4558 33652 4564
rect 33612 4282 33640 4558
rect 33600 4276 33652 4282
rect 33600 4218 33652 4224
rect 33704 4214 33732 4694
rect 33692 4208 33744 4214
rect 33692 4150 33744 4156
rect 34348 4154 34376 8366
rect 34808 7954 34836 8910
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34888 8424 34940 8430
rect 34888 8366 34940 8372
rect 34900 8090 34928 8366
rect 34888 8084 34940 8090
rect 34888 8026 34940 8032
rect 34796 7948 34848 7954
rect 34796 7890 34848 7896
rect 34808 6934 34836 7890
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35268 7154 35296 9590
rect 35544 9178 35572 9658
rect 35636 9586 35664 9998
rect 35728 9654 35756 10474
rect 35820 9994 35848 11591
rect 35900 11552 35952 11558
rect 35900 11494 35952 11500
rect 35808 9988 35860 9994
rect 35808 9930 35860 9936
rect 35912 9926 35940 11494
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 36096 10266 36124 10610
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 35900 9920 35952 9926
rect 35900 9862 35952 9868
rect 35716 9648 35768 9654
rect 35716 9590 35768 9596
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 35636 9178 35664 9522
rect 35728 9450 35756 9590
rect 35716 9444 35768 9450
rect 35716 9386 35768 9392
rect 35532 9172 35584 9178
rect 35532 9114 35584 9120
rect 35624 9172 35676 9178
rect 35624 9114 35676 9120
rect 35544 8430 35572 9114
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35544 7886 35572 8366
rect 35728 8022 35756 9386
rect 35716 8016 35768 8022
rect 35716 7958 35768 7964
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35440 7812 35492 7818
rect 35440 7754 35492 7760
rect 35176 7126 35296 7154
rect 34796 6928 34848 6934
rect 34796 6870 34848 6876
rect 35176 6866 35204 7126
rect 35256 6996 35308 7002
rect 35256 6938 35308 6944
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 34624 6458 34652 6802
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34612 6452 34664 6458
rect 34612 6394 34664 6400
rect 34624 5302 34652 6394
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34716 5234 34744 6734
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35268 6254 35296 6938
rect 35452 6934 35480 7754
rect 35728 7546 35756 7958
rect 35716 7540 35768 7546
rect 35716 7482 35768 7488
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 35440 6928 35492 6934
rect 35440 6870 35492 6876
rect 35256 6248 35308 6254
rect 35256 6190 35308 6196
rect 35452 5914 35480 6870
rect 35636 6458 35664 7346
rect 35716 7268 35768 7274
rect 35716 7210 35768 7216
rect 35624 6452 35676 6458
rect 35624 6394 35676 6400
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 34808 5098 34836 5850
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 34796 5092 34848 5098
rect 34796 5034 34848 5040
rect 35544 4826 35572 5170
rect 35532 4820 35584 4826
rect 35532 4762 35584 4768
rect 35728 4758 35756 7210
rect 35808 6928 35860 6934
rect 35808 6870 35860 6876
rect 35820 6118 35848 6870
rect 35808 6112 35860 6118
rect 35808 6054 35860 6060
rect 35716 4752 35768 4758
rect 35716 4694 35768 4700
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 33428 2990 33456 3538
rect 33704 3194 33732 4150
rect 34348 4126 34468 4154
rect 33692 3188 33744 3194
rect 33692 3130 33744 3136
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 34336 2984 34388 2990
rect 34336 2926 34388 2932
rect 33428 2514 33456 2926
rect 34348 2582 34376 2926
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 34440 2514 34468 4126
rect 34532 3641 34560 4422
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 35728 4214 35756 4694
rect 35716 4208 35768 4214
rect 35716 4150 35768 4156
rect 34612 3664 34664 3670
rect 34518 3632 34574 3641
rect 34612 3606 34664 3612
rect 34518 3567 34574 3576
rect 34624 3194 34652 3606
rect 35912 3602 35940 9862
rect 36372 9042 36400 13767
rect 36544 12708 36596 12714
rect 36544 12650 36596 12656
rect 36556 12306 36584 12650
rect 36544 12300 36596 12306
rect 36544 12242 36596 12248
rect 36452 12164 36504 12170
rect 36452 12106 36504 12112
rect 36464 10130 36492 12106
rect 36556 11898 36584 12242
rect 36636 12164 36688 12170
rect 36636 12106 36688 12112
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36648 10305 36676 12106
rect 36728 11688 36780 11694
rect 36728 11630 36780 11636
rect 36740 11354 36768 11630
rect 36728 11348 36780 11354
rect 36728 11290 36780 11296
rect 36634 10296 36690 10305
rect 36634 10231 36690 10240
rect 36452 10124 36504 10130
rect 36452 10066 36504 10072
rect 36464 9722 36492 10066
rect 36452 9716 36504 9722
rect 36452 9658 36504 9664
rect 36832 9217 36860 14758
rect 36924 14278 36952 14894
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 37188 13932 37240 13938
rect 37188 13874 37240 13880
rect 37004 13864 37056 13870
rect 37004 13806 37056 13812
rect 37016 13462 37044 13806
rect 37200 13734 37228 13874
rect 37188 13728 37240 13734
rect 37188 13670 37240 13676
rect 37004 13456 37056 13462
rect 37004 13398 37056 13404
rect 37292 13394 37320 14894
rect 37752 14822 37780 15506
rect 37832 14884 37884 14890
rect 37832 14826 37884 14832
rect 37740 14816 37792 14822
rect 37740 14758 37792 14764
rect 37844 14414 37872 14826
rect 38028 14550 38056 15846
rect 38292 15564 38344 15570
rect 38292 15506 38344 15512
rect 38304 15162 38332 15506
rect 38476 15428 38528 15434
rect 38476 15370 38528 15376
rect 38292 15156 38344 15162
rect 38292 15098 38344 15104
rect 38108 15088 38160 15094
rect 38108 15030 38160 15036
rect 38016 14544 38068 14550
rect 38016 14486 38068 14492
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37844 14074 37872 14350
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 38028 13938 38056 14486
rect 38016 13932 38068 13938
rect 38016 13874 38068 13880
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 37924 13388 37976 13394
rect 37924 13330 37976 13336
rect 37292 12986 37320 13330
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37292 12782 37320 12922
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 37292 12442 37320 12718
rect 37936 12714 37964 13330
rect 37556 12708 37608 12714
rect 37556 12650 37608 12656
rect 37924 12708 37976 12714
rect 37924 12650 37976 12656
rect 37280 12436 37332 12442
rect 37280 12378 37332 12384
rect 37280 11212 37332 11218
rect 37280 11154 37332 11160
rect 37292 10810 37320 11154
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 37004 10464 37056 10470
rect 37004 10406 37056 10412
rect 37016 9586 37044 10406
rect 37004 9580 37056 9586
rect 37004 9522 37056 9528
rect 36912 9376 36964 9382
rect 36912 9318 36964 9324
rect 36818 9208 36874 9217
rect 36818 9143 36874 9152
rect 36084 9036 36136 9042
rect 36084 8978 36136 8984
rect 36360 9036 36412 9042
rect 36360 8978 36412 8984
rect 36096 8294 36124 8978
rect 36084 8288 36136 8294
rect 36084 8230 36136 8236
rect 35992 7744 36044 7750
rect 35992 7686 36044 7692
rect 36004 7002 36032 7686
rect 35992 6996 36044 7002
rect 35992 6938 36044 6944
rect 36096 6390 36124 8230
rect 36372 8090 36400 8978
rect 36728 8968 36780 8974
rect 36728 8910 36780 8916
rect 36636 8424 36688 8430
rect 36636 8366 36688 8372
rect 36648 8294 36676 8366
rect 36636 8288 36688 8294
rect 36636 8230 36688 8236
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36740 7886 36768 8910
rect 36832 8430 36860 9143
rect 36820 8424 36872 8430
rect 36820 8366 36872 8372
rect 36832 8090 36860 8366
rect 36820 8084 36872 8090
rect 36820 8026 36872 8032
rect 36728 7880 36780 7886
rect 36924 7857 36952 9318
rect 37004 8288 37056 8294
rect 37004 8230 37056 8236
rect 36728 7822 36780 7828
rect 36910 7848 36966 7857
rect 36910 7783 36966 7792
rect 37016 7546 37044 8230
rect 37004 7540 37056 7546
rect 37004 7482 37056 7488
rect 36268 7268 36320 7274
rect 36268 7210 36320 7216
rect 36280 6905 36308 7210
rect 36266 6896 36322 6905
rect 36266 6831 36322 6840
rect 36280 6798 36308 6831
rect 36268 6792 36320 6798
rect 36268 6734 36320 6740
rect 36268 6656 36320 6662
rect 36188 6616 36268 6644
rect 36084 6384 36136 6390
rect 36084 6326 36136 6332
rect 36188 6186 36216 6616
rect 36268 6598 36320 6604
rect 36176 6180 36228 6186
rect 36176 6122 36228 6128
rect 36452 6180 36504 6186
rect 36452 6122 36504 6128
rect 36912 6180 36964 6186
rect 36912 6122 36964 6128
rect 36084 5024 36136 5030
rect 36084 4966 36136 4972
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 36004 3618 36032 4558
rect 36096 4078 36124 4966
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 36188 3913 36216 6122
rect 36360 5772 36412 5778
rect 36360 5714 36412 5720
rect 36372 5370 36400 5714
rect 36464 5370 36492 6122
rect 36820 5568 36872 5574
rect 36820 5510 36872 5516
rect 36360 5364 36412 5370
rect 36360 5306 36412 5312
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36832 4758 36860 5510
rect 36820 4752 36872 4758
rect 36820 4694 36872 4700
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36372 4010 36400 4150
rect 36924 4078 36952 6122
rect 37464 5704 37516 5710
rect 37464 5646 37516 5652
rect 37004 5568 37056 5574
rect 37004 5510 37056 5516
rect 37016 5234 37044 5510
rect 37096 5364 37148 5370
rect 37096 5306 37148 5312
rect 37004 5228 37056 5234
rect 37004 5170 37056 5176
rect 36912 4072 36964 4078
rect 36910 4040 36912 4049
rect 36964 4040 36966 4049
rect 36268 4004 36320 4010
rect 36268 3946 36320 3952
rect 36360 4004 36412 4010
rect 36910 3975 36966 3984
rect 36360 3946 36412 3952
rect 36924 3949 36952 3975
rect 36174 3904 36230 3913
rect 36174 3839 36230 3848
rect 36280 3738 36308 3946
rect 36268 3732 36320 3738
rect 36268 3674 36320 3680
rect 35900 3596 35952 3602
rect 36004 3590 36216 3618
rect 35900 3538 35952 3544
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 34624 2854 34652 3130
rect 34716 2990 34744 3334
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34704 2984 34756 2990
rect 34704 2926 34756 2932
rect 35072 2916 35124 2922
rect 35072 2858 35124 2864
rect 34612 2848 34664 2854
rect 34612 2790 34664 2796
rect 34624 2582 34652 2790
rect 34612 2576 34664 2582
rect 34612 2518 34664 2524
rect 35084 2514 35112 2858
rect 36004 2582 36032 3334
rect 36096 3126 36124 3470
rect 36188 3398 36216 3590
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36084 3120 36136 3126
rect 36084 3062 36136 3068
rect 36188 2650 36216 3334
rect 36556 3194 36584 3538
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 37016 2650 37044 5170
rect 37108 5098 37136 5306
rect 37096 5092 37148 5098
rect 37096 5034 37148 5040
rect 37476 4486 37504 5646
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 37476 4282 37504 4422
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37094 3768 37150 3777
rect 37094 3703 37150 3712
rect 37108 3670 37136 3703
rect 37568 3670 37596 12650
rect 38028 12646 38056 13874
rect 38120 12850 38148 15030
rect 38304 14958 38332 15098
rect 38488 14958 38516 15370
rect 38292 14952 38344 14958
rect 38292 14894 38344 14900
rect 38476 14952 38528 14958
rect 38476 14894 38528 14900
rect 38936 13728 38988 13734
rect 38936 13670 38988 13676
rect 38660 13320 38712 13326
rect 38660 13262 38712 13268
rect 38672 12850 38700 13262
rect 38108 12844 38160 12850
rect 38108 12786 38160 12792
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38844 12776 38896 12782
rect 38844 12718 38896 12724
rect 37648 12640 37700 12646
rect 37648 12582 37700 12588
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 37660 12102 37688 12582
rect 38028 12374 38056 12582
rect 38016 12368 38068 12374
rect 38016 12310 38068 12316
rect 37924 12232 37976 12238
rect 37924 12174 37976 12180
rect 37648 12096 37700 12102
rect 37648 12038 37700 12044
rect 37660 11762 37688 12038
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37660 11354 37688 11698
rect 37936 11626 37964 12174
rect 37924 11620 37976 11626
rect 37924 11562 37976 11568
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37648 11348 37700 11354
rect 37648 11290 37700 11296
rect 37844 11234 37872 11494
rect 37936 11354 37964 11562
rect 38028 11558 38056 12310
rect 38856 12170 38884 12718
rect 38844 12164 38896 12170
rect 38844 12106 38896 12112
rect 38016 11552 38068 11558
rect 38016 11494 38068 11500
rect 38568 11552 38620 11558
rect 38568 11494 38620 11500
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 37844 11206 37964 11234
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37740 11008 37792 11014
rect 37740 10950 37792 10956
rect 37752 9489 37780 10950
rect 37844 10674 37872 11086
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 10266 37872 10610
rect 37832 10260 37884 10266
rect 37832 10202 37884 10208
rect 37738 9480 37794 9489
rect 37738 9415 37794 9424
rect 37752 9382 37780 9415
rect 37740 9376 37792 9382
rect 37792 9336 37872 9364
rect 37740 9318 37792 9324
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37752 6390 37780 6802
rect 37740 6384 37792 6390
rect 37740 6326 37792 6332
rect 37648 5092 37700 5098
rect 37648 5034 37700 5040
rect 37740 5092 37792 5098
rect 37740 5034 37792 5040
rect 37660 4622 37688 5034
rect 37648 4616 37700 4622
rect 37648 4558 37700 4564
rect 37660 3777 37688 4558
rect 37646 3768 37702 3777
rect 37646 3703 37702 3712
rect 37096 3664 37148 3670
rect 37096 3606 37148 3612
rect 37556 3664 37608 3670
rect 37556 3606 37608 3612
rect 37568 2990 37596 3606
rect 37752 3097 37780 5034
rect 37844 3738 37872 9336
rect 37936 8945 37964 11206
rect 38028 10538 38056 11494
rect 38016 10532 38068 10538
rect 38016 10474 38068 10480
rect 38028 9178 38056 10474
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 37922 8936 37978 8945
rect 37922 8871 37978 8880
rect 37936 4554 37964 8871
rect 38028 8294 38056 9114
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8634 38148 8910
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 38016 8288 38068 8294
rect 38016 8230 38068 8236
rect 38028 7274 38056 8230
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 38488 7546 38516 7890
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38016 7268 38068 7274
rect 38016 7210 38068 7216
rect 38292 6656 38344 6662
rect 38292 6598 38344 6604
rect 38476 6656 38528 6662
rect 38580 6644 38608 11494
rect 38752 11280 38804 11286
rect 38752 11222 38804 11228
rect 38764 10606 38792 11222
rect 38752 10600 38804 10606
rect 38752 10542 38804 10548
rect 38752 10464 38804 10470
rect 38752 10406 38804 10412
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38672 9722 38700 9998
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 38764 9518 38792 10406
rect 38752 9512 38804 9518
rect 38752 9454 38804 9460
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38672 7342 38700 8774
rect 38752 8356 38804 8362
rect 38752 8298 38804 8304
rect 38764 8090 38792 8298
rect 38752 8084 38804 8090
rect 38752 8026 38804 8032
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 38528 6616 38608 6644
rect 38476 6598 38528 6604
rect 38304 6458 38332 6598
rect 38292 6452 38344 6458
rect 38292 6394 38344 6400
rect 38304 6254 38332 6394
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 38488 6236 38516 6598
rect 38568 6248 38620 6254
rect 38488 6208 38568 6236
rect 38016 5840 38068 5846
rect 38016 5782 38068 5788
rect 38028 5370 38056 5782
rect 38304 5370 38332 6190
rect 38016 5364 38068 5370
rect 38016 5306 38068 5312
rect 38292 5364 38344 5370
rect 38292 5306 38344 5312
rect 38304 5166 38332 5306
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38304 4690 38332 5102
rect 38488 4865 38516 6208
rect 38568 6190 38620 6196
rect 38474 4856 38530 4865
rect 38856 4826 38884 12106
rect 38948 11694 38976 13670
rect 39120 13456 39172 13462
rect 39120 13398 39172 13404
rect 39132 12102 39160 13398
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 39132 11694 39160 12038
rect 38936 11688 38988 11694
rect 38936 11630 38988 11636
rect 39120 11688 39172 11694
rect 39120 11630 39172 11636
rect 39028 10192 39080 10198
rect 39028 10134 39080 10140
rect 39040 9722 39068 10134
rect 39028 9716 39080 9722
rect 39028 9658 39080 9664
rect 39040 8412 39068 9658
rect 39120 8424 39172 8430
rect 39040 8384 39120 8412
rect 39120 8366 39172 8372
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39132 7546 39160 7822
rect 39120 7540 39172 7546
rect 39120 7482 39172 7488
rect 39028 7268 39080 7274
rect 39028 7210 39080 7216
rect 39040 6934 39068 7210
rect 39028 6928 39080 6934
rect 39028 6870 39080 6876
rect 39120 6928 39172 6934
rect 39120 6870 39172 6876
rect 39040 5914 39068 6870
rect 39132 6254 39160 6870
rect 39120 6248 39172 6254
rect 39120 6190 39172 6196
rect 39028 5908 39080 5914
rect 39028 5850 39080 5856
rect 38936 5840 38988 5846
rect 39132 5794 39160 6190
rect 38988 5788 39160 5794
rect 38936 5782 39160 5788
rect 38948 5766 39160 5782
rect 39120 5704 39172 5710
rect 39120 5646 39172 5652
rect 39028 5636 39080 5642
rect 39028 5578 39080 5584
rect 39040 5166 39068 5578
rect 39028 5160 39080 5166
rect 39028 5102 39080 5108
rect 38474 4791 38530 4800
rect 38844 4820 38896 4826
rect 38844 4762 38896 4768
rect 38292 4684 38344 4690
rect 38292 4626 38344 4632
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37936 4214 37964 4490
rect 38304 4282 38332 4626
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 38292 4276 38344 4282
rect 38292 4218 38344 4224
rect 37924 4208 37976 4214
rect 37924 4150 37976 4156
rect 38304 4078 38332 4218
rect 38292 4072 38344 4078
rect 38292 4014 38344 4020
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 38304 3602 38332 4014
rect 38580 3738 38608 4558
rect 38856 4078 38884 4762
rect 39132 4622 39160 5646
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 38844 4072 38896 4078
rect 38844 4014 38896 4020
rect 38568 3732 38620 3738
rect 38568 3674 38620 3680
rect 38292 3596 38344 3602
rect 38292 3538 38344 3544
rect 37738 3088 37794 3097
rect 38304 3058 38332 3538
rect 37738 3023 37794 3032
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 37556 2984 37608 2990
rect 37556 2926 37608 2932
rect 37832 2916 37884 2922
rect 37832 2858 37884 2864
rect 37844 2650 37872 2858
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 2650 38700 2790
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 37004 2644 37056 2650
rect 37004 2586 37056 2592
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 35992 2576 36044 2582
rect 35992 2518 36044 2524
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 34428 2508 34480 2514
rect 34428 2450 34480 2456
rect 35072 2508 35124 2514
rect 35072 2450 35124 2456
rect 34440 2310 34468 2450
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 32034 54 32168 82
rect 39118 82 39174 480
rect 39224 82 39252 18226
rect 39396 18216 39448 18222
rect 39396 18158 39448 18164
rect 39408 17746 39436 18158
rect 39396 17740 39448 17746
rect 39396 17682 39448 17688
rect 39408 17338 39436 17682
rect 39396 17332 39448 17338
rect 39396 17274 39448 17280
rect 39408 17134 39436 17274
rect 39396 17128 39448 17134
rect 39396 17070 39448 17076
rect 39408 16794 39436 17070
rect 39396 16788 39448 16794
rect 39396 16730 39448 16736
rect 39408 16182 39436 16730
rect 39592 16658 39620 22460
rect 39672 22442 39724 22448
rect 39856 22092 39908 22098
rect 39856 22034 39908 22040
rect 39868 21690 39896 22034
rect 39856 21684 39908 21690
rect 39856 21626 39908 21632
rect 39764 21412 39816 21418
rect 39764 21354 39816 21360
rect 39776 21010 39804 21354
rect 40328 21350 40356 23462
rect 40696 23322 40724 23666
rect 40684 23316 40736 23322
rect 40684 23258 40736 23264
rect 41248 23254 41276 23802
rect 42168 23474 42196 28070
rect 42524 27872 42576 27878
rect 42524 27814 42576 27820
rect 42536 26382 42564 27814
rect 42524 26376 42576 26382
rect 42524 26318 42576 26324
rect 42904 25809 42932 28966
rect 43088 28626 43116 29106
rect 43076 28620 43128 28626
rect 43076 28562 43128 28568
rect 43088 28218 43116 28562
rect 43168 28416 43220 28422
rect 43168 28358 43220 28364
rect 43076 28212 43128 28218
rect 43076 28154 43128 28160
rect 43076 27124 43128 27130
rect 43076 27066 43128 27072
rect 42890 25800 42946 25809
rect 42890 25735 42946 25744
rect 42432 24744 42484 24750
rect 42432 24686 42484 24692
rect 42444 24070 42472 24686
rect 42904 24070 42932 25735
rect 43088 24585 43116 27066
rect 43074 24576 43130 24585
rect 43074 24511 43130 24520
rect 42432 24064 42484 24070
rect 42432 24006 42484 24012
rect 42892 24064 42944 24070
rect 42892 24006 42944 24012
rect 42444 23662 42472 24006
rect 42432 23656 42484 23662
rect 42432 23598 42484 23604
rect 42168 23446 42472 23474
rect 41236 23248 41288 23254
rect 41236 23190 41288 23196
rect 40868 23180 40920 23186
rect 40868 23122 40920 23128
rect 40960 23180 41012 23186
rect 40960 23122 41012 23128
rect 40880 22506 40908 23122
rect 40868 22500 40920 22506
rect 40868 22442 40920 22448
rect 40776 22432 40828 22438
rect 40776 22374 40828 22380
rect 40788 21554 40816 22374
rect 40972 22234 41000 23122
rect 41604 22432 41656 22438
rect 41604 22374 41656 22380
rect 40960 22228 41012 22234
rect 40960 22170 41012 22176
rect 41420 22160 41472 22166
rect 41420 22102 41472 22108
rect 41052 22024 41104 22030
rect 41052 21966 41104 21972
rect 40776 21548 40828 21554
rect 40776 21490 40828 21496
rect 40500 21480 40552 21486
rect 40500 21422 40552 21428
rect 40316 21344 40368 21350
rect 40316 21286 40368 21292
rect 39764 21004 39816 21010
rect 39764 20946 39816 20952
rect 40328 20330 40356 21286
rect 40512 21146 40540 21422
rect 41064 21146 41092 21966
rect 41432 21690 41460 22102
rect 41512 22024 41564 22030
rect 41512 21966 41564 21972
rect 41420 21684 41472 21690
rect 41420 21626 41472 21632
rect 41420 21344 41472 21350
rect 41420 21286 41472 21292
rect 40500 21140 40552 21146
rect 40500 21082 40552 21088
rect 41052 21140 41104 21146
rect 41052 21082 41104 21088
rect 41432 21078 41460 21286
rect 41420 21072 41472 21078
rect 41420 21014 41472 21020
rect 41328 20936 41380 20942
rect 41328 20878 41380 20884
rect 40500 20392 40552 20398
rect 40500 20334 40552 20340
rect 40316 20324 40368 20330
rect 40316 20266 40368 20272
rect 40512 20058 40540 20334
rect 41340 20330 41368 20878
rect 41328 20324 41380 20330
rect 41328 20266 41380 20272
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 40040 19848 40092 19854
rect 40040 19790 40092 19796
rect 40052 18834 40080 19790
rect 41340 19514 41368 20266
rect 41432 20262 41460 21014
rect 41524 20874 41552 21966
rect 41512 20868 41564 20874
rect 41512 20810 41564 20816
rect 41420 20256 41472 20262
rect 41420 20198 41472 20204
rect 41420 19712 41472 19718
rect 41524 19700 41552 20810
rect 41616 19990 41644 22374
rect 42340 21548 42392 21554
rect 42340 21490 42392 21496
rect 42352 21146 42380 21490
rect 42340 21140 42392 21146
rect 42340 21082 42392 21088
rect 41880 20256 41932 20262
rect 41880 20198 41932 20204
rect 41892 19990 41920 20198
rect 41604 19984 41656 19990
rect 41604 19926 41656 19932
rect 41880 19984 41932 19990
rect 41880 19926 41932 19932
rect 41472 19672 41552 19700
rect 41420 19654 41472 19660
rect 41328 19508 41380 19514
rect 41328 19450 41380 19456
rect 41432 19242 41460 19654
rect 41420 19236 41472 19242
rect 41420 19178 41472 19184
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 40960 18896 41012 18902
rect 40960 18838 41012 18844
rect 39948 18828 40000 18834
rect 39948 18770 40000 18776
rect 40040 18828 40092 18834
rect 40040 18770 40092 18776
rect 39764 18624 39816 18630
rect 39764 18566 39816 18572
rect 39672 18216 39724 18222
rect 39672 18158 39724 18164
rect 39684 17814 39712 18158
rect 39672 17808 39724 17814
rect 39672 17750 39724 17756
rect 39580 16652 39632 16658
rect 39580 16594 39632 16600
rect 39592 16182 39620 16594
rect 39396 16176 39448 16182
rect 39396 16118 39448 16124
rect 39580 16176 39632 16182
rect 39580 16118 39632 16124
rect 39580 15496 39632 15502
rect 39580 15438 39632 15444
rect 39592 15162 39620 15438
rect 39580 15156 39632 15162
rect 39580 15098 39632 15104
rect 39672 14408 39724 14414
rect 39672 14350 39724 14356
rect 39684 14074 39712 14350
rect 39672 14068 39724 14074
rect 39672 14010 39724 14016
rect 39672 13184 39724 13190
rect 39672 13126 39724 13132
rect 39580 11620 39632 11626
rect 39580 11562 39632 11568
rect 39488 11144 39540 11150
rect 39488 11086 39540 11092
rect 39304 11076 39356 11082
rect 39304 11018 39356 11024
rect 39316 9926 39344 11018
rect 39500 10470 39528 11086
rect 39592 10674 39620 11562
rect 39580 10668 39632 10674
rect 39580 10610 39632 10616
rect 39488 10464 39540 10470
rect 39488 10406 39540 10412
rect 39304 9920 39356 9926
rect 39304 9862 39356 9868
rect 39500 9722 39528 10406
rect 39684 10130 39712 13126
rect 39672 10124 39724 10130
rect 39672 10066 39724 10072
rect 39488 9716 39540 9722
rect 39488 9658 39540 9664
rect 39488 8968 39540 8974
rect 39488 8910 39540 8916
rect 39500 8498 39528 8910
rect 39488 8492 39540 8498
rect 39488 8434 39540 8440
rect 39580 8288 39632 8294
rect 39580 8230 39632 8236
rect 39592 7478 39620 8230
rect 39580 7472 39632 7478
rect 39580 7414 39632 7420
rect 39580 5908 39632 5914
rect 39580 5850 39632 5856
rect 39304 5704 39356 5710
rect 39304 5646 39356 5652
rect 39316 5234 39344 5646
rect 39592 5370 39620 5850
rect 39684 5642 39712 10066
rect 39776 8566 39804 18566
rect 39960 17882 39988 18770
rect 40500 18624 40552 18630
rect 40500 18566 40552 18572
rect 40512 18222 40540 18566
rect 40500 18216 40552 18222
rect 40500 18158 40552 18164
rect 40972 18154 41000 18838
rect 41340 18426 41368 19110
rect 41616 18970 41644 19926
rect 41892 19514 41920 19926
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 41604 18964 41656 18970
rect 41604 18906 41656 18912
rect 41696 18828 41748 18834
rect 41696 18770 41748 18776
rect 41708 18426 41736 18770
rect 41328 18420 41380 18426
rect 41328 18362 41380 18368
rect 41696 18420 41748 18426
rect 41696 18362 41748 18368
rect 40684 18148 40736 18154
rect 40684 18090 40736 18096
rect 40960 18148 41012 18154
rect 40960 18090 41012 18096
rect 39948 17876 40000 17882
rect 39948 17818 40000 17824
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 39948 15632 40000 15638
rect 39948 15574 40000 15580
rect 39960 14822 39988 15574
rect 40052 15094 40080 17818
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40604 17270 40632 17614
rect 40592 17264 40644 17270
rect 40592 17206 40644 17212
rect 40224 16992 40276 16998
rect 40224 16934 40276 16940
rect 40316 16992 40368 16998
rect 40316 16934 40368 16940
rect 40236 16250 40264 16934
rect 40224 16244 40276 16250
rect 40224 16186 40276 16192
rect 40224 15972 40276 15978
rect 40224 15914 40276 15920
rect 40236 15162 40264 15914
rect 40328 15502 40356 16934
rect 40604 16794 40632 17206
rect 40696 17202 40724 18090
rect 40972 17814 41000 18090
rect 40960 17808 41012 17814
rect 40960 17750 41012 17756
rect 40684 17196 40736 17202
rect 40684 17138 40736 17144
rect 40972 16998 41000 17750
rect 41696 17196 41748 17202
rect 41696 17138 41748 17144
rect 40960 16992 41012 16998
rect 40960 16934 41012 16940
rect 40592 16788 40644 16794
rect 40592 16730 40644 16736
rect 40592 16516 40644 16522
rect 40592 16458 40644 16464
rect 40604 16114 40632 16458
rect 40592 16108 40644 16114
rect 40592 16050 40644 16056
rect 40776 16108 40828 16114
rect 40776 16050 40828 16056
rect 40316 15496 40368 15502
rect 40316 15438 40368 15444
rect 40224 15156 40276 15162
rect 40224 15098 40276 15104
rect 40040 15088 40092 15094
rect 40040 15030 40092 15036
rect 40236 14890 40264 15098
rect 40592 15020 40644 15026
rect 40592 14962 40644 14968
rect 40224 14884 40276 14890
rect 40224 14826 40276 14832
rect 39948 14816 40000 14822
rect 39948 14758 40000 14764
rect 39960 14550 39988 14758
rect 40604 14618 40632 14962
rect 40592 14612 40644 14618
rect 40592 14554 40644 14560
rect 39948 14544 40000 14550
rect 39948 14486 40000 14492
rect 39960 13938 39988 14486
rect 40788 14482 40816 16050
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40880 15026 40908 15438
rect 40868 15020 40920 15026
rect 40868 14962 40920 14968
rect 40776 14476 40828 14482
rect 40776 14418 40828 14424
rect 39948 13932 40000 13938
rect 39948 13874 40000 13880
rect 40972 13462 41000 16934
rect 41708 16794 41736 17138
rect 41696 16788 41748 16794
rect 41696 16730 41748 16736
rect 42444 16658 42472 23446
rect 43180 23050 43208 28358
rect 43272 27538 43300 30330
rect 43350 30288 43406 30297
rect 43350 30223 43406 30232
rect 43364 29714 43392 30223
rect 43352 29708 43404 29714
rect 43352 29650 43404 29656
rect 43364 29306 43392 29650
rect 43352 29300 43404 29306
rect 43352 29242 43404 29248
rect 43260 27532 43312 27538
rect 43312 27492 43392 27520
rect 43260 27474 43312 27480
rect 43260 27328 43312 27334
rect 43260 27270 43312 27276
rect 43272 26994 43300 27270
rect 43364 27130 43392 27492
rect 43352 27124 43404 27130
rect 43352 27066 43404 27072
rect 43260 26988 43312 26994
rect 43260 26930 43312 26936
rect 43640 26858 43668 33322
rect 43732 33134 43760 35430
rect 43812 34468 43864 34474
rect 43812 34410 43864 34416
rect 43824 34134 43852 34410
rect 43812 34128 43864 34134
rect 43812 34070 43864 34076
rect 43824 33658 43852 34070
rect 43812 33652 43864 33658
rect 43812 33594 43864 33600
rect 43732 33106 43852 33134
rect 43824 32978 43852 33106
rect 43812 32972 43864 32978
rect 43812 32914 43864 32920
rect 43824 32230 43852 32914
rect 43812 32224 43864 32230
rect 43812 32166 43864 32172
rect 43720 31204 43772 31210
rect 43720 31146 43772 31152
rect 43732 31113 43760 31146
rect 43718 31104 43774 31113
rect 43718 31039 43774 31048
rect 43720 27464 43772 27470
rect 43720 27406 43772 27412
rect 43536 26852 43588 26858
rect 43536 26794 43588 26800
rect 43628 26852 43680 26858
rect 43628 26794 43680 26800
rect 43548 26518 43576 26794
rect 43536 26512 43588 26518
rect 43536 26454 43588 26460
rect 43548 26042 43576 26454
rect 43732 26382 43760 27406
rect 43628 26376 43680 26382
rect 43628 26318 43680 26324
rect 43720 26376 43772 26382
rect 43720 26318 43772 26324
rect 43536 26036 43588 26042
rect 43536 25978 43588 25984
rect 43548 25770 43576 25978
rect 43640 25974 43668 26318
rect 43628 25968 43680 25974
rect 43628 25910 43680 25916
rect 43536 25764 43588 25770
rect 43536 25706 43588 25712
rect 43352 25696 43404 25702
rect 43732 25650 43760 26318
rect 43352 25638 43404 25644
rect 43260 24608 43312 24614
rect 43260 24550 43312 24556
rect 43272 23866 43300 24550
rect 43260 23860 43312 23866
rect 43260 23802 43312 23808
rect 43272 23576 43300 23802
rect 43364 23730 43392 25638
rect 43456 25622 43760 25650
rect 43456 25294 43484 25622
rect 43536 25424 43588 25430
rect 43824 25401 43852 32166
rect 43916 31346 43944 36518
rect 44364 36032 44416 36038
rect 44364 35974 44416 35980
rect 44376 35562 44404 35974
rect 44272 35556 44324 35562
rect 44272 35498 44324 35504
rect 44364 35556 44416 35562
rect 44364 35498 44416 35504
rect 44284 35290 44312 35498
rect 44272 35284 44324 35290
rect 44272 35226 44324 35232
rect 44376 34474 44404 35498
rect 44364 34468 44416 34474
rect 44364 34410 44416 34416
rect 44272 34400 44324 34406
rect 44272 34342 44324 34348
rect 44284 34202 44312 34342
rect 44272 34196 44324 34202
rect 44272 34138 44324 34144
rect 44088 33992 44140 33998
rect 44088 33934 44140 33940
rect 44100 33658 44128 33934
rect 44088 33652 44140 33658
rect 44088 33594 44140 33600
rect 44468 33134 44496 38694
rect 44640 38004 44692 38010
rect 44640 37946 44692 37952
rect 44548 34604 44600 34610
rect 44548 34546 44600 34552
rect 44560 34202 44588 34546
rect 44548 34196 44600 34202
rect 44548 34138 44600 34144
rect 44652 33134 44680 37946
rect 44732 37936 44784 37942
rect 44732 37878 44784 37884
rect 44744 37262 44772 37878
rect 44732 37256 44784 37262
rect 44732 37198 44784 37204
rect 44744 34474 44772 37198
rect 44836 34542 44864 44231
rect 44928 35193 44956 44775
rect 49528 44470 49556 48447
rect 49516 44464 49568 44470
rect 49516 44406 49568 44412
rect 49514 39128 49570 39137
rect 49514 39063 49570 39072
rect 46204 38344 46256 38350
rect 46204 38286 46256 38292
rect 45100 37392 45152 37398
rect 45100 37334 45152 37340
rect 45112 36854 45140 37334
rect 46216 37262 46244 38286
rect 45928 37256 45980 37262
rect 45928 37198 45980 37204
rect 46204 37256 46256 37262
rect 46204 37198 46256 37204
rect 45744 37120 45796 37126
rect 45744 37062 45796 37068
rect 45100 36848 45152 36854
rect 45100 36790 45152 36796
rect 45112 36310 45140 36790
rect 45192 36644 45244 36650
rect 45192 36586 45244 36592
rect 45100 36304 45152 36310
rect 45100 36246 45152 36252
rect 45112 35834 45140 36246
rect 45204 36174 45232 36586
rect 45192 36168 45244 36174
rect 45192 36110 45244 36116
rect 45100 35828 45152 35834
rect 45100 35770 45152 35776
rect 45008 35760 45060 35766
rect 45008 35702 45060 35708
rect 44914 35184 44970 35193
rect 44914 35119 44970 35128
rect 44824 34536 44876 34542
rect 44824 34478 44876 34484
rect 44732 34468 44784 34474
rect 44732 34410 44784 34416
rect 44836 33862 44864 34478
rect 44824 33856 44876 33862
rect 44824 33798 44876 33804
rect 45020 33658 45048 35702
rect 45204 35698 45232 36110
rect 45652 36032 45704 36038
rect 45652 35974 45704 35980
rect 45664 35834 45692 35974
rect 45652 35828 45704 35834
rect 45652 35770 45704 35776
rect 45192 35692 45244 35698
rect 45192 35634 45244 35640
rect 45100 35216 45152 35222
rect 45100 35158 45152 35164
rect 45112 34678 45140 35158
rect 45204 35086 45232 35634
rect 45192 35080 45244 35086
rect 45192 35022 45244 35028
rect 45204 34746 45232 35022
rect 45376 34944 45428 34950
rect 45376 34886 45428 34892
rect 45192 34740 45244 34746
rect 45192 34682 45244 34688
rect 45100 34672 45152 34678
rect 45100 34614 45152 34620
rect 45100 34400 45152 34406
rect 45100 34342 45152 34348
rect 45112 33998 45140 34342
rect 45388 34066 45416 34886
rect 45376 34060 45428 34066
rect 45376 34002 45428 34008
rect 45100 33992 45152 33998
rect 45100 33934 45152 33940
rect 45388 33658 45416 34002
rect 45008 33652 45060 33658
rect 45008 33594 45060 33600
rect 45376 33652 45428 33658
rect 45376 33594 45428 33600
rect 45020 33454 45048 33594
rect 45008 33448 45060 33454
rect 45008 33390 45060 33396
rect 44732 33312 44784 33318
rect 44732 33254 44784 33260
rect 44376 33106 44496 33134
rect 44560 33106 44680 33134
rect 43904 31340 43956 31346
rect 43904 31282 43956 31288
rect 44376 30394 44404 33106
rect 44456 32768 44508 32774
rect 44456 32710 44508 32716
rect 44468 32434 44496 32710
rect 44456 32428 44508 32434
rect 44456 32370 44508 32376
rect 44364 30388 44416 30394
rect 44364 30330 44416 30336
rect 44560 30240 44588 33106
rect 44744 32910 44772 33254
rect 44824 33040 44876 33046
rect 44824 32982 44876 32988
rect 44732 32904 44784 32910
rect 44732 32846 44784 32852
rect 44744 32026 44772 32846
rect 44836 32298 44864 32982
rect 45756 32978 45784 37062
rect 45940 36378 45968 37198
rect 46572 36576 46624 36582
rect 46572 36518 46624 36524
rect 46584 36378 46612 36518
rect 45928 36372 45980 36378
rect 45928 36314 45980 36320
rect 46572 36372 46624 36378
rect 46572 36314 46624 36320
rect 46388 36236 46440 36242
rect 46388 36178 46440 36184
rect 46400 35766 46428 36178
rect 46388 35760 46440 35766
rect 46388 35702 46440 35708
rect 46110 35456 46166 35465
rect 46110 35391 46166 35400
rect 46020 33856 46072 33862
rect 46020 33798 46072 33804
rect 45744 32972 45796 32978
rect 45744 32914 45796 32920
rect 45008 32904 45060 32910
rect 45008 32846 45060 32852
rect 44824 32292 44876 32298
rect 44824 32234 44876 32240
rect 44732 32020 44784 32026
rect 44732 31962 44784 31968
rect 45020 31958 45048 32846
rect 45560 32360 45612 32366
rect 45560 32302 45612 32308
rect 45192 32224 45244 32230
rect 45192 32166 45244 32172
rect 45204 31958 45232 32166
rect 45008 31952 45060 31958
rect 45008 31894 45060 31900
rect 45192 31952 45244 31958
rect 45192 31894 45244 31900
rect 44916 31748 44968 31754
rect 44916 31690 44968 31696
rect 44824 31136 44876 31142
rect 44824 31078 44876 31084
rect 44640 30864 44692 30870
rect 44640 30806 44692 30812
rect 44468 30212 44588 30240
rect 44364 28076 44416 28082
rect 44364 28018 44416 28024
rect 43904 27668 43956 27674
rect 43904 27610 43956 27616
rect 43916 26994 43944 27610
rect 44376 27538 44404 28018
rect 44468 28014 44496 30212
rect 44652 30122 44680 30806
rect 44548 30116 44600 30122
rect 44548 30058 44600 30064
rect 44640 30116 44692 30122
rect 44640 30058 44692 30064
rect 44560 28762 44588 30058
rect 44652 29850 44680 30058
rect 44640 29844 44692 29850
rect 44640 29786 44692 29792
rect 44652 29306 44680 29786
rect 44640 29300 44692 29306
rect 44640 29242 44692 29248
rect 44652 29034 44680 29242
rect 44836 29170 44864 31078
rect 44928 29170 44956 31690
rect 45020 30258 45048 31894
rect 45204 31482 45232 31894
rect 45192 31476 45244 31482
rect 45192 31418 45244 31424
rect 45284 31340 45336 31346
rect 45284 31282 45336 31288
rect 45296 31210 45324 31282
rect 45100 31204 45152 31210
rect 45100 31146 45152 31152
rect 45284 31204 45336 31210
rect 45284 31146 45336 31152
rect 45112 30870 45140 31146
rect 45100 30864 45152 30870
rect 45100 30806 45152 30812
rect 45100 30388 45152 30394
rect 45100 30330 45152 30336
rect 45008 30252 45060 30258
rect 45008 30194 45060 30200
rect 44824 29164 44876 29170
rect 44824 29106 44876 29112
rect 44916 29164 44968 29170
rect 44916 29106 44968 29112
rect 44640 29028 44692 29034
rect 44640 28970 44692 28976
rect 44836 28762 44864 29106
rect 44548 28756 44600 28762
rect 44548 28698 44600 28704
rect 44824 28756 44876 28762
rect 44824 28698 44876 28704
rect 44456 28008 44508 28014
rect 44456 27950 44508 27956
rect 44640 28008 44692 28014
rect 44640 27950 44692 27956
rect 44652 27878 44680 27950
rect 44640 27872 44692 27878
rect 44640 27814 44692 27820
rect 44456 27600 44508 27606
rect 44456 27542 44508 27548
rect 44364 27532 44416 27538
rect 44364 27474 44416 27480
rect 43904 26988 43956 26994
rect 43904 26930 43956 26936
rect 43916 26586 43944 26930
rect 44376 26586 44404 27474
rect 44468 26790 44496 27542
rect 44456 26784 44508 26790
rect 44456 26726 44508 26732
rect 43904 26580 43956 26586
rect 43904 26522 43956 26528
rect 44364 26580 44416 26586
rect 44364 26522 44416 26528
rect 43536 25366 43588 25372
rect 43810 25392 43866 25401
rect 43444 25288 43496 25294
rect 43444 25230 43496 25236
rect 43456 24954 43484 25230
rect 43444 24948 43496 24954
rect 43444 24890 43496 24896
rect 43548 24614 43576 25366
rect 43810 25327 43866 25336
rect 43628 25220 43680 25226
rect 43628 25162 43680 25168
rect 43536 24608 43588 24614
rect 43536 24550 43588 24556
rect 43548 24410 43576 24550
rect 43536 24404 43588 24410
rect 43536 24346 43588 24352
rect 43640 23730 43668 25162
rect 43916 24868 43944 26522
rect 44468 26466 44496 26726
rect 44376 26438 44496 26466
rect 43996 24880 44048 24886
rect 43916 24840 43996 24868
rect 43996 24822 44048 24828
rect 44376 24342 44404 26438
rect 44548 25152 44600 25158
rect 44548 25094 44600 25100
rect 44560 24818 44588 25094
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 44454 24576 44510 24585
rect 44454 24511 44510 24520
rect 44364 24336 44416 24342
rect 44364 24278 44416 24284
rect 44272 24200 44324 24206
rect 44272 24142 44324 24148
rect 43352 23724 43404 23730
rect 43352 23666 43404 23672
rect 43628 23724 43680 23730
rect 43628 23666 43680 23672
rect 43352 23588 43404 23594
rect 43272 23548 43352 23576
rect 43352 23530 43404 23536
rect 43640 23186 43668 23666
rect 44284 23322 44312 24142
rect 44376 23526 44404 24278
rect 44364 23520 44416 23526
rect 44364 23462 44416 23468
rect 44272 23316 44324 23322
rect 44272 23258 44324 23264
rect 43628 23180 43680 23186
rect 43628 23122 43680 23128
rect 43996 23180 44048 23186
rect 43996 23122 44048 23128
rect 43168 23044 43220 23050
rect 43168 22986 43220 22992
rect 43904 23044 43956 23050
rect 43904 22986 43956 22992
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42628 19258 42656 22918
rect 42708 22704 42760 22710
rect 42708 22646 42760 22652
rect 43168 22704 43220 22710
rect 43168 22646 43220 22652
rect 42720 21690 42748 22646
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 43088 22234 43116 22578
rect 43180 22506 43208 22646
rect 43168 22500 43220 22506
rect 43168 22442 43220 22448
rect 43444 22432 43496 22438
rect 43444 22374 43496 22380
rect 43076 22228 43128 22234
rect 43076 22170 43128 22176
rect 43352 22228 43404 22234
rect 43352 22170 43404 22176
rect 42984 21956 43036 21962
rect 42984 21898 43036 21904
rect 42708 21684 42760 21690
rect 42708 21626 42760 21632
rect 42892 21616 42944 21622
rect 42892 21558 42944 21564
rect 42798 21312 42854 21321
rect 42798 21247 42854 21256
rect 42628 19230 42748 19258
rect 42616 19168 42668 19174
rect 42616 19110 42668 19116
rect 42628 17338 42656 19110
rect 42616 17332 42668 17338
rect 42616 17274 42668 17280
rect 41144 16652 41196 16658
rect 41144 16594 41196 16600
rect 42432 16652 42484 16658
rect 42432 16594 42484 16600
rect 41156 15706 41184 16594
rect 42340 16584 42392 16590
rect 42340 16526 42392 16532
rect 42156 16448 42208 16454
rect 42156 16390 42208 16396
rect 42168 16046 42196 16390
rect 42156 16040 42208 16046
rect 42156 15982 42208 15988
rect 41144 15700 41196 15706
rect 41144 15642 41196 15648
rect 42352 15570 42380 16526
rect 42444 16250 42472 16594
rect 42432 16244 42484 16250
rect 42432 16186 42484 16192
rect 42340 15564 42392 15570
rect 42340 15506 42392 15512
rect 42248 15360 42300 15366
rect 42248 15302 42300 15308
rect 41972 14952 42024 14958
rect 41972 14894 42024 14900
rect 41696 14884 41748 14890
rect 41696 14826 41748 14832
rect 41604 14476 41656 14482
rect 41604 14418 41656 14424
rect 41616 14278 41644 14418
rect 41420 14272 41472 14278
rect 41420 14214 41472 14220
rect 41604 14272 41656 14278
rect 41604 14214 41656 14220
rect 41432 13938 41460 14214
rect 41420 13932 41472 13938
rect 41420 13874 41472 13880
rect 41432 13814 41460 13874
rect 41432 13786 41552 13814
rect 41524 13530 41552 13786
rect 41512 13524 41564 13530
rect 41512 13466 41564 13472
rect 40960 13456 41012 13462
rect 40880 13416 40960 13444
rect 39856 13388 39908 13394
rect 39856 13330 39908 13336
rect 39868 12918 39896 13330
rect 40316 13320 40368 13326
rect 40316 13262 40368 13268
rect 39856 12912 39908 12918
rect 39856 12854 39908 12860
rect 40328 12646 40356 13262
rect 40880 12918 40908 13416
rect 40960 13398 41012 13404
rect 40960 13184 41012 13190
rect 40960 13126 41012 13132
rect 40868 12912 40920 12918
rect 40868 12854 40920 12860
rect 40316 12640 40368 12646
rect 40316 12582 40368 12588
rect 40328 12442 40356 12582
rect 40316 12436 40368 12442
rect 40316 12378 40368 12384
rect 40880 12374 40908 12854
rect 40972 12782 41000 13126
rect 41616 12986 41644 14214
rect 41708 13734 41736 14826
rect 41880 14816 41932 14822
rect 41880 14758 41932 14764
rect 41696 13728 41748 13734
rect 41696 13670 41748 13676
rect 41892 13433 41920 14758
rect 41984 14550 42012 14894
rect 42260 14890 42288 15302
rect 42352 15162 42380 15506
rect 42340 15156 42392 15162
rect 42340 15098 42392 15104
rect 42248 14884 42300 14890
rect 42248 14826 42300 14832
rect 41972 14544 42024 14550
rect 41972 14486 42024 14492
rect 42064 14476 42116 14482
rect 42064 14418 42116 14424
rect 42076 13734 42104 14418
rect 41972 13728 42024 13734
rect 41972 13670 42024 13676
rect 42064 13728 42116 13734
rect 42064 13670 42116 13676
rect 41878 13424 41934 13433
rect 41878 13359 41934 13368
rect 41604 12980 41656 12986
rect 41604 12922 41656 12928
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 40868 12368 40920 12374
rect 40868 12310 40920 12316
rect 40592 12232 40644 12238
rect 40592 12174 40644 12180
rect 40500 11688 40552 11694
rect 40500 11630 40552 11636
rect 39948 11144 40000 11150
rect 39948 11086 40000 11092
rect 39856 10804 39908 10810
rect 39856 10746 39908 10752
rect 39868 9178 39896 10746
rect 39960 10470 39988 11086
rect 40512 11014 40540 11630
rect 40604 11558 40632 12174
rect 40880 11898 40908 12310
rect 40868 11892 40920 11898
rect 40868 11834 40920 11840
rect 40592 11552 40644 11558
rect 40592 11494 40644 11500
rect 40604 11354 40632 11494
rect 40592 11348 40644 11354
rect 40592 11290 40644 11296
rect 40880 11286 40908 11834
rect 40972 11694 41000 12718
rect 41984 12646 42012 13670
rect 41972 12640 42024 12646
rect 41972 12582 42024 12588
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 40960 11688 41012 11694
rect 40960 11630 41012 11636
rect 40868 11280 40920 11286
rect 40868 11222 40920 11228
rect 40500 11008 40552 11014
rect 40500 10950 40552 10956
rect 40880 10810 40908 11222
rect 40868 10804 40920 10810
rect 40868 10746 40920 10752
rect 40880 10538 40908 10746
rect 40868 10532 40920 10538
rect 40868 10474 40920 10480
rect 39948 10464 40000 10470
rect 39948 10406 40000 10412
rect 39960 10266 39988 10406
rect 39948 10260 40000 10266
rect 39948 10202 40000 10208
rect 40972 10130 41000 11630
rect 41604 11008 41656 11014
rect 41604 10950 41656 10956
rect 41616 10810 41644 10950
rect 41604 10804 41656 10810
rect 41604 10746 41656 10752
rect 41144 10668 41196 10674
rect 41144 10610 41196 10616
rect 41156 10266 41184 10610
rect 41144 10260 41196 10266
rect 41144 10202 41196 10208
rect 41800 10198 41828 12038
rect 41788 10192 41840 10198
rect 41788 10134 41840 10140
rect 40132 10124 40184 10130
rect 40132 10066 40184 10072
rect 40960 10124 41012 10130
rect 40960 10066 41012 10072
rect 40144 9654 40172 10066
rect 40972 9722 41000 10066
rect 40960 9716 41012 9722
rect 40960 9658 41012 9664
rect 40132 9648 40184 9654
rect 40132 9590 40184 9596
rect 41800 9178 41828 10134
rect 41880 9716 41932 9722
rect 41880 9658 41932 9664
rect 39856 9172 39908 9178
rect 39856 9114 39908 9120
rect 41788 9172 41840 9178
rect 41788 9114 41840 9120
rect 39764 8560 39816 8566
rect 39764 8502 39816 8508
rect 39868 8294 39896 9114
rect 41892 9110 41920 9658
rect 41984 9364 42012 12582
rect 42076 12442 42104 13670
rect 42156 13184 42208 13190
rect 42156 13126 42208 13132
rect 42168 12850 42196 13126
rect 42260 12850 42288 14826
rect 42432 14272 42484 14278
rect 42432 14214 42484 14220
rect 42340 13796 42392 13802
rect 42340 13738 42392 13744
rect 42156 12844 42208 12850
rect 42156 12786 42208 12792
rect 42248 12844 42300 12850
rect 42248 12786 42300 12792
rect 42168 12442 42196 12786
rect 42064 12436 42116 12442
rect 42064 12378 42116 12384
rect 42156 12436 42208 12442
rect 42156 12378 42208 12384
rect 42156 12300 42208 12306
rect 42156 12242 42208 12248
rect 42064 11552 42116 11558
rect 42064 11494 42116 11500
rect 42076 10742 42104 11494
rect 42168 11354 42196 12242
rect 42260 11898 42288 12786
rect 42248 11892 42300 11898
rect 42248 11834 42300 11840
rect 42260 11626 42288 11834
rect 42352 11762 42380 13738
rect 42444 11830 42472 14214
rect 42616 13388 42668 13394
rect 42616 13330 42668 13336
rect 42524 12844 42576 12850
rect 42524 12786 42576 12792
rect 42536 12646 42564 12786
rect 42524 12640 42576 12646
rect 42524 12582 42576 12588
rect 42628 12442 42656 13330
rect 42616 12436 42668 12442
rect 42616 12378 42668 12384
rect 42432 11824 42484 11830
rect 42432 11766 42484 11772
rect 42340 11756 42392 11762
rect 42340 11698 42392 11704
rect 42248 11620 42300 11626
rect 42248 11562 42300 11568
rect 42156 11348 42208 11354
rect 42156 11290 42208 11296
rect 42064 10736 42116 10742
rect 42064 10678 42116 10684
rect 42260 10606 42288 11562
rect 42248 10600 42300 10606
rect 42248 10542 42300 10548
rect 42260 10198 42288 10542
rect 42524 10464 42576 10470
rect 42524 10406 42576 10412
rect 42248 10192 42300 10198
rect 42248 10134 42300 10140
rect 42260 9722 42288 10134
rect 42248 9716 42300 9722
rect 42248 9658 42300 9664
rect 42536 9586 42564 10406
rect 42524 9580 42576 9586
rect 42524 9522 42576 9528
rect 42156 9376 42208 9382
rect 41984 9336 42156 9364
rect 42156 9318 42208 9324
rect 41880 9104 41932 9110
rect 41880 9046 41932 9052
rect 41788 8968 41840 8974
rect 41788 8910 41840 8916
rect 41800 8634 41828 8910
rect 41892 8634 41920 9046
rect 41788 8628 41840 8634
rect 41788 8570 41840 8576
rect 41880 8628 41932 8634
rect 41880 8570 41932 8576
rect 42168 8362 42196 9318
rect 42536 9178 42564 9522
rect 42524 9172 42576 9178
rect 42524 9114 42576 9120
rect 41512 8356 41564 8362
rect 41512 8298 41564 8304
rect 42156 8356 42208 8362
rect 42156 8298 42208 8304
rect 39856 8288 39908 8294
rect 39856 8230 39908 8236
rect 39868 8022 39896 8230
rect 39856 8016 39908 8022
rect 39856 7958 39908 7964
rect 39868 7206 39896 7958
rect 41524 7886 41552 8298
rect 41696 7948 41748 7954
rect 41696 7890 41748 7896
rect 42340 7948 42392 7954
rect 42340 7890 42392 7896
rect 41512 7880 41564 7886
rect 41512 7822 41564 7828
rect 40224 7812 40276 7818
rect 40224 7754 40276 7760
rect 39856 7200 39908 7206
rect 39856 7142 39908 7148
rect 40236 6934 40264 7754
rect 40684 7404 40736 7410
rect 40684 7346 40736 7352
rect 40696 6934 40724 7346
rect 40868 7200 40920 7206
rect 40868 7142 40920 7148
rect 41144 7200 41196 7206
rect 41144 7142 41196 7148
rect 40224 6928 40276 6934
rect 40224 6870 40276 6876
rect 40684 6928 40736 6934
rect 40684 6870 40736 6876
rect 40132 6180 40184 6186
rect 40132 6122 40184 6128
rect 39764 6112 39816 6118
rect 39764 6054 39816 6060
rect 39672 5636 39724 5642
rect 39672 5578 39724 5584
rect 39580 5364 39632 5370
rect 39580 5306 39632 5312
rect 39304 5228 39356 5234
rect 39304 5170 39356 5176
rect 39488 4752 39540 4758
rect 39488 4694 39540 4700
rect 39500 4282 39528 4694
rect 39488 4276 39540 4282
rect 39488 4218 39540 4224
rect 39396 4004 39448 4010
rect 39396 3946 39448 3952
rect 39408 3738 39436 3946
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39408 3058 39436 3674
rect 39592 3670 39620 5306
rect 39776 4758 39804 6054
rect 40144 5710 40172 6122
rect 40236 5914 40264 6870
rect 40696 6118 40724 6870
rect 40684 6112 40736 6118
rect 40684 6054 40736 6060
rect 40224 5908 40276 5914
rect 40224 5850 40276 5856
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 40144 5234 40172 5646
rect 40224 5568 40276 5574
rect 40224 5510 40276 5516
rect 40236 5370 40264 5510
rect 40224 5364 40276 5370
rect 40224 5306 40276 5312
rect 40696 5302 40724 6054
rect 40880 5914 40908 7142
rect 41052 6656 41104 6662
rect 41052 6598 41104 6604
rect 41064 6322 41092 6598
rect 41052 6316 41104 6322
rect 41052 6258 41104 6264
rect 41156 5914 41184 7142
rect 41512 6316 41564 6322
rect 41512 6258 41564 6264
rect 40868 5908 40920 5914
rect 40868 5850 40920 5856
rect 41144 5908 41196 5914
rect 41144 5850 41196 5856
rect 40880 5302 40908 5850
rect 41524 5710 41552 6258
rect 41708 6186 41736 7890
rect 42352 7546 42380 7890
rect 42616 7880 42668 7886
rect 42616 7822 42668 7828
rect 42628 7546 42656 7822
rect 42340 7540 42392 7546
rect 42340 7482 42392 7488
rect 42616 7540 42668 7546
rect 42616 7482 42668 7488
rect 42156 7336 42208 7342
rect 42156 7278 42208 7284
rect 42168 7002 42196 7278
rect 42352 7002 42380 7482
rect 42720 7041 42748 19230
rect 42812 18834 42840 21247
rect 42904 20602 42932 21558
rect 42996 21554 43024 21898
rect 42984 21548 43036 21554
rect 42984 21490 43036 21496
rect 42892 20596 42944 20602
rect 42892 20538 42944 20544
rect 42904 20262 42932 20538
rect 43168 20460 43220 20466
rect 43168 20402 43220 20408
rect 43076 20324 43128 20330
rect 43076 20266 43128 20272
rect 42892 20256 42944 20262
rect 42892 20198 42944 20204
rect 43088 20058 43116 20266
rect 43076 20052 43128 20058
rect 43076 19994 43128 20000
rect 42984 19236 43036 19242
rect 43180 19224 43208 20402
rect 43260 19372 43312 19378
rect 43260 19314 43312 19320
rect 43036 19196 43208 19224
rect 42984 19178 43036 19184
rect 43180 18970 43208 19196
rect 43168 18964 43220 18970
rect 43168 18906 43220 18912
rect 42800 18828 42852 18834
rect 42800 18770 42852 18776
rect 42812 18426 42840 18770
rect 42800 18420 42852 18426
rect 42800 18362 42852 18368
rect 43272 17746 43300 19314
rect 43364 18290 43392 22170
rect 43456 22166 43484 22374
rect 43444 22160 43496 22166
rect 43444 22102 43496 22108
rect 43536 22160 43588 22166
rect 43536 22102 43588 22108
rect 43456 21690 43484 22102
rect 43444 21684 43496 21690
rect 43444 21626 43496 21632
rect 43548 21554 43576 22102
rect 43536 21548 43588 21554
rect 43536 21490 43588 21496
rect 43720 19984 43772 19990
rect 43720 19926 43772 19932
rect 43444 19848 43496 19854
rect 43444 19790 43496 19796
rect 43628 19848 43680 19854
rect 43628 19790 43680 19796
rect 43456 19242 43484 19790
rect 43640 19378 43668 19790
rect 43628 19372 43680 19378
rect 43628 19314 43680 19320
rect 43444 19236 43496 19242
rect 43444 19178 43496 19184
rect 43732 19174 43760 19926
rect 43720 19168 43772 19174
rect 43720 19110 43772 19116
rect 43628 18896 43680 18902
rect 43628 18838 43680 18844
rect 43640 18630 43668 18838
rect 43732 18766 43760 19110
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43628 18624 43680 18630
rect 43628 18566 43680 18572
rect 43352 18284 43404 18290
rect 43352 18226 43404 18232
rect 43444 18216 43496 18222
rect 43444 18158 43496 18164
rect 43456 17882 43484 18158
rect 43640 18154 43668 18566
rect 43812 18284 43864 18290
rect 43812 18226 43864 18232
rect 43628 18148 43680 18154
rect 43628 18090 43680 18096
rect 43444 17876 43496 17882
rect 43444 17818 43496 17824
rect 43536 17876 43588 17882
rect 43536 17818 43588 17824
rect 43260 17740 43312 17746
rect 43180 17700 43260 17728
rect 43180 17270 43208 17700
rect 43260 17682 43312 17688
rect 43260 17536 43312 17542
rect 43260 17478 43312 17484
rect 43272 17338 43300 17478
rect 43260 17332 43312 17338
rect 43260 17274 43312 17280
rect 43168 17264 43220 17270
rect 43168 17206 43220 17212
rect 43272 16998 43300 17274
rect 43548 17066 43576 17818
rect 43824 17542 43852 18226
rect 43628 17536 43680 17542
rect 43628 17478 43680 17484
rect 43812 17536 43864 17542
rect 43812 17478 43864 17484
rect 43536 17060 43588 17066
rect 43536 17002 43588 17008
rect 43260 16992 43312 16998
rect 43260 16934 43312 16940
rect 43548 16794 43576 17002
rect 43536 16788 43588 16794
rect 43536 16730 43588 16736
rect 43444 16652 43496 16658
rect 43444 16594 43496 16600
rect 43456 16250 43484 16594
rect 43444 16244 43496 16250
rect 43444 16186 43496 16192
rect 43536 15972 43588 15978
rect 43536 15914 43588 15920
rect 43548 15638 43576 15914
rect 42892 15632 42944 15638
rect 42892 15574 42944 15580
rect 43536 15632 43588 15638
rect 43536 15574 43588 15580
rect 42904 15162 42932 15574
rect 43444 15496 43496 15502
rect 43444 15438 43496 15444
rect 42892 15156 42944 15162
rect 42892 15098 42944 15104
rect 42904 14006 42932 15098
rect 43456 14618 43484 15438
rect 43536 15088 43588 15094
rect 43536 15030 43588 15036
rect 43548 14890 43576 15030
rect 43536 14884 43588 14890
rect 43536 14826 43588 14832
rect 43548 14618 43576 14826
rect 43444 14612 43496 14618
rect 43444 14554 43496 14560
rect 43536 14612 43588 14618
rect 43536 14554 43588 14560
rect 42892 14000 42944 14006
rect 42892 13942 42944 13948
rect 43548 13814 43576 14554
rect 43456 13786 43576 13814
rect 43456 13462 43484 13786
rect 43444 13456 43496 13462
rect 43444 13398 43496 13404
rect 43456 12986 43484 13398
rect 43536 13184 43588 13190
rect 43536 13126 43588 13132
rect 43444 12980 43496 12986
rect 43444 12922 43496 12928
rect 43260 12300 43312 12306
rect 43260 12242 43312 12248
rect 43272 11898 43300 12242
rect 43456 11898 43484 12922
rect 43548 12714 43576 13126
rect 43536 12708 43588 12714
rect 43536 12650 43588 12656
rect 43548 12442 43576 12650
rect 43536 12436 43588 12442
rect 43536 12378 43588 12384
rect 43640 12238 43668 17478
rect 43824 16726 43852 17478
rect 43812 16720 43864 16726
rect 43812 16662 43864 16668
rect 43916 16658 43944 22986
rect 44008 22778 44036 23122
rect 43996 22772 44048 22778
rect 43996 22714 44048 22720
rect 44468 22574 44496 24511
rect 44560 23866 44588 24754
rect 44548 23860 44600 23866
rect 44548 23802 44600 23808
rect 44652 23186 44680 27814
rect 45112 26976 45140 30330
rect 45296 27062 45324 31146
rect 45468 30728 45520 30734
rect 45468 30670 45520 30676
rect 45480 30394 45508 30670
rect 45468 30388 45520 30394
rect 45468 30330 45520 30336
rect 45572 29646 45600 32302
rect 45756 32230 45784 32914
rect 45836 32768 45888 32774
rect 45836 32710 45888 32716
rect 45744 32224 45796 32230
rect 45744 32166 45796 32172
rect 45652 31272 45704 31278
rect 45652 31214 45704 31220
rect 45376 29640 45428 29646
rect 45376 29582 45428 29588
rect 45560 29640 45612 29646
rect 45560 29582 45612 29588
rect 45388 28422 45416 29582
rect 45376 28416 45428 28422
rect 45376 28358 45428 28364
rect 45388 28218 45416 28358
rect 45376 28212 45428 28218
rect 45376 28154 45428 28160
rect 45284 27056 45336 27062
rect 45284 26998 45336 27004
rect 45112 26948 45186 26976
rect 44732 26852 44784 26858
rect 45158 26840 45186 26948
rect 44732 26794 44784 26800
rect 45112 26812 45186 26840
rect 44744 25838 44772 26794
rect 44824 26376 44876 26382
rect 44824 26318 44876 26324
rect 44836 26042 44864 26318
rect 44824 26036 44876 26042
rect 44824 25978 44876 25984
rect 44732 25832 44784 25838
rect 44732 25774 44784 25780
rect 44824 24064 44876 24070
rect 44824 24006 44876 24012
rect 44640 23180 44692 23186
rect 44640 23122 44692 23128
rect 44456 22568 44508 22574
rect 44456 22510 44508 22516
rect 44548 21888 44600 21894
rect 44548 21830 44600 21836
rect 44560 21554 44588 21830
rect 44548 21548 44600 21554
rect 44548 21490 44600 21496
rect 44640 21412 44692 21418
rect 44640 21354 44692 21360
rect 44652 21146 44680 21354
rect 44640 21140 44692 21146
rect 44640 21082 44692 21088
rect 43996 21072 44048 21078
rect 43996 21014 44048 21020
rect 44008 20534 44036 21014
rect 44364 20936 44416 20942
rect 44364 20878 44416 20884
rect 44376 20602 44404 20878
rect 44732 20800 44784 20806
rect 44732 20742 44784 20748
rect 44364 20596 44416 20602
rect 44364 20538 44416 20544
rect 43996 20528 44048 20534
rect 43996 20470 44048 20476
rect 44744 18329 44772 20742
rect 44836 19922 44864 24006
rect 45112 23662 45140 26812
rect 45296 26790 45324 26998
rect 45284 26784 45336 26790
rect 45204 26744 45284 26772
rect 45204 24449 45232 26744
rect 45284 26726 45336 26732
rect 45560 26308 45612 26314
rect 45560 26250 45612 26256
rect 45376 25832 45428 25838
rect 45376 25774 45428 25780
rect 45468 25832 45520 25838
rect 45468 25774 45520 25780
rect 45284 25288 45336 25294
rect 45284 25230 45336 25236
rect 45190 24440 45246 24449
rect 45296 24410 45324 25230
rect 45190 24375 45246 24384
rect 45284 24404 45336 24410
rect 45284 24346 45336 24352
rect 45388 23730 45416 25774
rect 45480 24993 45508 25774
rect 45572 25294 45600 26250
rect 45560 25288 45612 25294
rect 45560 25230 45612 25236
rect 45466 24984 45522 24993
rect 45572 24954 45600 25230
rect 45466 24919 45522 24928
rect 45560 24948 45612 24954
rect 45480 24834 45508 24919
rect 45560 24890 45612 24896
rect 45480 24806 45600 24834
rect 45468 24404 45520 24410
rect 45468 24346 45520 24352
rect 45376 23724 45428 23730
rect 45376 23666 45428 23672
rect 45100 23656 45152 23662
rect 45100 23598 45152 23604
rect 45008 23180 45060 23186
rect 45008 23122 45060 23128
rect 45020 22438 45048 23122
rect 45008 22432 45060 22438
rect 45008 22374 45060 22380
rect 45020 21321 45048 22374
rect 45112 22001 45140 23598
rect 45480 23322 45508 24346
rect 45468 23316 45520 23322
rect 45468 23258 45520 23264
rect 45192 22500 45244 22506
rect 45192 22442 45244 22448
rect 45098 21992 45154 22001
rect 45098 21927 45154 21936
rect 45006 21312 45062 21321
rect 45006 21247 45062 21256
rect 44824 19916 44876 19922
rect 44824 19858 44876 19864
rect 44836 19514 44864 19858
rect 44824 19508 44876 19514
rect 44824 19450 44876 19456
rect 45008 19168 45060 19174
rect 45008 19110 45060 19116
rect 44916 18760 44968 18766
rect 44916 18702 44968 18708
rect 44928 18358 44956 18702
rect 45020 18426 45048 19110
rect 45112 18986 45140 21927
rect 45204 21418 45232 22442
rect 45376 22160 45428 22166
rect 45376 22102 45428 22108
rect 45284 22024 45336 22030
rect 45284 21966 45336 21972
rect 45296 21690 45324 21966
rect 45284 21684 45336 21690
rect 45284 21626 45336 21632
rect 45192 21412 45244 21418
rect 45192 21354 45244 21360
rect 45204 19242 45232 21354
rect 45388 21350 45416 22102
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45376 21344 45428 21350
rect 45376 21286 45428 21292
rect 45376 21072 45428 21078
rect 45376 21014 45428 21020
rect 45388 20534 45416 21014
rect 45376 20528 45428 20534
rect 45376 20470 45428 20476
rect 45284 19780 45336 19786
rect 45284 19722 45336 19728
rect 45192 19236 45244 19242
rect 45192 19178 45244 19184
rect 45112 18958 45232 18986
rect 45100 18896 45152 18902
rect 45100 18838 45152 18844
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 44916 18352 44968 18358
rect 44730 18320 44786 18329
rect 44916 18294 44968 18300
rect 44730 18255 44786 18264
rect 45112 18086 45140 18838
rect 45100 18080 45152 18086
rect 45100 18022 45152 18028
rect 44638 17912 44694 17921
rect 44638 17847 44694 17856
rect 44652 17066 44680 17847
rect 45112 17814 45140 18022
rect 44916 17808 44968 17814
rect 44916 17750 44968 17756
rect 45100 17808 45152 17814
rect 45100 17750 45152 17756
rect 44824 17672 44876 17678
rect 44824 17614 44876 17620
rect 44836 17338 44864 17614
rect 44824 17332 44876 17338
rect 44824 17274 44876 17280
rect 44640 17060 44692 17066
rect 44640 17002 44692 17008
rect 44652 16658 44680 17002
rect 44836 16794 44864 17274
rect 44928 17202 44956 17750
rect 44916 17196 44968 17202
rect 44916 17138 44968 17144
rect 45204 17134 45232 18958
rect 45192 17128 45244 17134
rect 45192 17070 45244 17076
rect 44824 16788 44876 16794
rect 44824 16730 44876 16736
rect 43904 16652 43956 16658
rect 43904 16594 43956 16600
rect 44640 16652 44692 16658
rect 44640 16594 44692 16600
rect 44272 16516 44324 16522
rect 44272 16458 44324 16464
rect 43720 16448 43772 16454
rect 43720 16390 43772 16396
rect 43732 14482 43760 16390
rect 44284 16046 44312 16458
rect 44652 16250 44680 16594
rect 44640 16244 44692 16250
rect 44640 16186 44692 16192
rect 44272 16040 44324 16046
rect 44272 15982 44324 15988
rect 44284 15706 44312 15982
rect 44272 15700 44324 15706
rect 44272 15642 44324 15648
rect 43996 15428 44048 15434
rect 43996 15370 44048 15376
rect 44008 15094 44036 15370
rect 43996 15088 44048 15094
rect 43996 15030 44048 15036
rect 44008 14550 44036 15030
rect 43996 14544 44048 14550
rect 43996 14486 44048 14492
rect 45192 14544 45244 14550
rect 45192 14486 45244 14492
rect 43720 14476 43772 14482
rect 43720 14418 43772 14424
rect 43732 14074 43760 14418
rect 45204 14074 45232 14486
rect 43720 14068 43772 14074
rect 43720 14010 43772 14016
rect 45192 14068 45244 14074
rect 45192 14010 45244 14016
rect 43812 14000 43864 14006
rect 43812 13942 43864 13948
rect 43824 13802 43852 13942
rect 45296 13814 45324 19722
rect 45480 17814 45508 21966
rect 45572 21078 45600 24806
rect 45664 23662 45692 31214
rect 45756 28626 45784 32166
rect 45848 31822 45876 32710
rect 45836 31816 45888 31822
rect 45836 31758 45888 31764
rect 45848 31482 45876 31758
rect 45836 31476 45888 31482
rect 45836 31418 45888 31424
rect 45928 30796 45980 30802
rect 45928 30738 45980 30744
rect 45940 30326 45968 30738
rect 45928 30320 45980 30326
rect 45928 30262 45980 30268
rect 45744 28620 45796 28626
rect 45744 28562 45796 28568
rect 45756 27878 45784 28562
rect 45744 27872 45796 27878
rect 45744 27814 45796 27820
rect 45756 24721 45784 27814
rect 45836 27328 45888 27334
rect 45836 27270 45888 27276
rect 45848 26790 45876 27270
rect 45836 26784 45888 26790
rect 45836 26726 45888 26732
rect 45848 26518 45876 26726
rect 45836 26512 45888 26518
rect 45836 26454 45888 26460
rect 45848 26042 45876 26454
rect 45926 26344 45982 26353
rect 45926 26279 45982 26288
rect 45836 26036 45888 26042
rect 45836 25978 45888 25984
rect 45742 24712 45798 24721
rect 45742 24647 45798 24656
rect 45836 24336 45888 24342
rect 45836 24278 45888 24284
rect 45848 23866 45876 24278
rect 45836 23860 45888 23866
rect 45836 23802 45888 23808
rect 45836 23724 45888 23730
rect 45836 23666 45888 23672
rect 45652 23656 45704 23662
rect 45652 23598 45704 23604
rect 45664 22234 45692 23598
rect 45848 22574 45876 23666
rect 45836 22568 45888 22574
rect 45836 22510 45888 22516
rect 45848 22409 45876 22510
rect 45834 22400 45890 22409
rect 45834 22335 45890 22344
rect 45652 22228 45704 22234
rect 45652 22170 45704 22176
rect 45744 21888 45796 21894
rect 45744 21830 45796 21836
rect 45652 21616 45704 21622
rect 45652 21558 45704 21564
rect 45560 21072 45612 21078
rect 45560 21014 45612 21020
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 45572 18902 45600 20878
rect 45560 18896 45612 18902
rect 45560 18838 45612 18844
rect 45468 17808 45520 17814
rect 45468 17750 45520 17756
rect 45560 16652 45612 16658
rect 45560 16594 45612 16600
rect 45572 16522 45600 16594
rect 45560 16516 45612 16522
rect 45560 16458 45612 16464
rect 45572 16250 45600 16458
rect 45560 16244 45612 16250
rect 45560 16186 45612 16192
rect 45560 14544 45612 14550
rect 45560 14486 45612 14492
rect 43812 13796 43864 13802
rect 43812 13738 43864 13744
rect 44364 13796 44416 13802
rect 44364 13738 44416 13744
rect 45204 13786 45324 13814
rect 43720 13320 43772 13326
rect 43720 13262 43772 13268
rect 43732 12850 43760 13262
rect 43720 12844 43772 12850
rect 43720 12786 43772 12792
rect 43628 12232 43680 12238
rect 43628 12174 43680 12180
rect 43628 12096 43680 12102
rect 43628 12038 43680 12044
rect 43260 11892 43312 11898
rect 43260 11834 43312 11840
rect 43444 11892 43496 11898
rect 43444 11834 43496 11840
rect 43272 11558 43300 11834
rect 43456 11558 43484 11834
rect 43640 11626 43668 12038
rect 43628 11620 43680 11626
rect 43628 11562 43680 11568
rect 43260 11552 43312 11558
rect 43260 11494 43312 11500
rect 43444 11552 43496 11558
rect 43444 11494 43496 11500
rect 43076 10192 43128 10198
rect 43076 10134 43128 10140
rect 43088 9654 43116 10134
rect 43076 9648 43128 9654
rect 43076 9590 43128 9596
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43272 9110 43300 9522
rect 43260 9104 43312 9110
rect 43260 9046 43312 9052
rect 43536 9104 43588 9110
rect 43536 9046 43588 9052
rect 43444 8968 43496 8974
rect 43444 8910 43496 8916
rect 43456 8566 43484 8910
rect 43548 8634 43576 9046
rect 43640 8956 43668 11562
rect 43720 10804 43772 10810
rect 43824 10792 43852 13738
rect 44376 13326 44404 13738
rect 44364 13320 44416 13326
rect 44364 13262 44416 13268
rect 44456 12708 44508 12714
rect 44456 12650 44508 12656
rect 44468 11626 44496 12650
rect 44732 12232 44784 12238
rect 44732 12174 44784 12180
rect 44456 11620 44508 11626
rect 44456 11562 44508 11568
rect 44548 11620 44600 11626
rect 44548 11562 44600 11568
rect 43996 11552 44048 11558
rect 43996 11494 44048 11500
rect 44008 11286 44036 11494
rect 43996 11280 44048 11286
rect 43996 11222 44048 11228
rect 43904 11144 43956 11150
rect 43904 11086 43956 11092
rect 43916 10810 43944 11086
rect 43772 10764 43852 10792
rect 43904 10804 43956 10810
rect 43720 10746 43772 10752
rect 43904 10746 43956 10752
rect 43812 10532 43864 10538
rect 43812 10474 43864 10480
rect 43824 10266 43852 10474
rect 43812 10260 43864 10266
rect 43812 10202 43864 10208
rect 43824 9926 43852 10202
rect 43916 10198 43944 10746
rect 44008 10742 44036 11222
rect 43996 10736 44048 10742
rect 43996 10678 44048 10684
rect 44088 10668 44140 10674
rect 44088 10610 44140 10616
rect 44100 10538 44128 10610
rect 44088 10532 44140 10538
rect 44088 10474 44140 10480
rect 44100 10198 44128 10474
rect 43904 10192 43956 10198
rect 43904 10134 43956 10140
rect 44088 10192 44140 10198
rect 44088 10134 44140 10140
rect 43904 10056 43956 10062
rect 43904 9998 43956 10004
rect 43812 9920 43864 9926
rect 43812 9862 43864 9868
rect 43916 9586 43944 9998
rect 44100 9722 44128 10134
rect 44468 9994 44496 11562
rect 44560 11150 44588 11562
rect 44548 11144 44600 11150
rect 44548 11086 44600 11092
rect 44560 10742 44588 11086
rect 44548 10736 44600 10742
rect 44548 10678 44600 10684
rect 44456 9988 44508 9994
rect 44456 9930 44508 9936
rect 44088 9716 44140 9722
rect 44088 9658 44140 9664
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 44088 9444 44140 9450
rect 44088 9386 44140 9392
rect 44100 9178 44128 9386
rect 44088 9172 44140 9178
rect 44088 9114 44140 9120
rect 43720 8968 43772 8974
rect 43640 8928 43720 8956
rect 43720 8910 43772 8916
rect 43536 8628 43588 8634
rect 43536 8570 43588 8576
rect 43444 8560 43496 8566
rect 43444 8502 43496 8508
rect 43732 8498 43760 8910
rect 43720 8492 43772 8498
rect 43720 8434 43772 8440
rect 44272 8424 44324 8430
rect 44272 8366 44324 8372
rect 43812 8356 43864 8362
rect 43812 8298 43864 8304
rect 43824 7954 43852 8298
rect 44284 8090 44312 8366
rect 44364 8288 44416 8294
rect 44364 8230 44416 8236
rect 44272 8084 44324 8090
rect 44272 8026 44324 8032
rect 43812 7948 43864 7954
rect 43812 7890 43864 7896
rect 43824 7546 43852 7890
rect 43904 7812 43956 7818
rect 43904 7754 43956 7760
rect 43812 7540 43864 7546
rect 43812 7482 43864 7488
rect 43916 7478 43944 7754
rect 44376 7546 44404 8230
rect 44456 7880 44508 7886
rect 44456 7822 44508 7828
rect 44468 7750 44496 7822
rect 44456 7744 44508 7750
rect 44456 7686 44508 7692
rect 44364 7540 44416 7546
rect 44364 7482 44416 7488
rect 43904 7472 43956 7478
rect 43904 7414 43956 7420
rect 44376 7206 44404 7482
rect 44364 7200 44416 7206
rect 44364 7142 44416 7148
rect 42706 7032 42762 7041
rect 42156 6996 42208 7002
rect 42156 6938 42208 6944
rect 42340 6996 42392 7002
rect 42706 6967 42762 6976
rect 42340 6938 42392 6944
rect 42720 6866 42748 6967
rect 44376 6934 44404 7142
rect 43536 6928 43588 6934
rect 43442 6896 43498 6905
rect 42156 6860 42208 6866
rect 42156 6802 42208 6808
rect 42708 6860 42760 6866
rect 43536 6870 43588 6876
rect 44364 6928 44416 6934
rect 44364 6870 44416 6876
rect 43442 6831 43498 6840
rect 42708 6802 42760 6808
rect 42168 6458 42196 6802
rect 43456 6798 43484 6831
rect 43444 6792 43496 6798
rect 43444 6734 43496 6740
rect 42616 6724 42668 6730
rect 42616 6666 42668 6672
rect 42340 6656 42392 6662
rect 42340 6598 42392 6604
rect 42156 6452 42208 6458
rect 42156 6394 42208 6400
rect 41696 6180 41748 6186
rect 41696 6122 41748 6128
rect 41972 6180 42024 6186
rect 41972 6122 42024 6128
rect 41880 5840 41932 5846
rect 41880 5782 41932 5788
rect 41512 5704 41564 5710
rect 41512 5646 41564 5652
rect 41524 5302 41552 5646
rect 41892 5302 41920 5782
rect 40684 5296 40736 5302
rect 40684 5238 40736 5244
rect 40868 5296 40920 5302
rect 40868 5238 40920 5244
rect 41512 5296 41564 5302
rect 41512 5238 41564 5244
rect 41880 5296 41932 5302
rect 41880 5238 41932 5244
rect 40132 5228 40184 5234
rect 40132 5170 40184 5176
rect 40696 5098 40724 5238
rect 40684 5092 40736 5098
rect 40684 5034 40736 5040
rect 41604 5092 41656 5098
rect 41604 5034 41656 5040
rect 39764 4752 39816 4758
rect 39764 4694 39816 4700
rect 39776 4214 39804 4694
rect 41328 4684 41380 4690
rect 41328 4626 41380 4632
rect 40776 4480 40828 4486
rect 40776 4422 40828 4428
rect 39764 4208 39816 4214
rect 39764 4150 39816 4156
rect 40788 4078 40816 4422
rect 41340 4154 41368 4626
rect 41616 4282 41644 5034
rect 41788 4548 41840 4554
rect 41788 4490 41840 4496
rect 41696 4480 41748 4486
rect 41696 4422 41748 4428
rect 41604 4276 41656 4282
rect 41604 4218 41656 4224
rect 41248 4126 41368 4154
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 39764 3528 39816 3534
rect 39764 3470 39816 3476
rect 39776 3058 39804 3470
rect 39960 3126 39988 3606
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 39960 2922 39988 3062
rect 39948 2916 40000 2922
rect 39948 2858 40000 2864
rect 40052 2650 40080 3538
rect 40500 3052 40552 3058
rect 40500 2994 40552 3000
rect 40512 2650 40540 2994
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 40788 2514 40816 4014
rect 41248 3942 41276 4126
rect 41616 3942 41644 4218
rect 41052 3936 41104 3942
rect 41052 3878 41104 3884
rect 41236 3936 41288 3942
rect 41236 3878 41288 3884
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 41064 2650 41092 3878
rect 41248 3194 41276 3878
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 41708 3058 41736 4422
rect 41800 3670 41828 4490
rect 41880 4480 41932 4486
rect 41880 4422 41932 4428
rect 41892 4010 41920 4422
rect 41880 4004 41932 4010
rect 41880 3946 41932 3952
rect 41788 3664 41840 3670
rect 41788 3606 41840 3612
rect 41696 3052 41748 3058
rect 41696 2994 41748 3000
rect 41052 2644 41104 2650
rect 41052 2586 41104 2592
rect 40776 2508 40828 2514
rect 40776 2450 40828 2456
rect 41892 2378 41920 3946
rect 41984 3670 42012 6122
rect 42352 5370 42380 6598
rect 42628 6458 42656 6666
rect 43456 6458 43484 6734
rect 42616 6452 42668 6458
rect 42616 6394 42668 6400
rect 43444 6452 43496 6458
rect 43444 6394 43496 6400
rect 43548 6186 43576 6870
rect 43904 6792 43956 6798
rect 43904 6734 43956 6740
rect 43916 6322 43944 6734
rect 44088 6656 44140 6662
rect 44088 6598 44140 6604
rect 43904 6316 43956 6322
rect 43904 6258 43956 6264
rect 43444 6180 43496 6186
rect 43444 6122 43496 6128
rect 43536 6180 43588 6186
rect 43536 6122 43588 6128
rect 43456 5846 43484 6122
rect 43444 5840 43496 5846
rect 43444 5782 43496 5788
rect 43076 5704 43128 5710
rect 43076 5646 43128 5652
rect 42340 5364 42392 5370
rect 42340 5306 42392 5312
rect 43088 4826 43116 5646
rect 43456 5370 43484 5782
rect 43444 5364 43496 5370
rect 43444 5306 43496 5312
rect 43076 4820 43128 4826
rect 43076 4762 43128 4768
rect 43456 4758 43484 5306
rect 43548 5098 43576 6122
rect 43916 5914 43944 6258
rect 43904 5908 43956 5914
rect 43904 5850 43956 5856
rect 44100 5710 44128 6598
rect 44088 5704 44140 5710
rect 44088 5646 44140 5652
rect 43812 5568 43864 5574
rect 43812 5510 43864 5516
rect 43824 5234 43852 5510
rect 43812 5228 43864 5234
rect 43812 5170 43864 5176
rect 43536 5092 43588 5098
rect 43536 5034 43588 5040
rect 43444 4752 43496 4758
rect 43444 4694 43496 4700
rect 42800 4684 42852 4690
rect 42800 4626 42852 4632
rect 42616 4140 42668 4146
rect 42616 4082 42668 4088
rect 42524 4004 42576 4010
rect 42524 3946 42576 3952
rect 42064 3936 42116 3942
rect 42064 3878 42116 3884
rect 41972 3664 42024 3670
rect 41972 3606 42024 3612
rect 41984 3194 42012 3606
rect 42076 3194 42104 3878
rect 42536 3670 42564 3946
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 42628 3602 42656 4082
rect 42812 3942 42840 4626
rect 43456 4282 43484 4694
rect 43444 4276 43496 4282
rect 43444 4218 43496 4224
rect 43456 3992 43484 4218
rect 43548 4154 43576 5034
rect 43720 4616 43772 4622
rect 43720 4558 43772 4564
rect 43548 4126 43668 4154
rect 43536 4004 43588 4010
rect 43456 3964 43536 3992
rect 43536 3946 43588 3952
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42812 3738 42840 3878
rect 42800 3732 42852 3738
rect 42800 3674 42852 3680
rect 43640 3670 43668 4126
rect 43732 4049 43760 4558
rect 43824 4554 43852 5170
rect 43812 4548 43864 4554
rect 43812 4490 43864 4496
rect 43996 4208 44048 4214
rect 43996 4150 44048 4156
rect 43718 4040 43774 4049
rect 43718 3975 43774 3984
rect 43904 4004 43956 4010
rect 43732 3738 43760 3975
rect 43904 3946 43956 3952
rect 43916 3913 43944 3946
rect 43902 3904 43958 3913
rect 43902 3839 43958 3848
rect 43902 3768 43958 3777
rect 43720 3732 43772 3738
rect 43902 3703 43958 3712
rect 43720 3674 43772 3680
rect 43628 3664 43680 3670
rect 43628 3606 43680 3612
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 41972 3188 42024 3194
rect 41972 3130 42024 3136
rect 42064 3188 42116 3194
rect 42064 3130 42116 3136
rect 42432 3188 42484 3194
rect 42432 3130 42484 3136
rect 41984 2582 42012 3130
rect 42340 3052 42392 3058
rect 42340 2994 42392 3000
rect 42064 2984 42116 2990
rect 42064 2926 42116 2932
rect 41972 2576 42024 2582
rect 41972 2518 42024 2524
rect 42076 2446 42104 2926
rect 42064 2440 42116 2446
rect 42064 2382 42116 2388
rect 41880 2372 41932 2378
rect 41880 2314 41932 2320
rect 42352 2310 42380 2994
rect 42444 2922 42472 3130
rect 42628 3058 42656 3538
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42432 2916 42484 2922
rect 42432 2858 42484 2864
rect 43456 2582 43484 3470
rect 43640 3194 43668 3606
rect 43628 3188 43680 3194
rect 43628 3130 43680 3136
rect 43640 2854 43668 3130
rect 43916 3058 43944 3703
rect 44008 3466 44036 4150
rect 43996 3460 44048 3466
rect 43996 3402 44048 3408
rect 44100 3058 44128 5646
rect 44468 5098 44496 7686
rect 44548 7268 44600 7274
rect 44548 7210 44600 7216
rect 44560 6662 44588 7210
rect 44548 6656 44600 6662
rect 44548 6598 44600 6604
rect 44744 6254 44772 12174
rect 45204 11218 45232 13786
rect 45468 13728 45520 13734
rect 45572 13716 45600 14486
rect 45520 13688 45600 13716
rect 45468 13670 45520 13676
rect 45480 13462 45508 13670
rect 45376 13456 45428 13462
rect 45376 13398 45428 13404
rect 45468 13456 45520 13462
rect 45468 13398 45520 13404
rect 45284 13320 45336 13326
rect 45284 13262 45336 13268
rect 45296 12442 45324 13262
rect 45388 12646 45416 13398
rect 45376 12640 45428 12646
rect 45376 12582 45428 12588
rect 45284 12436 45336 12442
rect 45284 12378 45336 12384
rect 45480 12374 45508 13398
rect 45468 12368 45520 12374
rect 45468 12310 45520 12316
rect 45376 12232 45428 12238
rect 45376 12174 45428 12180
rect 45388 11626 45416 12174
rect 45480 11898 45508 12310
rect 45468 11892 45520 11898
rect 45468 11834 45520 11840
rect 45376 11620 45428 11626
rect 45376 11562 45428 11568
rect 45192 11212 45244 11218
rect 45192 11154 45244 11160
rect 45204 10810 45232 11154
rect 45192 10804 45244 10810
rect 45192 10746 45244 10752
rect 45664 8401 45692 21558
rect 45756 21078 45784 21830
rect 45744 21072 45796 21078
rect 45744 21014 45796 21020
rect 45836 21072 45888 21078
rect 45836 21014 45888 21020
rect 45756 20602 45784 21014
rect 45848 20602 45876 21014
rect 45744 20596 45796 20602
rect 45744 20538 45796 20544
rect 45836 20596 45888 20602
rect 45836 20538 45888 20544
rect 45848 20482 45876 20538
rect 45756 20454 45876 20482
rect 45756 20262 45784 20454
rect 45744 20256 45796 20262
rect 45744 20198 45796 20204
rect 45834 20224 45890 20233
rect 45756 20058 45784 20198
rect 45834 20159 45890 20168
rect 45744 20052 45796 20058
rect 45744 19994 45796 20000
rect 45848 19922 45876 20159
rect 45836 19916 45888 19922
rect 45836 19858 45888 19864
rect 45848 19514 45876 19858
rect 45836 19508 45888 19514
rect 45836 19450 45888 19456
rect 45940 18222 45968 26279
rect 45928 18216 45980 18222
rect 45928 18158 45980 18164
rect 45836 15496 45888 15502
rect 45836 15438 45888 15444
rect 45848 14550 45876 15438
rect 45836 14544 45888 14550
rect 45836 14486 45888 14492
rect 45848 13258 45876 14486
rect 46032 14482 46060 33798
rect 46124 31929 46152 35391
rect 46940 35148 46992 35154
rect 46940 35090 46992 35096
rect 46952 34406 46980 35090
rect 46940 34400 46992 34406
rect 46940 34342 46992 34348
rect 46952 33522 46980 34342
rect 46940 33516 46992 33522
rect 46940 33458 46992 33464
rect 49528 33425 49556 39063
rect 49514 33416 49570 33425
rect 49514 33351 49570 33360
rect 46664 32428 46716 32434
rect 46664 32370 46716 32376
rect 46676 32026 46704 32370
rect 47582 32328 47638 32337
rect 46848 32292 46900 32298
rect 47582 32263 47638 32272
rect 46848 32234 46900 32240
rect 46664 32020 46716 32026
rect 46664 31962 46716 31968
rect 46110 31920 46166 31929
rect 46110 31855 46166 31864
rect 46388 31884 46440 31890
rect 46124 31278 46152 31855
rect 46388 31826 46440 31832
rect 46112 31272 46164 31278
rect 46112 31214 46164 31220
rect 46400 31210 46428 31826
rect 46388 31204 46440 31210
rect 46388 31146 46440 31152
rect 46296 31136 46348 31142
rect 46296 31078 46348 31084
rect 46308 29617 46336 31078
rect 46860 30870 46888 32234
rect 46848 30864 46900 30870
rect 46848 30806 46900 30812
rect 47032 30592 47084 30598
rect 47032 30534 47084 30540
rect 46940 30252 46992 30258
rect 46940 30194 46992 30200
rect 46388 30048 46440 30054
rect 46388 29990 46440 29996
rect 46294 29608 46350 29617
rect 46294 29543 46350 29552
rect 46400 28529 46428 29990
rect 46952 29714 46980 30194
rect 47044 30190 47072 30534
rect 47596 30394 47624 32263
rect 47584 30388 47636 30394
rect 47584 30330 47636 30336
rect 47032 30184 47084 30190
rect 47032 30126 47084 30132
rect 46940 29708 46992 29714
rect 46940 29650 46992 29656
rect 46848 29504 46900 29510
rect 46848 29446 46900 29452
rect 46860 28801 46888 29446
rect 46952 29238 46980 29650
rect 47044 29306 47072 30126
rect 49514 29744 49570 29753
rect 47216 29708 47268 29714
rect 49514 29679 49570 29688
rect 47216 29650 47268 29656
rect 47032 29300 47084 29306
rect 47032 29242 47084 29248
rect 46940 29232 46992 29238
rect 46940 29174 46992 29180
rect 47228 29102 47256 29650
rect 47216 29096 47268 29102
rect 47216 29038 47268 29044
rect 46846 28792 46902 28801
rect 46846 28727 46902 28736
rect 47124 28620 47176 28626
rect 47124 28562 47176 28568
rect 46386 28520 46442 28529
rect 46386 28455 46442 28464
rect 46204 28416 46256 28422
rect 46204 28358 46256 28364
rect 46756 28416 46808 28422
rect 46756 28358 46808 28364
rect 46216 28082 46244 28358
rect 46204 28076 46256 28082
rect 46204 28018 46256 28024
rect 46480 28076 46532 28082
rect 46480 28018 46532 28024
rect 46204 27940 46256 27946
rect 46204 27882 46256 27888
rect 46216 27606 46244 27882
rect 46492 27878 46520 28018
rect 46480 27872 46532 27878
rect 46768 27849 46796 28358
rect 47136 27878 47164 28562
rect 47228 28422 47256 29038
rect 47216 28416 47268 28422
rect 47216 28358 47268 28364
rect 48228 28416 48280 28422
rect 48228 28358 48280 28364
rect 47124 27872 47176 27878
rect 46480 27814 46532 27820
rect 46754 27840 46810 27849
rect 46204 27600 46256 27606
rect 46204 27542 46256 27548
rect 46388 27464 46440 27470
rect 46388 27406 46440 27412
rect 46400 27130 46428 27406
rect 46388 27124 46440 27130
rect 46388 27066 46440 27072
rect 46204 26852 46256 26858
rect 46204 26794 46256 26800
rect 46216 26586 46244 26794
rect 46204 26580 46256 26586
rect 46204 26522 46256 26528
rect 46216 26042 46244 26522
rect 46204 26036 46256 26042
rect 46204 25978 46256 25984
rect 46296 25424 46348 25430
rect 46296 25366 46348 25372
rect 46204 25288 46256 25294
rect 46204 25230 46256 25236
rect 46216 24818 46244 25230
rect 46308 25158 46336 25366
rect 46296 25152 46348 25158
rect 46296 25094 46348 25100
rect 46204 24812 46256 24818
rect 46204 24754 46256 24760
rect 46308 24682 46336 25094
rect 46386 24712 46442 24721
rect 46296 24676 46348 24682
rect 46386 24647 46442 24656
rect 46296 24618 46348 24624
rect 46308 24342 46336 24618
rect 46296 24336 46348 24342
rect 46296 24278 46348 24284
rect 46112 24200 46164 24206
rect 46112 24142 46164 24148
rect 46124 23798 46152 24142
rect 46112 23792 46164 23798
rect 46112 23734 46164 23740
rect 46124 23322 46152 23734
rect 46400 23474 46428 24647
rect 46492 24206 46520 27814
rect 47124 27814 47176 27820
rect 46754 27775 46810 27784
rect 46756 27056 46808 27062
rect 46756 26998 46808 27004
rect 46768 25786 46796 26998
rect 47136 26897 47164 27814
rect 47122 26888 47178 26897
rect 47122 26823 47178 26832
rect 46848 26580 46900 26586
rect 46848 26522 46900 26528
rect 46584 25758 46796 25786
rect 46584 25702 46612 25758
rect 46572 25696 46624 25702
rect 46572 25638 46624 25644
rect 46664 25696 46716 25702
rect 46664 25638 46716 25644
rect 46676 25401 46704 25638
rect 46662 25392 46718 25401
rect 46662 25327 46718 25336
rect 46480 24200 46532 24206
rect 46480 24142 46532 24148
rect 46400 23446 46520 23474
rect 46112 23316 46164 23322
rect 46112 23258 46164 23264
rect 46492 22098 46520 23446
rect 46480 22092 46532 22098
rect 46480 22034 46532 22040
rect 46676 21350 46704 25327
rect 46768 24886 46796 25758
rect 46756 24880 46808 24886
rect 46756 24822 46808 24828
rect 46756 22092 46808 22098
rect 46756 22034 46808 22040
rect 46768 21622 46796 22034
rect 46756 21616 46808 21622
rect 46756 21558 46808 21564
rect 46664 21344 46716 21350
rect 46664 21286 46716 21292
rect 46204 20324 46256 20330
rect 46204 20266 46256 20272
rect 46216 20058 46244 20266
rect 46204 20052 46256 20058
rect 46204 19994 46256 20000
rect 46480 18896 46532 18902
rect 46480 18838 46532 18844
rect 46572 18896 46624 18902
rect 46572 18838 46624 18844
rect 46204 18080 46256 18086
rect 46204 18022 46256 18028
rect 46216 17882 46244 18022
rect 46492 17882 46520 18838
rect 46584 18086 46612 18838
rect 46572 18080 46624 18086
rect 46572 18022 46624 18028
rect 46676 17898 46704 21286
rect 46860 20806 46888 26522
rect 47124 26444 47176 26450
rect 47124 26386 47176 26392
rect 47032 25832 47084 25838
rect 47032 25774 47084 25780
rect 47044 24070 47072 25774
rect 47136 25702 47164 26386
rect 47124 25696 47176 25702
rect 47124 25638 47176 25644
rect 47582 24440 47638 24449
rect 47582 24375 47638 24384
rect 47032 24064 47084 24070
rect 47032 24006 47084 24012
rect 47596 21486 47624 24375
rect 46940 21480 46992 21486
rect 46940 21422 46992 21428
rect 47584 21480 47636 21486
rect 47584 21422 47636 21428
rect 46848 20800 46900 20806
rect 46848 20742 46900 20748
rect 46848 20324 46900 20330
rect 46848 20266 46900 20272
rect 46756 19236 46808 19242
rect 46756 19178 46808 19184
rect 46768 18766 46796 19178
rect 46756 18760 46808 18766
rect 46756 18702 46808 18708
rect 46860 18290 46888 20266
rect 46848 18284 46900 18290
rect 46848 18226 46900 18232
rect 46952 18170 46980 21422
rect 47032 20528 47084 20534
rect 47032 20470 47084 20476
rect 46204 17876 46256 17882
rect 46204 17818 46256 17824
rect 46480 17876 46532 17882
rect 46480 17818 46532 17824
rect 46584 17870 46704 17898
rect 46768 18142 46980 18170
rect 46388 16992 46440 16998
rect 46388 16934 46440 16940
rect 46296 16448 46348 16454
rect 46296 16390 46348 16396
rect 46112 15972 46164 15978
rect 46112 15914 46164 15920
rect 46124 15638 46152 15914
rect 46112 15632 46164 15638
rect 46112 15574 46164 15580
rect 46124 15162 46152 15574
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 46112 15156 46164 15162
rect 46112 15098 46164 15104
rect 46216 15026 46244 15302
rect 46204 15020 46256 15026
rect 46204 14962 46256 14968
rect 46020 14476 46072 14482
rect 46020 14418 46072 14424
rect 45836 13252 45888 13258
rect 45836 13194 45888 13200
rect 46216 12850 46244 14962
rect 46308 14890 46336 16390
rect 46400 16046 46428 16934
rect 46388 16040 46440 16046
rect 46388 15982 46440 15988
rect 46480 15496 46532 15502
rect 46480 15438 46532 15444
rect 46492 15026 46520 15438
rect 46480 15020 46532 15026
rect 46480 14962 46532 14968
rect 46296 14884 46348 14890
rect 46296 14826 46348 14832
rect 46308 14618 46336 14826
rect 46296 14612 46348 14618
rect 46296 14554 46348 14560
rect 46584 13814 46612 17870
rect 46768 13814 46796 18142
rect 46848 14476 46900 14482
rect 46848 14418 46900 14424
rect 46860 14074 46888 14418
rect 46940 14272 46992 14278
rect 46940 14214 46992 14220
rect 46848 14068 46900 14074
rect 46848 14010 46900 14016
rect 46860 13870 46888 14010
rect 46492 13786 46612 13814
rect 46676 13786 46796 13814
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 46296 13184 46348 13190
rect 46296 13126 46348 13132
rect 46020 12844 46072 12850
rect 46020 12786 46072 12792
rect 46204 12844 46256 12850
rect 46204 12786 46256 12792
rect 46032 12374 46060 12786
rect 46204 12708 46256 12714
rect 46308 12696 46336 13126
rect 46256 12668 46336 12696
rect 46204 12650 46256 12656
rect 46020 12368 46072 12374
rect 46020 12310 46072 12316
rect 46020 11008 46072 11014
rect 46020 10950 46072 10956
rect 46032 10130 46060 10950
rect 46112 10532 46164 10538
rect 46112 10474 46164 10480
rect 46020 10124 46072 10130
rect 46020 10066 46072 10072
rect 45928 10056 45980 10062
rect 45928 9998 45980 10004
rect 45940 9722 45968 9998
rect 45928 9716 45980 9722
rect 45928 9658 45980 9664
rect 45940 9382 45968 9658
rect 46032 9654 46060 10066
rect 46020 9648 46072 9654
rect 46020 9590 46072 9596
rect 45928 9376 45980 9382
rect 45928 9318 45980 9324
rect 46124 9110 46152 10474
rect 46388 9580 46440 9586
rect 46388 9522 46440 9528
rect 46112 9104 46164 9110
rect 46112 9046 46164 9052
rect 45744 8968 45796 8974
rect 45744 8910 45796 8916
rect 46020 8968 46072 8974
rect 46020 8910 46072 8916
rect 45756 8634 45784 8910
rect 45928 8832 45980 8838
rect 45928 8774 45980 8780
rect 45744 8628 45796 8634
rect 45744 8570 45796 8576
rect 45650 8392 45706 8401
rect 45650 8327 45706 8336
rect 45756 8022 45784 8570
rect 45008 8016 45060 8022
rect 45008 7958 45060 7964
rect 45744 8016 45796 8022
rect 45744 7958 45796 7964
rect 45020 7546 45048 7958
rect 45008 7540 45060 7546
rect 45008 7482 45060 7488
rect 45756 7410 45784 7958
rect 45940 7954 45968 8774
rect 46032 8537 46060 8910
rect 46018 8528 46074 8537
rect 46124 8498 46152 9046
rect 46296 8560 46348 8566
rect 46296 8502 46348 8508
rect 46018 8463 46074 8472
rect 46112 8492 46164 8498
rect 46112 8434 46164 8440
rect 46204 8424 46256 8430
rect 46204 8366 46256 8372
rect 46112 8356 46164 8362
rect 46112 8298 46164 8304
rect 45928 7948 45980 7954
rect 45928 7890 45980 7896
rect 46124 7546 46152 8298
rect 46216 8022 46244 8366
rect 46308 8090 46336 8502
rect 46296 8084 46348 8090
rect 46296 8026 46348 8032
rect 46204 8016 46256 8022
rect 46204 7958 46256 7964
rect 46216 7818 46244 7958
rect 46204 7812 46256 7818
rect 46204 7754 46256 7760
rect 46112 7540 46164 7546
rect 46112 7482 46164 7488
rect 45744 7404 45796 7410
rect 45744 7346 45796 7352
rect 46124 7206 46152 7482
rect 46400 7410 46428 9522
rect 46388 7404 46440 7410
rect 46388 7346 46440 7352
rect 46204 7268 46256 7274
rect 46204 7210 46256 7216
rect 46112 7200 46164 7206
rect 46112 7142 46164 7148
rect 45192 6928 45244 6934
rect 45192 6870 45244 6876
rect 45204 6458 45232 6870
rect 46216 6866 46244 7210
rect 46294 7032 46350 7041
rect 46294 6967 46350 6976
rect 46308 6866 46336 6967
rect 46400 6934 46428 7346
rect 46388 6928 46440 6934
rect 46388 6870 46440 6876
rect 46204 6860 46256 6866
rect 46204 6802 46256 6808
rect 46296 6860 46348 6866
rect 46296 6802 46348 6808
rect 45192 6452 45244 6458
rect 45192 6394 45244 6400
rect 44732 6248 44784 6254
rect 44732 6190 44784 6196
rect 46112 6248 46164 6254
rect 46112 6190 46164 6196
rect 44744 6118 44772 6190
rect 44732 6112 44784 6118
rect 44732 6054 44784 6060
rect 45376 6112 45428 6118
rect 45376 6054 45428 6060
rect 45008 5772 45060 5778
rect 45008 5714 45060 5720
rect 45020 5370 45048 5714
rect 45008 5364 45060 5370
rect 45008 5306 45060 5312
rect 44456 5092 44508 5098
rect 44456 5034 44508 5040
rect 44468 4758 44496 5034
rect 45020 4826 45048 5306
rect 45008 4820 45060 4826
rect 45008 4762 45060 4768
rect 44456 4752 44508 4758
rect 44456 4694 44508 4700
rect 45388 4690 45416 6054
rect 46124 5914 46152 6190
rect 46112 5908 46164 5914
rect 46112 5850 46164 5856
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 45388 4214 45416 4626
rect 46216 4282 46244 6802
rect 46308 6458 46336 6802
rect 46296 6452 46348 6458
rect 46296 6394 46348 6400
rect 46204 4276 46256 4282
rect 46204 4218 46256 4224
rect 45376 4208 45428 4214
rect 45376 4150 45428 4156
rect 45744 4072 45796 4078
rect 45744 4014 45796 4020
rect 45756 3641 45784 4014
rect 45742 3632 45798 3641
rect 45742 3567 45798 3576
rect 43904 3052 43956 3058
rect 43904 2994 43956 3000
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 43628 2848 43680 2854
rect 43628 2790 43680 2796
rect 43444 2576 43496 2582
rect 43444 2518 43496 2524
rect 42340 2304 42392 2310
rect 42340 2246 42392 2252
rect 46492 1873 46520 13786
rect 46572 13728 46624 13734
rect 46572 13670 46624 13676
rect 46584 12306 46612 13670
rect 46572 12300 46624 12306
rect 46572 12242 46624 12248
rect 46584 11898 46612 12242
rect 46572 11892 46624 11898
rect 46572 11834 46624 11840
rect 46676 5273 46704 13786
rect 46952 13394 46980 14214
rect 46940 13388 46992 13394
rect 46940 13330 46992 13336
rect 46848 12708 46900 12714
rect 46848 12650 46900 12656
rect 46860 12374 46888 12650
rect 46848 12368 46900 12374
rect 46848 12310 46900 12316
rect 47044 11529 47072 20470
rect 47308 16720 47360 16726
rect 47308 16662 47360 16668
rect 47216 16652 47268 16658
rect 47216 16594 47268 16600
rect 47228 16182 47256 16594
rect 47216 16176 47268 16182
rect 47216 16118 47268 16124
rect 47320 15570 47348 16662
rect 47308 15564 47360 15570
rect 47308 15506 47360 15512
rect 47320 15162 47348 15506
rect 47308 15156 47360 15162
rect 47308 15098 47360 15104
rect 48240 14657 48268 28358
rect 49528 26586 49556 29679
rect 49516 26580 49568 26586
rect 49516 26522 49568 26528
rect 49514 20360 49570 20369
rect 49514 20295 49570 20304
rect 49528 19417 49556 20295
rect 49514 19408 49570 19417
rect 49514 19343 49570 19352
rect 48226 14648 48282 14657
rect 48226 14583 48282 14592
rect 47124 13388 47176 13394
rect 47124 13330 47176 13336
rect 47136 12986 47164 13330
rect 47124 12980 47176 12986
rect 47124 12922 47176 12928
rect 47030 11520 47086 11529
rect 47030 11455 47086 11464
rect 47492 10804 47544 10810
rect 47492 10746 47544 10752
rect 46756 10600 46808 10606
rect 46756 10542 46808 10548
rect 46768 10266 46796 10542
rect 46756 10260 46808 10266
rect 46756 10202 46808 10208
rect 47504 10130 47532 10746
rect 47492 10124 47544 10130
rect 47492 10066 47544 10072
rect 47504 9722 47532 10066
rect 47492 9716 47544 9722
rect 47492 9658 47544 9664
rect 46848 9444 46900 9450
rect 46848 9386 46900 9392
rect 46860 8974 46888 9386
rect 47216 9036 47268 9042
rect 47216 8978 47268 8984
rect 46848 8968 46900 8974
rect 46848 8910 46900 8916
rect 47228 8294 47256 8978
rect 47492 8900 47544 8906
rect 47492 8842 47544 8848
rect 47216 8288 47268 8294
rect 47216 8230 47268 8236
rect 47124 7948 47176 7954
rect 47124 7890 47176 7896
rect 47136 7546 47164 7890
rect 47228 7857 47256 8230
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47214 7848 47270 7857
rect 47214 7783 47270 7792
rect 47124 7540 47176 7546
rect 47124 7482 47176 7488
rect 47412 7478 47440 7890
rect 47504 7886 47532 8842
rect 47492 7880 47544 7886
rect 47492 7822 47544 7828
rect 47400 7472 47452 7478
rect 47400 7414 47452 7420
rect 46662 5264 46718 5273
rect 46662 5199 46718 5208
rect 46478 1864 46534 1873
rect 46478 1799 46534 1808
rect 39118 54 39252 82
rect 24858 0 24914 54
rect 32034 0 32090 54
rect 39118 0 39174 54
rect 46294 0 46350 480
<< via2 >>
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 22282 45328 22338 45384
rect 6090 44104 6146 44160
rect 19062 44104 19118 44160
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 14922 41520 14978 41576
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 12714 29688 12770 29744
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 15934 40568 15990 40624
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19246 43696 19302 43752
rect 19062 42880 19118 42936
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 17498 35572 17500 35592
rect 17500 35572 17552 35592
rect 17552 35572 17554 35592
rect 17498 35536 17554 35572
rect 18602 42064 18658 42120
rect 18602 34720 18658 34776
rect 17222 32816 17278 32872
rect 15842 31864 15898 31920
rect 14370 28600 14426 28656
rect 13542 25744 13598 25800
rect 14370 26016 14426 26072
rect 14186 25200 14242 25256
rect 14278 25064 14334 25120
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 14094 23704 14150 23760
rect 14646 23976 14702 24032
rect 14278 23568 14334 23624
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 16118 26968 16174 27024
rect 15750 25880 15806 25936
rect 18510 34040 18566 34096
rect 19430 42880 19486 42936
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 18970 40432 19026 40488
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19062 33632 19118 33688
rect 18970 33224 19026 33280
rect 18234 31864 18290 31920
rect 18970 33088 19026 33144
rect 17222 26832 17278 26888
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 3790 1944 3846 2000
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19430 31456 19486 31512
rect 19246 28464 19302 28520
rect 17590 23840 17646 23896
rect 16486 21392 16542 21448
rect 17222 22616 17278 22672
rect 22650 35264 22706 35320
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19890 28328 19946 28384
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19062 24248 19118 24304
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 20442 23704 20498 23760
rect 20626 29688 20682 29744
rect 19246 21664 19302 21720
rect 20902 28736 20958 28792
rect 21362 32952 21418 33008
rect 21270 23568 21326 23624
rect 20810 21392 20866 21448
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 18142 16496 18198 16552
rect 17958 13796 18014 13832
rect 17958 13776 17960 13796
rect 17960 13776 18012 13796
rect 18012 13776 18014 13796
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 13818 8880 13874 8936
rect 17130 1944 17186 2000
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19062 13640 19118 13696
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 20074 16496 20130 16552
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19246 13776 19302 13832
rect 19292 13640 19348 13696
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19430 13368 19486 13424
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 21546 22752 21602 22808
rect 23570 34720 23626 34776
rect 22834 34484 22836 34504
rect 22836 34484 22888 34504
rect 22888 34484 22890 34504
rect 22834 34448 22890 34484
rect 22742 32816 22798 32872
rect 24490 40704 24546 40760
rect 24490 40568 24546 40624
rect 24674 40704 24730 40760
rect 28446 45328 28502 45384
rect 27066 43696 27122 43752
rect 26790 42608 26846 42664
rect 26790 42064 26846 42120
rect 26514 40568 26570 40624
rect 26514 40296 26570 40352
rect 23754 32952 23810 33008
rect 22742 30232 22798 30288
rect 23478 28464 23534 28520
rect 22834 25744 22890 25800
rect 23662 23976 23718 24032
rect 23938 25880 23994 25936
rect 23662 21800 23718 21856
rect 23110 19252 23112 19272
rect 23112 19252 23164 19272
rect 23164 19252 23166 19272
rect 23110 19216 23166 19252
rect 23386 19080 23442 19136
rect 23110 16360 23166 16416
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 21822 10240 21878 10296
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19982 8472 20038 8528
rect 21454 8880 21510 8936
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 20534 5616 20590 5672
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 23754 19216 23810 19272
rect 23938 19216 23994 19272
rect 23754 9152 23810 9208
rect 24122 27784 24178 27840
rect 24858 26832 24914 26888
rect 24122 21392 24178 21448
rect 25042 26016 25098 26072
rect 24950 25744 25006 25800
rect 25594 34040 25650 34096
rect 27894 38256 27950 38312
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 28814 40568 28870 40624
rect 29826 40432 29882 40488
rect 26882 35672 26938 35728
rect 24858 22752 24914 22808
rect 25042 22616 25098 22672
rect 26054 33632 26110 33688
rect 28078 35536 28134 35592
rect 28262 35264 28318 35320
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 32954 43832 33010 43888
rect 29734 35264 29790 35320
rect 28446 34448 28502 34504
rect 22282 4800 22338 4856
rect 24858 9424 24914 9480
rect 24398 3712 24454 3768
rect 22098 3032 22154 3088
rect 26422 26968 26478 27024
rect 26330 24248 26386 24304
rect 28630 30912 28686 30968
rect 27342 23840 27398 23896
rect 27434 23296 27490 23352
rect 27342 23160 27398 23216
rect 27894 25472 27950 25528
rect 28722 25880 28778 25936
rect 29734 28736 29790 28792
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34610 42608 34666 42664
rect 32310 40976 32366 41032
rect 32402 40568 32458 40624
rect 34150 42064 34206 42120
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 36266 45328 36322 45384
rect 34150 40704 34206 40760
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34242 40296 34298 40352
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 33414 38256 33470 38312
rect 31482 32136 31538 32192
rect 31850 32544 31906 32600
rect 32586 32952 32642 33008
rect 30286 27784 30342 27840
rect 31850 29008 31906 29064
rect 28538 22888 28594 22944
rect 28538 21936 28594 21992
rect 30194 24384 30250 24440
rect 30838 25200 30894 25256
rect 30746 21800 30802 21856
rect 27986 19352 28042 19408
rect 26330 12688 26386 12744
rect 27894 11600 27950 11656
rect 28630 10512 28686 10568
rect 27250 5616 27306 5672
rect 31206 23160 31262 23216
rect 31022 22752 31078 22808
rect 31390 22344 31446 22400
rect 31298 19080 31354 19136
rect 30930 16360 30986 16416
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 35806 38664 35862 38720
rect 33782 35672 33838 35728
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 33414 34448 33470 34504
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34610 33380 34666 33416
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 35622 35164 35624 35184
rect 35624 35164 35676 35184
rect 35676 35164 35678 35184
rect 35622 35128 35678 35164
rect 37830 44240 37886 44296
rect 34610 33360 34612 33380
rect 34612 33360 34664 33380
rect 34664 33360 34666 33380
rect 35346 33088 35402 33144
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34794 32544 34850 32600
rect 32218 30232 32274 30288
rect 32862 28600 32918 28656
rect 32034 23296 32090 23352
rect 32310 20168 32366 20224
rect 32586 23568 32642 23624
rect 32862 23568 32918 23624
rect 31206 16496 31262 16552
rect 32770 19080 32826 19136
rect 32034 15000 32090 15056
rect 35070 31864 35126 31920
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 33598 26832 33654 26888
rect 34242 28600 34298 28656
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 36818 34584 36874 34640
rect 36266 32136 36322 32192
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 33598 25880 33654 25936
rect 33874 25472 33930 25528
rect 33690 25336 33746 25392
rect 34242 24520 34298 24576
rect 32954 18808 33010 18864
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34794 25744 34850 25800
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 35346 24384 35402 24440
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 36358 29008 36414 29064
rect 36082 28464 36138 28520
rect 36174 24928 36230 24984
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 35990 21936 36046 21992
rect 37094 28736 37150 28792
rect 37278 24656 37334 24712
rect 36174 19352 36230 19408
rect 36358 19352 36414 19408
rect 34518 18808 34574 18864
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 33874 13776 33930 13832
rect 33874 12688 33930 12744
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35806 18264 35862 18320
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 49514 48456 49570 48512
rect 39762 42064 39818 42120
rect 39486 40568 39542 40624
rect 37554 30232 37610 30288
rect 37462 29552 37518 29608
rect 37830 34448 37886 34504
rect 38198 33088 38254 33144
rect 41878 43832 41934 43888
rect 42522 40976 42578 41032
rect 38474 26832 38530 26888
rect 37830 25356 37886 25392
rect 37830 25336 37832 25356
rect 37832 25336 37884 25356
rect 37884 25336 37886 25356
rect 37738 21256 37794 21312
rect 37370 17856 37426 17912
rect 35806 16904 35862 16960
rect 38658 23604 38660 23624
rect 38660 23604 38712 23624
rect 38712 23604 38714 23624
rect 38658 23568 38714 23604
rect 40314 30912 40370 30968
rect 44914 44784 44970 44840
rect 43350 40976 43406 41032
rect 43810 38664 43866 38720
rect 42062 31048 42118 31104
rect 44822 44240 44878 44296
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 36358 13776 36414 13832
rect 35806 11600 35862 11656
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34610 10512 34666 10568
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34518 3576 34574 3632
rect 36634 10240 36690 10296
rect 36818 9152 36874 9208
rect 36910 7792 36966 7848
rect 36266 6840 36322 6896
rect 36910 4020 36912 4040
rect 36912 4020 36964 4040
rect 36964 4020 36966 4040
rect 36910 3984 36966 4020
rect 36174 3848 36230 3904
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 37094 3712 37150 3768
rect 37738 9424 37794 9480
rect 37646 3712 37702 3768
rect 37922 8880 37978 8936
rect 38474 4800 38530 4856
rect 37738 3032 37794 3088
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 42890 25744 42946 25800
rect 43074 24520 43130 24576
rect 43350 30232 43406 30288
rect 43718 31048 43774 31104
rect 49514 39072 49570 39128
rect 44914 35128 44970 35184
rect 46110 35400 46166 35456
rect 43810 25336 43866 25392
rect 44454 24520 44510 24576
rect 42798 21256 42854 21312
rect 41878 13368 41934 13424
rect 45190 24384 45246 24440
rect 45466 24928 45522 24984
rect 45098 21936 45154 21992
rect 45006 21256 45062 21312
rect 44730 18264 44786 18320
rect 44638 17856 44694 17912
rect 45926 26288 45982 26344
rect 45742 24656 45798 24712
rect 45834 22344 45890 22400
rect 42706 6976 42762 7032
rect 43442 6840 43498 6896
rect 43718 3984 43774 4040
rect 43902 3848 43958 3904
rect 43902 3712 43958 3768
rect 45834 20168 45890 20224
rect 49514 33360 49570 33416
rect 47582 32272 47638 32328
rect 46110 31864 46166 31920
rect 46294 29552 46350 29608
rect 49514 29688 49570 29744
rect 46846 28736 46902 28792
rect 46386 28464 46442 28520
rect 46386 24656 46442 24712
rect 46754 27784 46810 27840
rect 47122 26832 47178 26888
rect 46662 25336 46718 25392
rect 47582 24384 47638 24440
rect 45650 8336 45706 8392
rect 46018 8472 46074 8528
rect 46294 6976 46350 7032
rect 45742 3576 45798 3632
rect 49514 20304 49570 20360
rect 49514 19352 49570 19408
rect 48226 14592 48282 14648
rect 47030 11464 47086 11520
rect 47214 7792 47270 7848
rect 46662 5208 46718 5264
rect 46478 1808 46534 1864
<< metal3 >>
rect 49520 48517 50000 48544
rect 49509 48514 50000 48517
rect 49428 48512 50000 48514
rect 49428 48456 49514 48512
rect 49570 48456 50000 48512
rect 49428 48454 50000 48456
rect 49509 48451 50000 48454
rect 49520 48424 50000 48451
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 22277 45386 22343 45389
rect 28441 45386 28507 45389
rect 36261 45386 36327 45389
rect 22277 45384 36327 45386
rect 22277 45328 22282 45384
rect 22338 45328 28446 45384
rect 28502 45328 36266 45384
rect 36322 45328 36327 45384
rect 22277 45326 36327 45328
rect 22277 45323 22343 45326
rect 28441 45323 28507 45326
rect 36261 45323 36327 45326
rect 49520 45296 50000 45416
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 44909 44842 44975 44845
rect 49558 44842 49618 45296
rect 44909 44840 49618 44842
rect 44909 44784 44914 44840
rect 44970 44784 49618 44840
rect 44909 44782 49618 44784
rect 44909 44779 44975 44782
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 37825 44298 37891 44301
rect 44817 44298 44883 44301
rect 37825 44296 44883 44298
rect 37825 44240 37830 44296
rect 37886 44240 44822 44296
rect 44878 44240 44883 44296
rect 37825 44238 44883 44240
rect 37825 44235 37891 44238
rect 44817 44235 44883 44238
rect 6085 44162 6151 44165
rect 19057 44162 19123 44165
rect 6085 44160 19123 44162
rect 6085 44104 6090 44160
rect 6146 44104 19062 44160
rect 19118 44104 19123 44160
rect 6085 44102 19123 44104
rect 6085 44099 6151 44102
rect 19057 44099 19123 44102
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 32949 43890 33015 43893
rect 41873 43890 41939 43893
rect 32949 43888 41939 43890
rect 32949 43832 32954 43888
rect 33010 43832 41878 43888
rect 41934 43832 41939 43888
rect 32949 43830 41939 43832
rect 32949 43827 33015 43830
rect 41873 43827 41939 43830
rect 19241 43754 19307 43757
rect 27061 43754 27127 43757
rect 19241 43752 27127 43754
rect 19241 43696 19246 43752
rect 19302 43696 27066 43752
rect 27122 43696 27127 43752
rect 19241 43694 27127 43696
rect 19241 43691 19307 43694
rect 27061 43691 27127 43694
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 19057 42938 19123 42941
rect 19425 42938 19491 42941
rect 19057 42936 19491 42938
rect 19057 42880 19062 42936
rect 19118 42880 19430 42936
rect 19486 42880 19491 42936
rect 19057 42878 19491 42880
rect 19057 42875 19123 42878
rect 19425 42875 19491 42878
rect 26785 42666 26851 42669
rect 34605 42666 34671 42669
rect 26785 42664 34671 42666
rect 26785 42608 26790 42664
rect 26846 42608 34610 42664
rect 34666 42608 34671 42664
rect 26785 42606 34671 42608
rect 26785 42603 26851 42606
rect 34605 42603 34671 42606
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 49520 42260 50000 42288
rect 49520 42258 49556 42260
rect 49428 42198 49556 42258
rect 49520 42196 49556 42198
rect 49620 42196 50000 42260
rect 49520 42168 50000 42196
rect 18597 42122 18663 42125
rect 26785 42122 26851 42125
rect 18597 42120 26851 42122
rect 18597 42064 18602 42120
rect 18658 42064 26790 42120
rect 26846 42064 26851 42120
rect 18597 42062 26851 42064
rect 18597 42059 18663 42062
rect 26785 42059 26851 42062
rect 34145 42122 34211 42125
rect 39757 42122 39823 42125
rect 34145 42120 39823 42122
rect 34145 42064 34150 42120
rect 34206 42064 39762 42120
rect 39818 42064 39823 42120
rect 34145 42062 39823 42064
rect 34145 42059 34211 42062
rect 39757 42059 39823 42062
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 0 41716 480 41744
rect 0 41652 60 41716
rect 124 41652 480 41716
rect 0 41624 480 41652
rect 14917 41578 14983 41581
rect 614 41576 14983 41578
rect 614 41520 14922 41576
rect 14978 41520 14983 41576
rect 614 41518 14983 41520
rect 54 41380 60 41444
rect 124 41442 130 41444
rect 614 41442 674 41518
rect 14917 41515 14983 41518
rect 124 41382 674 41442
rect 124 41380 130 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 32305 41034 32371 41037
rect 42517 41034 42583 41037
rect 43345 41034 43411 41037
rect 32305 41032 43411 41034
rect 32305 40976 32310 41032
rect 32366 40976 42522 41032
rect 42578 40976 43350 41032
rect 43406 40976 43411 41032
rect 32305 40974 43411 40976
rect 32305 40971 32371 40974
rect 42517 40971 42583 40974
rect 43345 40971 43411 40974
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 24485 40762 24551 40765
rect 24669 40762 24735 40765
rect 34145 40762 34211 40765
rect 24485 40760 34211 40762
rect 24485 40704 24490 40760
rect 24546 40704 24674 40760
rect 24730 40704 34150 40760
rect 34206 40704 34211 40760
rect 24485 40702 34211 40704
rect 24485 40699 24551 40702
rect 24669 40699 24735 40702
rect 34145 40699 34211 40702
rect 15929 40626 15995 40629
rect 24485 40626 24551 40629
rect 26509 40626 26575 40629
rect 15929 40624 26575 40626
rect 15929 40568 15934 40624
rect 15990 40568 24490 40624
rect 24546 40568 26514 40624
rect 26570 40568 26575 40624
rect 15929 40566 26575 40568
rect 15929 40563 15995 40566
rect 24485 40563 24551 40566
rect 26509 40563 26575 40566
rect 28809 40626 28875 40629
rect 32397 40626 32463 40629
rect 39481 40626 39547 40629
rect 28809 40624 39547 40626
rect 28809 40568 28814 40624
rect 28870 40568 32402 40624
rect 32458 40568 39486 40624
rect 39542 40568 39547 40624
rect 28809 40566 39547 40568
rect 28809 40563 28875 40566
rect 32397 40563 32463 40566
rect 39481 40563 39547 40566
rect 18965 40490 19031 40493
rect 29821 40490 29887 40493
rect 18965 40488 29887 40490
rect 18965 40432 18970 40488
rect 19026 40432 29826 40488
rect 29882 40432 29887 40488
rect 18965 40430 29887 40432
rect 18965 40427 19031 40430
rect 29821 40427 29887 40430
rect 26509 40354 26575 40357
rect 34237 40354 34303 40357
rect 26509 40352 34303 40354
rect 26509 40296 26514 40352
rect 26570 40296 34242 40352
rect 34298 40296 34303 40352
rect 26509 40294 34303 40296
rect 26509 40291 26575 40294
rect 34237 40291 34303 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 49520 39133 50000 39160
rect 49509 39130 50000 39133
rect 49428 39128 50000 39130
rect 49428 39072 49514 39128
rect 49570 39072 50000 39128
rect 49428 39070 50000 39072
rect 49509 39067 50000 39070
rect 49520 39040 50000 39067
rect 35801 38722 35867 38725
rect 43805 38722 43871 38725
rect 35801 38720 43871 38722
rect 35801 38664 35806 38720
rect 35862 38664 43810 38720
rect 43866 38664 43871 38720
rect 35801 38662 43871 38664
rect 35801 38659 35867 38662
rect 43805 38659 43871 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 27889 38314 27955 38317
rect 33409 38314 33475 38317
rect 27889 38312 33475 38314
rect 27889 38256 27894 38312
rect 27950 38256 33414 38312
rect 33470 38256 33475 38312
rect 27889 38254 33475 38256
rect 27889 38251 27955 38254
rect 33409 38251 33475 38254
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 49520 35912 50000 36032
rect 34928 35871 35248 35872
rect 26877 35730 26943 35733
rect 33777 35730 33843 35733
rect 26877 35728 33843 35730
rect 26877 35672 26882 35728
rect 26938 35672 33782 35728
rect 33838 35672 33843 35728
rect 26877 35670 33843 35672
rect 26877 35667 26943 35670
rect 33777 35667 33843 35670
rect 17493 35594 17559 35597
rect 28073 35594 28139 35597
rect 17493 35592 28139 35594
rect 17493 35536 17498 35592
rect 17554 35536 28078 35592
rect 28134 35536 28139 35592
rect 17493 35534 28139 35536
rect 17493 35531 17559 35534
rect 28073 35531 28139 35534
rect 46105 35458 46171 35461
rect 49558 35458 49618 35912
rect 46105 35456 49618 35458
rect 46105 35400 46110 35456
rect 46166 35400 49618 35456
rect 46105 35398 49618 35400
rect 46105 35395 46171 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 22645 35322 22711 35325
rect 28257 35322 28323 35325
rect 29729 35322 29795 35325
rect 22645 35320 29795 35322
rect 22645 35264 22650 35320
rect 22706 35264 28262 35320
rect 28318 35264 29734 35320
rect 29790 35264 29795 35320
rect 22645 35262 29795 35264
rect 22645 35259 22711 35262
rect 28257 35259 28323 35262
rect 29729 35259 29795 35262
rect 35617 35186 35683 35189
rect 44909 35186 44975 35189
rect 35617 35184 44975 35186
rect 35617 35128 35622 35184
rect 35678 35128 44914 35184
rect 44970 35128 44975 35184
rect 35617 35126 44975 35128
rect 35617 35123 35683 35126
rect 44909 35123 44975 35126
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 18597 34778 18663 34781
rect 23565 34778 23631 34781
rect 18597 34776 23631 34778
rect 18597 34720 18602 34776
rect 18658 34720 23570 34776
rect 23626 34720 23631 34776
rect 18597 34718 23631 34720
rect 18597 34715 18663 34718
rect 23565 34715 23631 34718
rect 36813 34642 36879 34645
rect 49550 34642 49556 34644
rect 36813 34640 49556 34642
rect 36813 34584 36818 34640
rect 36874 34584 49556 34640
rect 36813 34582 49556 34584
rect 36813 34579 36879 34582
rect 49550 34580 49556 34582
rect 49620 34580 49626 34644
rect 22829 34506 22895 34509
rect 28441 34506 28507 34509
rect 22829 34504 28507 34506
rect 22829 34448 22834 34504
rect 22890 34448 28446 34504
rect 28502 34448 28507 34504
rect 22829 34446 28507 34448
rect 22829 34443 22895 34446
rect 28441 34443 28507 34446
rect 33409 34506 33475 34509
rect 37825 34506 37891 34509
rect 33409 34504 37891 34506
rect 33409 34448 33414 34504
rect 33470 34448 37830 34504
rect 37886 34448 37891 34504
rect 33409 34446 37891 34448
rect 33409 34443 33475 34446
rect 37825 34443 37891 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 18505 34098 18571 34101
rect 25589 34098 25655 34101
rect 18505 34096 25655 34098
rect 18505 34040 18510 34096
rect 18566 34040 25594 34096
rect 25650 34040 25655 34096
rect 18505 34038 25655 34040
rect 18505 34035 18571 34038
rect 25589 34035 25655 34038
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 19057 33690 19123 33693
rect 26049 33690 26115 33693
rect 19057 33688 26115 33690
rect 19057 33632 19062 33688
rect 19118 33632 26054 33688
rect 26110 33632 26115 33688
rect 19057 33630 26115 33632
rect 19057 33627 19123 33630
rect 26049 33627 26115 33630
rect 34605 33418 34671 33421
rect 49509 33418 49575 33421
rect 34605 33416 49575 33418
rect 34605 33360 34610 33416
rect 34666 33360 49514 33416
rect 49570 33360 49575 33416
rect 34605 33358 49575 33360
rect 34605 33355 34671 33358
rect 49509 33355 49575 33358
rect 18965 33282 19031 33285
rect 19190 33282 19196 33284
rect 18965 33280 19196 33282
rect 18965 33224 18970 33280
rect 19026 33224 19196 33280
rect 18965 33222 19196 33224
rect 18965 33219 19031 33222
rect 19190 33220 19196 33222
rect 19260 33220 19266 33284
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 18965 33146 19031 33149
rect 35341 33146 35407 33149
rect 38193 33146 38259 33149
rect 18965 33144 19396 33146
rect 18965 33088 18970 33144
rect 19026 33088 19396 33144
rect 18965 33086 19396 33088
rect 18965 33083 19031 33086
rect 19336 33010 19396 33086
rect 35341 33144 38259 33146
rect 35341 33088 35346 33144
rect 35402 33088 38198 33144
rect 38254 33088 38259 33144
rect 35341 33086 38259 33088
rect 35341 33083 35407 33086
rect 38193 33083 38259 33086
rect 21357 33010 21423 33013
rect 19336 33008 21423 33010
rect 19336 32952 21362 33008
rect 21418 32952 21423 33008
rect 19336 32950 21423 32952
rect 21357 32947 21423 32950
rect 23749 33010 23815 33013
rect 32581 33010 32647 33013
rect 23749 33008 32647 33010
rect 23749 32952 23754 33008
rect 23810 32952 32586 33008
rect 32642 32952 32647 33008
rect 23749 32950 32647 32952
rect 23749 32947 23815 32950
rect 32581 32947 32647 32950
rect 17217 32874 17283 32877
rect 22737 32874 22803 32877
rect 17217 32872 22803 32874
rect 17217 32816 17222 32872
rect 17278 32816 22742 32872
rect 22798 32816 22803 32872
rect 17217 32814 22803 32816
rect 17217 32811 17283 32814
rect 22737 32811 22803 32814
rect 49520 32784 50000 32904
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 31845 32602 31911 32605
rect 34789 32602 34855 32605
rect 31845 32600 34855 32602
rect 31845 32544 31850 32600
rect 31906 32544 34794 32600
rect 34850 32544 34855 32600
rect 31845 32542 34855 32544
rect 31845 32539 31911 32542
rect 34789 32539 34855 32542
rect 47577 32330 47643 32333
rect 49558 32330 49618 32784
rect 47577 32328 49618 32330
rect 47577 32272 47582 32328
rect 47638 32272 49618 32328
rect 47577 32270 49618 32272
rect 47577 32267 47643 32270
rect 31477 32194 31543 32197
rect 36261 32194 36327 32197
rect 31477 32192 36327 32194
rect 31477 32136 31482 32192
rect 31538 32136 36266 32192
rect 36322 32136 36327 32192
rect 31477 32134 36327 32136
rect 31477 32131 31543 32134
rect 36261 32131 36327 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 15837 31922 15903 31925
rect 18229 31922 18295 31925
rect 15837 31920 18295 31922
rect 15837 31864 15842 31920
rect 15898 31864 18234 31920
rect 18290 31864 18295 31920
rect 15837 31862 18295 31864
rect 15837 31859 15903 31862
rect 18229 31859 18295 31862
rect 35065 31922 35131 31925
rect 46105 31922 46171 31925
rect 35065 31920 46171 31922
rect 35065 31864 35070 31920
rect 35126 31864 46110 31920
rect 46166 31864 46171 31920
rect 35065 31862 46171 31864
rect 35065 31859 35131 31862
rect 46105 31859 46171 31862
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19190 31452 19196 31516
rect 19260 31514 19266 31516
rect 19425 31514 19491 31517
rect 19260 31512 19491 31514
rect 19260 31456 19430 31512
rect 19486 31456 19491 31512
rect 19260 31454 19491 31456
rect 19260 31452 19266 31454
rect 19425 31451 19491 31454
rect 42057 31106 42123 31109
rect 43713 31106 43779 31109
rect 42057 31104 43779 31106
rect 42057 31048 42062 31104
rect 42118 31048 43718 31104
rect 43774 31048 43779 31104
rect 42057 31046 43779 31048
rect 42057 31043 42123 31046
rect 43713 31043 43779 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 28625 30970 28691 30973
rect 40309 30970 40375 30973
rect 28625 30968 40375 30970
rect 28625 30912 28630 30968
rect 28686 30912 40314 30968
rect 40370 30912 40375 30968
rect 28625 30910 40375 30912
rect 28625 30907 28691 30910
rect 40309 30907 40375 30910
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 22737 30290 22803 30293
rect 32213 30290 32279 30293
rect 22737 30288 32279 30290
rect 22737 30232 22742 30288
rect 22798 30232 32218 30288
rect 32274 30232 32279 30288
rect 22737 30230 32279 30232
rect 22737 30227 22803 30230
rect 32213 30227 32279 30230
rect 37549 30290 37615 30293
rect 43345 30290 43411 30293
rect 37549 30288 43411 30290
rect 37549 30232 37554 30288
rect 37610 30232 43350 30288
rect 43406 30232 43411 30288
rect 37549 30230 43411 30232
rect 37549 30227 37615 30230
rect 43345 30227 43411 30230
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 49520 29749 50000 29776
rect 12709 29746 12775 29749
rect 20621 29746 20687 29749
rect 49509 29746 50000 29749
rect 12709 29744 20687 29746
rect 12709 29688 12714 29744
rect 12770 29688 20626 29744
rect 20682 29688 20687 29744
rect 12709 29686 20687 29688
rect 49428 29744 50000 29746
rect 49428 29688 49514 29744
rect 49570 29688 50000 29744
rect 49428 29686 50000 29688
rect 12709 29683 12775 29686
rect 20621 29683 20687 29686
rect 49509 29683 50000 29686
rect 49520 29656 50000 29683
rect 37457 29610 37523 29613
rect 46289 29610 46355 29613
rect 37457 29608 46355 29610
rect 37457 29552 37462 29608
rect 37518 29552 46294 29608
rect 46350 29552 46355 29608
rect 37457 29550 46355 29552
rect 37457 29547 37523 29550
rect 46289 29547 46355 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 31845 29066 31911 29069
rect 36353 29066 36419 29069
rect 31845 29064 36419 29066
rect 31845 29008 31850 29064
rect 31906 29008 36358 29064
rect 36414 29008 36419 29064
rect 31845 29006 36419 29008
rect 31845 29003 31911 29006
rect 36353 29003 36419 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 20897 28794 20963 28797
rect 29729 28794 29795 28797
rect 20897 28792 29795 28794
rect 20897 28736 20902 28792
rect 20958 28736 29734 28792
rect 29790 28736 29795 28792
rect 20897 28734 29795 28736
rect 20897 28731 20963 28734
rect 29729 28731 29795 28734
rect 37089 28794 37155 28797
rect 46841 28794 46907 28797
rect 37089 28792 46907 28794
rect 37089 28736 37094 28792
rect 37150 28736 46846 28792
rect 46902 28736 46907 28792
rect 37089 28734 46907 28736
rect 37089 28731 37155 28734
rect 46841 28731 46907 28734
rect 14365 28658 14431 28661
rect 32857 28658 32923 28661
rect 34237 28658 34303 28661
rect 14365 28656 34303 28658
rect 14365 28600 14370 28656
rect 14426 28600 32862 28656
rect 32918 28600 34242 28656
rect 34298 28600 34303 28656
rect 14365 28598 34303 28600
rect 14365 28595 14431 28598
rect 32857 28595 32923 28598
rect 34237 28595 34303 28598
rect 19241 28522 19307 28525
rect 23473 28522 23539 28525
rect 19241 28520 23539 28522
rect 19241 28464 19246 28520
rect 19302 28464 23478 28520
rect 23534 28464 23539 28520
rect 19241 28462 23539 28464
rect 19241 28459 19307 28462
rect 23473 28459 23539 28462
rect 36077 28522 36143 28525
rect 46381 28522 46447 28525
rect 36077 28520 46447 28522
rect 36077 28464 36082 28520
rect 36138 28464 46386 28520
rect 46442 28464 46447 28520
rect 36077 28462 46447 28464
rect 36077 28459 36143 28462
rect 46381 28459 46447 28462
rect 19374 28324 19380 28388
rect 19444 28386 19450 28388
rect 19885 28386 19951 28389
rect 19444 28384 19951 28386
rect 19444 28328 19890 28384
rect 19946 28328 19951 28384
rect 19444 28326 19951 28328
rect 19444 28324 19450 28326
rect 19885 28323 19951 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 24117 27842 24183 27845
rect 30281 27842 30347 27845
rect 46749 27842 46815 27845
rect 24117 27840 46815 27842
rect 24117 27784 24122 27840
rect 24178 27784 30286 27840
rect 30342 27784 46754 27840
rect 46810 27784 46815 27840
rect 24117 27782 46815 27784
rect 24117 27779 24183 27782
rect 30281 27779 30347 27782
rect 46749 27779 46815 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 16113 27026 16179 27029
rect 26417 27026 26483 27029
rect 16113 27024 26483 27026
rect 16113 26968 16118 27024
rect 16174 26968 26422 27024
rect 26478 26968 26483 27024
rect 16113 26966 26483 26968
rect 16113 26963 16179 26966
rect 26417 26963 26483 26966
rect 17217 26890 17283 26893
rect 24853 26890 24919 26893
rect 17217 26888 24919 26890
rect 17217 26832 17222 26888
rect 17278 26832 24858 26888
rect 24914 26832 24919 26888
rect 17217 26830 24919 26832
rect 17217 26827 17283 26830
rect 24853 26827 24919 26830
rect 33593 26890 33659 26893
rect 38469 26890 38535 26893
rect 47117 26890 47183 26893
rect 33593 26888 47183 26890
rect 33593 26832 33598 26888
rect 33654 26832 38474 26888
rect 38530 26832 47122 26888
rect 47178 26832 47183 26888
rect 33593 26830 47183 26832
rect 33593 26827 33659 26830
rect 38469 26827 38535 26830
rect 47117 26827 47183 26830
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 49520 26528 50000 26648
rect 45921 26346 45987 26349
rect 49558 26346 49618 26528
rect 45921 26344 49618 26346
rect 45921 26288 45926 26344
rect 45982 26288 49618 26344
rect 45921 26286 49618 26288
rect 45921 26283 45987 26286
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 14365 26074 14431 26077
rect 25037 26074 25103 26077
rect 14365 26072 25103 26074
rect 14365 26016 14370 26072
rect 14426 26016 25042 26072
rect 25098 26016 25103 26072
rect 14365 26014 25103 26016
rect 14365 26011 14431 26014
rect 25037 26011 25103 26014
rect 15745 25938 15811 25941
rect 23933 25938 23999 25941
rect 28717 25938 28783 25941
rect 33593 25938 33659 25941
rect 15745 25936 23999 25938
rect 15745 25880 15750 25936
rect 15806 25880 23938 25936
rect 23994 25880 23999 25936
rect 15745 25878 23999 25880
rect 15745 25875 15811 25878
rect 23933 25875 23999 25878
rect 27294 25936 33659 25938
rect 27294 25880 28722 25936
rect 28778 25880 33598 25936
rect 33654 25880 33659 25936
rect 27294 25878 33659 25880
rect 13537 25802 13603 25805
rect 22829 25802 22895 25805
rect 24945 25802 25011 25805
rect 27294 25802 27354 25878
rect 28717 25875 28783 25878
rect 33593 25875 33659 25878
rect 13537 25800 13830 25802
rect 13537 25744 13542 25800
rect 13598 25744 13830 25800
rect 13537 25742 13830 25744
rect 13537 25739 13603 25742
rect 13770 25258 13830 25742
rect 22829 25800 27354 25802
rect 22829 25744 22834 25800
rect 22890 25744 24950 25800
rect 25006 25744 27354 25800
rect 22829 25742 27354 25744
rect 34789 25802 34855 25805
rect 42885 25802 42951 25805
rect 34789 25800 42951 25802
rect 34789 25744 34794 25800
rect 34850 25744 42890 25800
rect 42946 25744 42951 25800
rect 34789 25742 42951 25744
rect 22829 25739 22895 25742
rect 24945 25739 25011 25742
rect 34789 25739 34855 25742
rect 42885 25739 42951 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 27889 25530 27955 25533
rect 33869 25530 33935 25533
rect 27889 25528 33935 25530
rect 27889 25472 27894 25528
rect 27950 25472 33874 25528
rect 33930 25472 33935 25528
rect 27889 25470 33935 25472
rect 27889 25467 27955 25470
rect 33869 25467 33935 25470
rect 33685 25394 33751 25397
rect 37825 25394 37891 25397
rect 43805 25394 43871 25397
rect 46657 25394 46723 25397
rect 33685 25392 46723 25394
rect 33685 25336 33690 25392
rect 33746 25336 37830 25392
rect 37886 25336 43810 25392
rect 43866 25336 46662 25392
rect 46718 25336 46723 25392
rect 33685 25334 46723 25336
rect 33685 25331 33751 25334
rect 37825 25331 37891 25334
rect 43805 25331 43871 25334
rect 46657 25331 46723 25334
rect 62 25198 13830 25258
rect 62 25016 122 25198
rect 13770 25122 13830 25198
rect 14181 25258 14247 25261
rect 30833 25258 30899 25261
rect 14181 25256 30899 25258
rect 14181 25200 14186 25256
rect 14242 25200 30838 25256
rect 30894 25200 30899 25256
rect 14181 25198 30899 25200
rect 14181 25195 14247 25198
rect 30833 25195 30899 25198
rect 14273 25122 14339 25125
rect 13770 25120 14339 25122
rect 13770 25064 14278 25120
rect 14334 25064 14339 25120
rect 13770 25062 14339 25064
rect 14273 25059 14339 25062
rect 4208 25056 4528 25057
rect 0 24896 480 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 36169 24986 36235 24989
rect 45461 24986 45527 24989
rect 36169 24984 45527 24986
rect 36169 24928 36174 24984
rect 36230 24928 45466 24984
rect 45522 24928 45527 24984
rect 36169 24926 45527 24928
rect 36169 24923 36235 24926
rect 45461 24923 45527 24926
rect 37273 24714 37339 24717
rect 45737 24714 45803 24717
rect 46381 24714 46447 24717
rect 37273 24712 46447 24714
rect 37273 24656 37278 24712
rect 37334 24656 45742 24712
rect 45798 24656 46386 24712
rect 46442 24656 46447 24712
rect 37273 24654 46447 24656
rect 37273 24651 37339 24654
rect 45737 24651 45803 24654
rect 46381 24651 46447 24654
rect 34237 24578 34303 24581
rect 43069 24578 43135 24581
rect 44449 24578 44515 24581
rect 34237 24576 44515 24578
rect 34237 24520 34242 24576
rect 34298 24520 43074 24576
rect 43130 24520 44454 24576
rect 44510 24520 44515 24576
rect 34237 24518 44515 24520
rect 34237 24515 34303 24518
rect 43069 24515 43135 24518
rect 44449 24515 44515 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 30189 24442 30255 24445
rect 35341 24442 35407 24445
rect 45185 24442 45251 24445
rect 47577 24442 47643 24445
rect 30189 24440 47643 24442
rect 30189 24384 30194 24440
rect 30250 24384 35346 24440
rect 35402 24384 45190 24440
rect 45246 24384 47582 24440
rect 47638 24384 47643 24440
rect 30189 24382 47643 24384
rect 30189 24379 30255 24382
rect 35341 24379 35407 24382
rect 45185 24379 45251 24382
rect 47577 24379 47643 24382
rect 19057 24306 19123 24309
rect 26325 24306 26391 24309
rect 19057 24304 26391 24306
rect 19057 24248 19062 24304
rect 19118 24248 26330 24304
rect 26386 24248 26391 24304
rect 19057 24246 26391 24248
rect 19057 24243 19123 24246
rect 26325 24243 26391 24246
rect 14641 24034 14707 24037
rect 23657 24034 23723 24037
rect 14641 24032 23723 24034
rect 14641 23976 14646 24032
rect 14702 23976 23662 24032
rect 23718 23976 23723 24032
rect 14641 23974 23723 23976
rect 14641 23971 14707 23974
rect 23657 23971 23723 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 17585 23898 17651 23901
rect 27337 23898 27403 23901
rect 17585 23896 27403 23898
rect 17585 23840 17590 23896
rect 17646 23840 27342 23896
rect 27398 23840 27403 23896
rect 17585 23838 27403 23840
rect 17585 23835 17651 23838
rect 27337 23835 27403 23838
rect 14089 23762 14155 23765
rect 20437 23762 20503 23765
rect 14089 23760 23490 23762
rect 14089 23704 14094 23760
rect 14150 23704 20442 23760
rect 20498 23704 23490 23760
rect 14089 23702 23490 23704
rect 14089 23699 14155 23702
rect 20437 23699 20503 23702
rect 14273 23626 14339 23629
rect 21265 23626 21331 23629
rect 14273 23624 21331 23626
rect 14273 23568 14278 23624
rect 14334 23568 21270 23624
rect 21326 23568 21331 23624
rect 14273 23566 21331 23568
rect 14273 23563 14339 23566
rect 21265 23563 21331 23566
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 23430 23354 23490 23702
rect 32581 23626 32647 23629
rect 32857 23626 32923 23629
rect 38653 23626 38719 23629
rect 32581 23624 38719 23626
rect 32581 23568 32586 23624
rect 32642 23568 32862 23624
rect 32918 23568 38658 23624
rect 38714 23568 38719 23624
rect 32581 23566 38719 23568
rect 32581 23563 32647 23566
rect 32857 23563 32923 23566
rect 38653 23563 38719 23566
rect 49520 23462 50000 23520
rect 49520 23460 49556 23462
rect 49428 23400 49556 23460
rect 49550 23398 49556 23400
rect 49620 23400 50000 23462
rect 49620 23398 49626 23400
rect 27429 23354 27495 23357
rect 32029 23354 32095 23357
rect 23430 23352 32095 23354
rect 23430 23296 27434 23352
rect 27490 23296 32034 23352
rect 32090 23296 32095 23352
rect 23430 23294 32095 23296
rect 27429 23291 27495 23294
rect 32029 23291 32095 23294
rect 27337 23218 27403 23221
rect 31201 23218 31267 23221
rect 27337 23216 31267 23218
rect 27337 23160 27342 23216
rect 27398 23160 31206 23216
rect 31262 23160 31267 23216
rect 27337 23158 31267 23160
rect 27337 23155 27403 23158
rect 31201 23155 31267 23158
rect 28533 22946 28599 22949
rect 23430 22944 28599 22946
rect 23430 22888 28538 22944
rect 28594 22888 28599 22944
rect 23430 22886 28599 22888
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 21541 22810 21607 22813
rect 23430 22810 23490 22886
rect 28533 22883 28599 22886
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 21541 22808 23490 22810
rect 21541 22752 21546 22808
rect 21602 22752 23490 22808
rect 21541 22750 23490 22752
rect 24853 22810 24919 22813
rect 31017 22810 31083 22813
rect 24853 22808 31083 22810
rect 24853 22752 24858 22808
rect 24914 22752 31022 22808
rect 31078 22752 31083 22808
rect 24853 22750 31083 22752
rect 21541 22747 21607 22750
rect 24853 22747 24919 22750
rect 31017 22747 31083 22750
rect 17217 22674 17283 22677
rect 25037 22674 25103 22677
rect 17217 22672 25103 22674
rect 17217 22616 17222 22672
rect 17278 22616 25042 22672
rect 25098 22616 25103 22672
rect 17217 22614 25103 22616
rect 17217 22611 17283 22614
rect 25037 22611 25103 22614
rect 31385 22402 31451 22405
rect 45829 22402 45895 22405
rect 31385 22400 45895 22402
rect 31385 22344 31390 22400
rect 31446 22344 45834 22400
rect 45890 22344 45895 22400
rect 31385 22342 45895 22344
rect 31385 22339 31451 22342
rect 45829 22339 45895 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 28533 21994 28599 21997
rect 32254 21994 32260 21996
rect 28533 21992 32260 21994
rect 28533 21936 28538 21992
rect 28594 21936 32260 21992
rect 28533 21934 32260 21936
rect 28533 21931 28599 21934
rect 32254 21932 32260 21934
rect 32324 21994 32330 21996
rect 35985 21994 36051 21997
rect 45093 21994 45159 21997
rect 32324 21992 45159 21994
rect 32324 21936 35990 21992
rect 36046 21936 45098 21992
rect 45154 21936 45159 21992
rect 32324 21934 45159 21936
rect 32324 21932 32330 21934
rect 35985 21931 36051 21934
rect 45093 21931 45159 21934
rect 23657 21858 23723 21861
rect 30741 21858 30807 21861
rect 23657 21856 30807 21858
rect 23657 21800 23662 21856
rect 23718 21800 30746 21856
rect 30802 21800 30807 21856
rect 23657 21798 30807 21800
rect 23657 21795 23723 21798
rect 30741 21795 30807 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 19241 21722 19307 21725
rect 19374 21722 19380 21724
rect 19241 21720 19380 21722
rect 19241 21664 19246 21720
rect 19302 21664 19380 21720
rect 19241 21662 19380 21664
rect 19241 21659 19307 21662
rect 19374 21660 19380 21662
rect 19444 21660 19450 21724
rect 16481 21450 16547 21453
rect 20805 21450 20871 21453
rect 24117 21450 24183 21453
rect 16481 21448 24183 21450
rect 16481 21392 16486 21448
rect 16542 21392 20810 21448
rect 20866 21392 24122 21448
rect 24178 21392 24183 21448
rect 16481 21390 24183 21392
rect 16481 21387 16547 21390
rect 20805 21387 20871 21390
rect 24117 21387 24183 21390
rect 37733 21314 37799 21317
rect 42793 21314 42859 21317
rect 45001 21314 45067 21317
rect 37733 21312 45067 21314
rect 37733 21256 37738 21312
rect 37794 21256 42798 21312
rect 42854 21256 45006 21312
rect 45062 21256 45067 21312
rect 37733 21254 45067 21256
rect 37733 21251 37799 21254
rect 42793 21251 42859 21254
rect 45001 21251 45067 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 49520 20365 50000 20392
rect 49509 20362 50000 20365
rect 49428 20360 50000 20362
rect 49428 20304 49514 20360
rect 49570 20304 50000 20360
rect 49428 20302 50000 20304
rect 49509 20299 50000 20302
rect 49520 20272 50000 20299
rect 32305 20226 32371 20229
rect 45829 20226 45895 20229
rect 32305 20224 45895 20226
rect 32305 20168 32310 20224
rect 32366 20168 45834 20224
rect 45890 20168 45895 20224
rect 32305 20166 45895 20168
rect 32305 20163 32371 20166
rect 45829 20163 45895 20166
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 27981 19410 28047 19413
rect 36169 19410 36235 19413
rect 27981 19408 36235 19410
rect 27981 19352 27986 19408
rect 28042 19352 36174 19408
rect 36230 19352 36235 19408
rect 27981 19350 36235 19352
rect 27981 19347 28047 19350
rect 36169 19347 36235 19350
rect 36353 19410 36419 19413
rect 49509 19410 49575 19413
rect 36353 19408 49575 19410
rect 36353 19352 36358 19408
rect 36414 19352 49514 19408
rect 49570 19352 49575 19408
rect 36353 19350 49575 19352
rect 36353 19347 36419 19350
rect 49509 19347 49575 19350
rect 23105 19274 23171 19277
rect 23749 19274 23815 19277
rect 23105 19272 23815 19274
rect 23105 19216 23110 19272
rect 23166 19216 23754 19272
rect 23810 19216 23815 19272
rect 23105 19214 23815 19216
rect 23105 19211 23171 19214
rect 23749 19211 23815 19214
rect 23933 19272 23999 19277
rect 23933 19216 23938 19272
rect 23994 19216 23999 19272
rect 23933 19211 23999 19216
rect 23381 19138 23447 19141
rect 23936 19138 23996 19211
rect 23381 19136 23996 19138
rect 23381 19080 23386 19136
rect 23442 19080 23996 19136
rect 23381 19078 23996 19080
rect 31293 19138 31359 19141
rect 32765 19138 32831 19141
rect 31293 19136 32831 19138
rect 31293 19080 31298 19136
rect 31354 19080 32770 19136
rect 32826 19080 32831 19136
rect 31293 19078 32831 19080
rect 23381 19075 23447 19078
rect 31293 19075 31359 19078
rect 32765 19075 32831 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 32949 18866 33015 18869
rect 34513 18866 34579 18869
rect 49550 18866 49556 18868
rect 32949 18864 49556 18866
rect 32949 18808 32954 18864
rect 33010 18808 34518 18864
rect 34574 18808 49556 18864
rect 32949 18806 49556 18808
rect 32949 18803 33015 18806
rect 34513 18803 34579 18806
rect 49550 18804 49556 18806
rect 49620 18804 49626 18868
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 35801 18322 35867 18325
rect 44725 18322 44791 18325
rect 35801 18320 44791 18322
rect 35801 18264 35806 18320
rect 35862 18264 44730 18320
rect 44786 18264 44791 18320
rect 35801 18262 44791 18264
rect 35801 18259 35867 18262
rect 44725 18259 44791 18262
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 37365 17914 37431 17917
rect 44633 17914 44699 17917
rect 37365 17912 44699 17914
rect 37365 17856 37370 17912
rect 37426 17856 44638 17912
rect 44694 17856 44699 17912
rect 37365 17854 44699 17856
rect 37365 17851 37431 17854
rect 44633 17851 44699 17854
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 49520 17144 50000 17264
rect 35801 16962 35867 16965
rect 49558 16962 49618 17144
rect 35801 16960 49618 16962
rect 35801 16904 35806 16960
rect 35862 16904 49618 16960
rect 35801 16902 49618 16904
rect 35801 16899 35867 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 18137 16554 18203 16557
rect 20069 16554 20135 16557
rect 31201 16554 31267 16557
rect 18137 16552 31267 16554
rect 18137 16496 18142 16552
rect 18198 16496 20074 16552
rect 20130 16496 31206 16552
rect 31262 16496 31267 16552
rect 18137 16494 31267 16496
rect 18137 16491 18203 16494
rect 20069 16491 20135 16494
rect 31201 16491 31267 16494
rect 23105 16418 23171 16421
rect 30925 16418 30991 16421
rect 23105 16416 30991 16418
rect 23105 16360 23110 16416
rect 23166 16360 30930 16416
rect 30986 16360 30991 16416
rect 23105 16358 30991 16360
rect 23105 16355 23171 16358
rect 30925 16355 30991 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 32029 15058 32095 15061
rect 32254 15058 32260 15060
rect 32029 15056 32260 15058
rect 32029 15000 32034 15056
rect 32090 15000 32260 15056
rect 32029 14998 32260 15000
rect 32029 14995 32095 14998
rect 32254 14996 32260 14998
rect 32324 14996 32330 15060
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 48221 14650 48287 14653
rect 48221 14648 49618 14650
rect 48221 14592 48226 14648
rect 48282 14592 49618 14648
rect 48221 14590 49618 14592
rect 48221 14587 48287 14590
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 49558 14136 49618 14590
rect 34928 14111 35248 14112
rect 49520 14016 50000 14136
rect 17953 13834 18019 13837
rect 19241 13834 19307 13837
rect 17953 13832 19307 13834
rect 17953 13776 17958 13832
rect 18014 13776 19246 13832
rect 19302 13776 19307 13832
rect 17953 13774 19307 13776
rect 17953 13771 18019 13774
rect 19241 13771 19307 13774
rect 33869 13834 33935 13837
rect 36353 13834 36419 13837
rect 33869 13832 36419 13834
rect 33869 13776 33874 13832
rect 33930 13776 36358 13832
rect 36414 13776 36419 13832
rect 33869 13774 36419 13776
rect 33869 13771 33935 13774
rect 36353 13771 36419 13774
rect 19057 13698 19123 13701
rect 19287 13698 19353 13701
rect 19057 13696 19353 13698
rect 19057 13640 19062 13696
rect 19118 13640 19292 13696
rect 19348 13640 19353 13696
rect 19057 13638 19353 13640
rect 19057 13635 19123 13638
rect 19287 13635 19353 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 19425 13426 19491 13429
rect 41873 13426 41939 13429
rect 19425 13424 41939 13426
rect 19425 13368 19430 13424
rect 19486 13368 41878 13424
rect 41934 13368 41939 13424
rect 19425 13366 41939 13368
rect 19425 13363 19491 13366
rect 41873 13363 41939 13366
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 26325 12746 26391 12749
rect 33869 12746 33935 12749
rect 26325 12744 33935 12746
rect 26325 12688 26330 12744
rect 26386 12688 33874 12744
rect 33930 12688 33935 12744
rect 26325 12686 33935 12688
rect 26325 12683 26391 12686
rect 33869 12683 33935 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 27889 11658 27955 11661
rect 35801 11658 35867 11661
rect 27889 11656 35867 11658
rect 27889 11600 27894 11656
rect 27950 11600 35806 11656
rect 35862 11600 35867 11656
rect 27889 11598 35867 11600
rect 27889 11595 27955 11598
rect 35801 11595 35867 11598
rect 47025 11522 47091 11525
rect 47025 11520 49618 11522
rect 47025 11464 47030 11520
rect 47086 11464 49618 11520
rect 47025 11462 49618 11464
rect 47025 11459 47091 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 49558 11008 49618 11462
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 49520 10888 50000 11008
rect 34928 10847 35248 10848
rect 28625 10570 28691 10573
rect 34605 10570 34671 10573
rect 28625 10568 34671 10570
rect 28625 10512 28630 10568
rect 28686 10512 34610 10568
rect 34666 10512 34671 10568
rect 28625 10510 34671 10512
rect 28625 10507 28691 10510
rect 34605 10507 34671 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 21817 10298 21883 10301
rect 36629 10298 36695 10301
rect 21817 10296 36695 10298
rect 21817 10240 21822 10296
rect 21878 10240 36634 10296
rect 36690 10240 36695 10296
rect 21817 10238 36695 10240
rect 21817 10235 21883 10238
rect 36629 10235 36695 10238
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 24853 9482 24919 9485
rect 37733 9482 37799 9485
rect 24853 9480 37799 9482
rect 24853 9424 24858 9480
rect 24914 9424 37738 9480
rect 37794 9424 37799 9480
rect 24853 9422 37799 9424
rect 24853 9419 24919 9422
rect 37733 9419 37799 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 23749 9210 23815 9213
rect 36813 9210 36879 9213
rect 23749 9208 36879 9210
rect 23749 9152 23754 9208
rect 23810 9152 36818 9208
rect 36874 9152 36879 9208
rect 23749 9150 36879 9152
rect 23749 9147 23815 9150
rect 36813 9147 36879 9150
rect 13813 8938 13879 8941
rect 62 8936 13879 8938
rect 62 8880 13818 8936
rect 13874 8880 13879 8936
rect 62 8878 13879 8880
rect 62 8424 122 8878
rect 13813 8875 13879 8878
rect 21449 8938 21515 8941
rect 37917 8938 37983 8941
rect 21449 8936 37983 8938
rect 21449 8880 21454 8936
rect 21510 8880 37922 8936
rect 37978 8880 37983 8936
rect 21449 8878 37983 8880
rect 21449 8875 21515 8878
rect 37917 8875 37983 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 19977 8530 20043 8533
rect 46013 8530 46079 8533
rect 19977 8528 46079 8530
rect 19977 8472 19982 8528
rect 20038 8472 46018 8528
rect 46074 8472 46079 8528
rect 19977 8470 46079 8472
rect 19977 8467 20043 8470
rect 46013 8467 46079 8470
rect 0 8304 480 8424
rect 45645 8394 45711 8397
rect 45645 8392 49618 8394
rect 45645 8336 45650 8392
rect 45706 8336 49618 8392
rect 45645 8334 49618 8336
rect 45645 8331 45711 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 49558 7880 49618 8334
rect 36905 7850 36971 7853
rect 47209 7850 47275 7853
rect 36905 7848 47275 7850
rect 36905 7792 36910 7848
rect 36966 7792 47214 7848
rect 47270 7792 47275 7848
rect 36905 7790 47275 7792
rect 36905 7787 36971 7790
rect 47209 7787 47275 7790
rect 49520 7760 50000 7880
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 42701 7034 42767 7037
rect 46289 7034 46355 7037
rect 42701 7032 46355 7034
rect 42701 6976 42706 7032
rect 42762 6976 46294 7032
rect 46350 6976 46355 7032
rect 42701 6974 46355 6976
rect 42701 6971 42767 6974
rect 46289 6971 46355 6974
rect 36261 6898 36327 6901
rect 43437 6898 43503 6901
rect 36261 6896 43503 6898
rect 36261 6840 36266 6896
rect 36322 6840 43442 6896
rect 43498 6840 43503 6896
rect 36261 6838 43503 6840
rect 36261 6835 36327 6838
rect 43437 6835 43503 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 20529 5674 20595 5677
rect 27245 5674 27311 5677
rect 20529 5672 27311 5674
rect 20529 5616 20534 5672
rect 20590 5616 27250 5672
rect 27306 5616 27311 5672
rect 20529 5614 27311 5616
rect 20529 5611 20595 5614
rect 27245 5611 27311 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 46657 5266 46723 5269
rect 46657 5264 49618 5266
rect 46657 5208 46662 5264
rect 46718 5208 49618 5264
rect 46657 5206 49618 5208
rect 46657 5203 46723 5206
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 22277 4858 22343 4861
rect 38469 4858 38535 4861
rect 22277 4856 38535 4858
rect 22277 4800 22282 4856
rect 22338 4800 38474 4856
rect 38530 4800 38535 4856
rect 22277 4798 38535 4800
rect 22277 4795 22343 4798
rect 38469 4795 38535 4798
rect 49558 4752 49618 5206
rect 49520 4632 50000 4752
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 36905 4042 36971 4045
rect 43713 4042 43779 4045
rect 36905 4040 43779 4042
rect 36905 3984 36910 4040
rect 36966 3984 43718 4040
rect 43774 3984 43779 4040
rect 36905 3982 43779 3984
rect 36905 3979 36971 3982
rect 43713 3979 43779 3982
rect 36169 3906 36235 3909
rect 43897 3906 43963 3909
rect 36169 3904 43963 3906
rect 36169 3848 36174 3904
rect 36230 3848 43902 3904
rect 43958 3848 43963 3904
rect 36169 3846 43963 3848
rect 36169 3843 36235 3846
rect 43897 3843 43963 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 24393 3770 24459 3773
rect 37089 3770 37155 3773
rect 24393 3768 37155 3770
rect 24393 3712 24398 3768
rect 24454 3712 37094 3768
rect 37150 3712 37155 3768
rect 24393 3710 37155 3712
rect 24393 3707 24459 3710
rect 37089 3707 37155 3710
rect 37641 3770 37707 3773
rect 43897 3770 43963 3773
rect 37641 3768 43963 3770
rect 37641 3712 37646 3768
rect 37702 3712 43902 3768
rect 43958 3712 43963 3768
rect 37641 3710 43963 3712
rect 37641 3707 37707 3710
rect 43897 3707 43963 3710
rect 34513 3634 34579 3637
rect 45737 3634 45803 3637
rect 34513 3632 45803 3634
rect 34513 3576 34518 3632
rect 34574 3576 45742 3632
rect 45798 3576 45803 3632
rect 34513 3574 45803 3576
rect 34513 3571 34579 3574
rect 45737 3571 45803 3574
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 22093 3090 22159 3093
rect 37733 3090 37799 3093
rect 22093 3088 37799 3090
rect 22093 3032 22098 3088
rect 22154 3032 37738 3088
rect 37794 3032 37799 3088
rect 22093 3030 37799 3032
rect 22093 3027 22159 3030
rect 37733 3027 37799 3030
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 3785 2002 3851 2005
rect 17125 2002 17191 2005
rect 3785 2000 17191 2002
rect 3785 1944 3790 2000
rect 3846 1944 17130 2000
rect 17186 1944 17191 2000
rect 3785 1942 17191 1944
rect 3785 1939 3851 1942
rect 17125 1939 17191 1942
rect 46473 1866 46539 1869
rect 46473 1864 49618 1866
rect 46473 1808 46478 1864
rect 46534 1808 49618 1864
rect 46473 1806 49618 1808
rect 46473 1803 46539 1806
rect 49558 1624 49618 1806
rect 49520 1504 50000 1624
<< via3 >>
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 49556 42196 49620 42260
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 60 41652 124 41716
rect 60 41380 124 41444
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 49556 34580 49620 34644
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19196 33220 19260 33284
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19196 31452 19260 31516
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 19380 28324 19444 28388
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 49556 23398 49620 23462
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 32260 21932 32324 21996
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19380 21660 19444 21724
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 49556 18804 49620 18868
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 32260 14996 32324 15060
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 46816 4528 47376
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 59 41716 125 41717
rect 59 41652 60 41716
rect 124 41652 125 41716
rect 59 41651 125 41652
rect 62 41445 122 41651
rect 59 41444 125 41445
rect 59 41380 60 41444
rect 124 41380 125 41444
rect 59 41379 125 41380
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 19568 47360 19888 47376
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19195 33284 19261 33285
rect 19195 33220 19196 33284
rect 19260 33220 19261 33284
rect 19195 33219 19261 33220
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 19198 31517 19258 33219
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19195 31516 19261 31517
rect 19195 31452 19196 31516
rect 19260 31452 19261 31516
rect 19195 31451 19261 31452
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19379 28388 19445 28389
rect 19379 28324 19380 28388
rect 19444 28324 19445 28388
rect 19379 28323 19445 28324
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 19382 21725 19442 28323
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19379 21724 19445 21725
rect 19379 21660 19380 21724
rect 19444 21660 19445 21724
rect 19379 21659 19445 21660
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 21248 19888 22272
rect 34928 46816 35248 47376
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 49555 42260 49621 42261
rect 49555 42196 49556 42260
rect 49620 42196 49621 42260
rect 49555 42195 49621 42196
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 49558 34645 49618 42195
rect 49555 34644 49621 34645
rect 49555 34580 49556 34644
rect 49620 34580 49621 34644
rect 49555 34579 49621 34580
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 49555 23462 49621 23463
rect 49555 23398 49556 23462
rect 49620 23398 49621 23462
rect 49555 23397 49621 23398
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 32259 21996 32325 21997
rect 32259 21932 32260 21996
rect 32324 21932 32325 21996
rect 32259 21931 32325 21932
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 32262 15061 32322 21931
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 49558 18869 49618 23397
rect 49555 18868 49621 18869
rect 49555 18804 49556 18868
rect 49620 18804 49621 18868
rect 49555 18803 49621 18804
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 32259 15060 32325 15061
rect 32259 14996 32260 15060
rect 32324 14996 32325 15060
rect 32259 14995 32325 14996
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__594__B
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__594__A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_222 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _594_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_234
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_246
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__591__A
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__591__B
timestamp 1586364061
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_278
timestamp 1586364061
transform 1 0 26680 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_282
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_289
timestamp 1586364061
transform 1 0 27692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_283
timestamp 1586364061
transform 1 0 27140 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__586__B
timestamp 1586364061
transform 1 0 27508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__586__A
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _586_
timestamp 1586364061
transform 1 0 28060 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__587__B
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_314
timestamp 1586364061
transform 1 0 29992 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_309
timestamp 1586364061
transform 1 0 29532 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__584__B
timestamp 1586364061
transform 1 0 29808 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__587__A
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__584__A
timestamp 1586364061
transform 1 0 30176 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_nor2_4  _587_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_324
timestamp 1586364061
transform 1 0 30912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31096 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_333
timestamp 1586364061
transform 1 0 31740 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__251__B
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_345
timestamp 1586364061
transform 1 0 32844 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_345
timestamp 1586364061
transform 1 0 32844 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__262__B
timestamp 1586364061
transform 1 0 32660 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 33028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_358
timestamp 1586364061
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_351
timestamp 1586364061
transform 1 0 33396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 33212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _262_
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _251_
timestamp 1586364061
transform 1 0 33580 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_362
timestamp 1586364061
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__251__A
timestamp 1586364061
transform 1 0 34592 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_1_382
timestamp 1586364061
transform 1 0 36248 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_378
timestamp 1586364061
transform 1 0 35880 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_384
timestamp 1586364061
transform 1 0 36432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36064 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_387
timestamp 1586364061
transform 1 0 36708 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_395
timestamp 1586364061
transform 1 0 37444 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_388
timestamp 1586364061
transform 1 0 36800 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 36892 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37168 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _285_
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_400
timestamp 1586364061
transform 1 0 37904 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_399
timestamp 1586364061
transform 1 0 37812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 38088 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_404
timestamp 1586364061
transform 1 0 38272 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38640 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 38824 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 38640 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_423
timestamp 1586364061
transform 1 0 40020 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_419
timestamp 1586364061
transform 1 0 39652 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_425
timestamp 1586364061
transform 1 0 40204 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_421
timestamp 1586364061
transform 1 0 39836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_439
timestamp 1586364061
transform 1 0 41492 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_430
timestamp 1586364061
transform 1 0 40664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_443
timestamp 1586364061
transform 1 0 41860 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 41676 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_456
timestamp 1586364061
transform 1 0 43056 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_454
timestamp 1586364061
transform 1 0 42872 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_450
timestamp 1586364061
transform 1 0 42504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43240 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_458
timestamp 1586364061
transform 1 0 43240 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_461
timestamp 1586364061
transform 1 0 43516 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_460
timestamp 1586364061
transform 1 0 43424 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_469
timestamp 1586364061
transform 1 0 44252 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 866 592
use scs8hd_decap_8  FILLER_1_477
timestamp 1586364061
transform 1 0 44988 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_473
timestamp 1586364061
transform 1 0 44620 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_473
timestamp 1586364061
transform 1 0 44620 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44804 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44436 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_485
timestamp 1586364061
transform 1 0 45724 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_493
timestamp 1586364061
transform 1 0 46460 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_1_485
timestamp 1586364061
transform 1 0 45724 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 48852 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 48852 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_515
timestamp 1586364061
transform 1 0 48484 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__593__B
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_221
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_225
timestamp 1586364061
transform 1 0 21804 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _591_
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23920 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_250
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 28152 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27508 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_285
timestamp 1586364061
transform 1 0 27324 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_289
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _584_
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29348 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_309
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_317
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__266__B
timestamp 1586364061
transform 1 0 33120 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32660 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_327
timestamp 1586364061
transform 1 0 31188 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_340
timestamp 1586364061
transform 1 0 32384 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_345
timestamp 1586364061
transform 1 0 32844 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _266_
timestamp 1586364061
transform 1 0 33304 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 34868 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34684 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_359
timestamp 1586364061
transform 1 0 34132 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_378
timestamp 1586364061
transform 1 0 35880 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36064 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_382
timestamp 1586364061
transform 1 0 36248 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_389
timestamp 1586364061
transform 1 0 36892 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_393
timestamp 1586364061
transform 1 0 37260 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__285__B
timestamp 1586364061
transform 1 0 37076 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__281__B
timestamp 1586364061
transform 1 0 38088 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _281_
timestamp 1586364061
transform 1 0 38272 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 39836 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_413
timestamp 1586364061
transform 1 0 39100 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_417
timestamp 1586364061
transform 1 0 39468 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_432
timestamp 1586364061
transform 1 0 40848 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_438
timestamp 1586364061
transform 1 0 41400 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_450
timestamp 1586364061
transform 1 0 42504 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_468
timestamp 1586364061
transform 1 0 44160 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_472
timestamp 1586364061
transform 1 0 44528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_484
timestamp 1586364061
transform 1 0 45632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_496
timestamp 1586364061
transform 1 0 46736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_508
timestamp 1586364061
transform 1 0 47840 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 48852 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_nor2_4  _593_
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__593__A
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__592__A
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _592_
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__622__A
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_279
timestamp 1586364061
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_283
timestamp 1586364061
transform 1 0 27140 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_291
timestamp 1586364061
transform 1 0 27876 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_322
timestamp 1586364061
transform 1 0 30728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_319
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_315
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30544 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32660 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_335
timestamp 1586364061
transform 1 0 31924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_339
timestamp 1586364061
transform 1 0 32292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_352
timestamp 1586364061
transform 1 0 33488 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_356
timestamp 1586364061
transform 1 0 33856 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34040 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_360
timestamp 1586364061
transform 1 0 34224 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_373
timestamp 1586364061
transform 1 0 35420 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35144 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35604 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36156 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__292__A
timestamp 1586364061
transform 1 0 37996 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__292__B
timestamp 1586364061
transform 1 0 37628 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_377
timestamp 1586364061
transform 1 0 35788 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_390
timestamp 1586364061
transform 1 0 36984 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_396
timestamp 1586364061
transform 1 0 37536 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_399
timestamp 1586364061
transform 1 0 37812 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__289__A
timestamp 1586364061
transform 1 0 38456 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _289_
timestamp 1586364061
transform 1 0 38640 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_421
timestamp 1586364061
transform 1 0 39836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_417
timestamp 1586364061
transform 1 0 39468 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39652 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_425
timestamp 1586364061
transform 1 0 40204 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40020 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40756 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41768 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41216 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_434
timestamp 1586364061
transform 1 0 41032 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_438
timestamp 1586364061
transform 1 0 41400 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_451
timestamp 1586364061
transform 1 0 42596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_455
timestamp 1586364061
transform 1 0 42964 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43148 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_472
timestamp 1586364061
transform 1 0 44528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_468
timestamp 1586364061
transform 1 0 44160 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_483
timestamp 1586364061
transform 1 0 45540 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_479
timestamp 1586364061
transform 1 0 45172 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45356 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45724 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_487
timestamp 1586364061
transform 1 0 45908 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__590__B
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_236
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23552 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__592__B
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_267
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _622_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_293
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30360 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28520 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__583__B
timestamp 1586364061
transform 1 0 29532 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_307
timestamp 1586364061
transform 1 0 29348 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_311
timestamp 1586364061
transform 1 0 29716 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_317
timestamp 1586364061
transform 1 0 30268 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_321
timestamp 1586364061
transform 1 0 30636 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_325
timestamp 1586364061
transform 1 0 31004 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31188 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__582__B
timestamp 1586364061
transform 1 0 30820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_335
timestamp 1586364061
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_329
timestamp 1586364061
transform 1 0 31372 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_340
timestamp 1586364061
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__B
timestamp 1586364061
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_344
timestamp 1586364061
transform 1 0 32752 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__257__B
timestamp 1586364061
transform 1 0 33028 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 33580 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 35144 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35512 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_364
timestamp 1586364061
transform 1 0 34592 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_372
timestamp 1586364061
transform 1 0 35328 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _292_
timestamp 1586364061
transform 1 0 37996 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_376
timestamp 1586364061
transform 1 0 35696 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_389
timestamp 1586364061
transform 1 0 36892 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_3  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39560 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__289__B
timestamp 1586364061
transform 1 0 39008 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_410
timestamp 1586364061
transform 1 0 38824 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_414
timestamp 1586364061
transform 1 0 39192 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_427
timestamp 1586364061
transform 1 0 40388 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_433
timestamp 1586364061
transform 1 0 40940 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40756 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_438
timestamp 1586364061
transform 1 0 41400 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41768 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_449
timestamp 1586364061
transform 1 0 42412 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_444
timestamp 1586364061
transform 1 0 41952 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_455
timestamp 1586364061
transform 1 0 42964 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45172 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_482
timestamp 1586364061
transform 1 0 45448 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_494
timestamp 1586364061
transform 1 0 46552 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_506
timestamp 1586364061
transform 1 0 47656 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 48852 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_514
timestamp 1586364061
transform 1 0 48392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _590_
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__590__A
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27784 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28152 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_288
timestamp 1586364061
transform 1 0 27600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_292
timestamp 1586364061
transform 1 0 27968 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _583_
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__582__A
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__583__A
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_296
timestamp 1586364061
transform 1 0 28336 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_300
timestamp 1586364061
transform 1 0 28704 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _257_
timestamp 1586364061
transform 1 0 33028 0 1 4896
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 31004 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 32844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__A
timestamp 1586364061
transform 1 0 32200 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_336
timestamp 1586364061
transform 1 0 32016 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_340
timestamp 1586364061
transform 1 0 32384 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_344
timestamp 1586364061
transform 1 0 32752 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 35144 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_356
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_360
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36892 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_385
timestamp 1586364061
transform 1 0 36524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_398
timestamp 1586364061
transform 1 0 37720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_402
timestamp 1586364061
transform 1 0 38088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 38272 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _277_
timestamp 1586364061
transform 1 0 38456 0 1 4896
box -38 -48 866 592
use scs8hd_fill_2  FILLER_5_419
timestamp 1586364061
transform 1 0 39652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_415
timestamp 1586364061
transform 1 0 39284 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 39468 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_423
timestamp 1586364061
transform 1 0 40020 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42412 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40848 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 41860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40664 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_441
timestamp 1586364061
transform 1 0 41676 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_445
timestamp 1586364061
transform 1 0 42044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43700 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__631__A
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_457
timestamp 1586364061
transform 1 0 43148 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_461
timestamp 1586364061
transform 1 0 43516 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_472
timestamp 1586364061
transform 1 0 44528 0 1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_5_478
timestamp 1586364061
transform 1 0 45080 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_486
timestamp 1586364061
transform 1 0 45816 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _624_
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__624__A
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_223
timestamp 1586364061
transform 1 0 21620 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__589__A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_229
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__589__B
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _589_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_271
timestamp 1586364061
transform 1 0 26036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_288
timestamp 1586364061
transform 1 0 27600 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26772 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_292
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_294
timestamp 1586364061
transform 1 0 28152 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_290
timestamp 1586364061
transform 1 0 27784 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_303
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_299
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__581__A
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 28520 0 -1 5984
box -38 -48 1050 592
use scs8hd_buf_1  _581_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_316
timestamp 1586364061
transform 1 0 30176 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_313
timestamp 1586364061
transform 1 0 29900 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_309
timestamp 1586364061
transform 1 0 29532 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_309
timestamp 1586364061
transform 1 0 29532 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29992 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _582_
timestamp 1586364061
transform 1 0 30268 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 30544 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_331
timestamp 1586364061
transform 1 0 31556 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_330
timestamp 1586364061
transform 1 0 31464 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_326
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31740 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _585_
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_348
timestamp 1586364061
transform 1 0 33120 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_344
timestamp 1586364061
transform 1 0 32752 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_346
timestamp 1586364061
transform 1 0 32936 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__244__B
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 32936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_359
timestamp 1586364061
transform 1 0 34132 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_351
timestamp 1586364061
transform 1 0 33396 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _244_
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_370
timestamp 1586364061
transform 1 0 35144 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__248__B
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 34408 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35512 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_384
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_377
timestamp 1586364061
transform 1 0 35788 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36156 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_389
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_6_391
timestamp 1586364061
transform 1 0 37076 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_388
timestamp 1586364061
transform 1 0 36800 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_400
timestamp 1586364061
transform 1 0 37904 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_397
timestamp 1586364061
transform 1 0 37628 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 37720 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_411
timestamp 1586364061
transform 1 0 38916 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_407
timestamp 1586364061
transform 1 0 38548 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__277__B
timestamp 1586364061
transform 1 0 38732 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 38272 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _273_
timestamp 1586364061
transform 1 0 38456 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_419
timestamp 1586364061
transform 1 0 39652 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_415
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_426
timestamp 1586364061
transform 1 0 40296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39468 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 39284 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40480 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_442
timestamp 1586364061
transform 1 0 41768 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_430
timestamp 1586364061
transform 1 0 40664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 41032 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_453
timestamp 1586364061
transform 1 0 42780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_447
timestamp 1586364061
transform 1 0 42228 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_445
timestamp 1586364061
transform 1 0 42044 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 42044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_466
timestamp 1586364061
transform 1 0 43976 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_457
timestamp 1586364061
transform 1 0 43148 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43148 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_470
timestamp 1586364061
transform 1 0 44344 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_472
timestamp 1586364061
transform 1 0 44528 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_468
timestamp 1586364061
transform 1 0 44160 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44712 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44528 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44160 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 44712 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_481
timestamp 1586364061
transform 1 0 45356 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_477
timestamp 1586364061
transform 1 0 44988 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 45540 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45172 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _631_
timestamp 1586364061
transform 1 0 44896 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_485
timestamp 1586364061
transform 1 0 45724 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_491
timestamp 1586364061
transform 1 0 46276 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_485
timestamp 1586364061
transform 1 0 45724 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__630__A
timestamp 1586364061
transform 1 0 46092 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_inv_8  _630_
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 866 592
use scs8hd_decap_12  FILLER_7_502
timestamp 1586364061
transform 1 0 47288 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_498
timestamp 1586364061
transform 1 0 46920 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_503
timestamp 1586364061
transform 1 0 47380 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47104 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 48852 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 48852 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_515
timestamp 1586364061
transform 1 0 48484 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_514
timestamp 1586364061
transform 1 0 48392 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__625__A
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 590 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_293
timestamp 1586364061
transform 1 0 28060 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28796 0 -1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_310
timestamp 1586364061
transform 1 0 29624 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_314
timestamp 1586364061
transform 1 0 29992 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_318
timestamp 1586364061
transform 1 0 30360 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _234_
timestamp 1586364061
transform 1 0 32936 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__298__B
timestamp 1586364061
transform 1 0 32660 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_6  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_345
timestamp 1586364061
transform 1 0 32844 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _248_
timestamp 1586364061
transform 1 0 33948 0 -1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35512 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34960 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35328 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_366
timestamp 1586364061
transform 1 0 34776 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_370
timestamp 1586364061
transform 1 0 35144 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _267_
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_383
timestamp 1586364061
transform 1 0 36340 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_387
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_395
timestamp 1586364061
transform 1 0 37444 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_401
timestamp 1586364061
transform 1 0 37996 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38916 0 -1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__273__B
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_405
timestamp 1586364061
transform 1 0 38364 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_408
timestamp 1586364061
transform 1 0 38640 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_420
timestamp 1586364061
transform 1 0 39744 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 42044 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_437
timestamp 1586364061
transform 1 0 41308 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_441
timestamp 1586364061
transform 1 0 41676 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_448
timestamp 1586364061
transform 1 0 42320 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_456
timestamp 1586364061
transform 1 0 43056 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44896 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_468
timestamp 1586364061
transform 1 0 44160 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_473
timestamp 1586364061
transform 1 0 44620 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46460 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46092 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_485
timestamp 1586364061
transform 1 0 45724 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_491
timestamp 1586364061
transform 1 0 46276 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_496
timestamp 1586364061
transform 1 0 46736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_508
timestamp 1586364061
transform 1 0 47840 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 48852 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _625_
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__621__A
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_228
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_255
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__588__A
timestamp 1586364061
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _588_
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _623_
timestamp 1586364061
transform 1 0 26128 0 1 7072
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28152 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__623__A
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_285
timestamp 1586364061
transform 1 0 27324 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_292
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_300
timestamp 1586364061
transform 1 0 28704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_296
timestamp 1586364061
transform 1 0 28336 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28888 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28520 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_314
timestamp 1586364061
transform 1 0 29992 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29532 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29716 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30544 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30176 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30728 0 1 7072
box -38 -48 866 592
use scs8hd_nor2_4  _298_
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__298__A
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_331
timestamp 1586364061
transform 1 0 31556 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_339
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_356
timestamp 1586364061
transform 1 0 33856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_352
timestamp 1586364061
transform 1 0 33488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_360
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_371
timestamp 1586364061
transform 1 0 35236 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35052 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35512 0 1 7072
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 37536 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 37352 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36524 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_383
timestamp 1586364061
transform 1 0 36340 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_387
timestamp 1586364061
transform 1 0 36708 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_392
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_407
timestamp 1586364061
transform 1 0 38548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_411
timestamp 1586364061
transform 1 0 38916 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39100 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39284 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_418
timestamp 1586364061
transform 1 0 39560 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 39744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_422
timestamp 1586364061
transform 1 0 39928 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_426
timestamp 1586364061
transform 1 0 40296 0 1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_435
timestamp 1586364061
transform 1 0 41124 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_431
timestamp 1586364061
transform 1 0 40756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__628__A
timestamp 1586364061
transform 1 0 41308 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _628_
timestamp 1586364061
transform 1 0 41492 0 1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_9_448
timestamp 1586364061
transform 1 0 42320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_452
timestamp 1586364061
transform 1 0 42688 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42872 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__629__A
timestamp 1586364061
transform 1 0 42504 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43056 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44252 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45448 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 43792 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_459
timestamp 1586364061
transform 1 0 43332 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_463
timestamp 1586364061
transform 1 0 43700 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_466
timestamp 1586364061
transform 1 0 43976 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_480
timestamp 1586364061
transform 1 0 45264 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47104 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_484
timestamp 1586364061
transform 1 0 45632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_498
timestamp 1586364061
transform 1 0 46920 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_502
timestamp 1586364061
transform 1 0 47288 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_506
timestamp 1586364061
transform 1 0 47656 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 48852 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_514
timestamp 1586364061
transform 1 0 48392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _621_
timestamp 1586364061
transform 1 0 23184 0 -1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_236
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_257
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_289
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29624 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_302
timestamp 1586364061
transform 1 0 28888 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_321
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_325
timestamp 1586364061
transform 1 0 31004 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_330
timestamp 1586364061
transform 1 0 31464 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_342
timestamp 1586364061
transform 1 0 32568 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32292 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_346
timestamp 1586364061
transform 1 0 32936 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__295__B
timestamp 1586364061
transform 1 0 32752 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 33304 0 -1 8160
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__532__A
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__530__B
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__301__B
timestamp 1586364061
transform 1 0 36708 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__304__B
timestamp 1586364061
transform 1 0 36248 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_384
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_6  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38272 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 39376 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38732 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_407
timestamp 1586364061
transform 1 0 38548 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_411
timestamp 1586364061
transform 1 0 38916 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_415
timestamp 1586364061
transform 1 0 39284 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_427
timestamp 1586364061
transform 1 0 40388 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_8  _629_
timestamp 1586364061
transform 1 0 41676 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41400 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_435
timestamp 1586364061
transform 1 0 41124 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_440
timestamp 1586364061
transform 1 0 41584 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_450
timestamp 1586364061
transform 1 0 42504 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 43792 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44804 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__633__A
timestamp 1586364061
transform 1 0 44252 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_463
timestamp 1586364061
transform 1 0 43700 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_467
timestamp 1586364061
transform 1 0 44068 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_471
timestamp 1586364061
transform 1 0 44436 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46368 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 47380 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__632__A
timestamp 1586364061
transform 1 0 46092 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_484
timestamp 1586364061
transform 1 0 45632 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_488
timestamp 1586364061
transform 1 0 46000 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_491
timestamp 1586364061
transform 1 0 46276 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_495
timestamp 1586364061
transform 1 0 46644 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_8  FILLER_10_506
timestamp 1586364061
transform 1 0 47656 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 48852 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_514
timestamp 1586364061
transform 1 0 48392 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__627__A
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__620__A
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23736 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27508 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__595__B
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_279
timestamp 1586364061
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_283
timestamp 1586364061
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_290
timestamp 1586364061
transform 1 0 27784 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_294
timestamp 1586364061
transform 1 0 28152 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29532 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__595__A
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_320
timestamp 1586364061
transform 1 0 30544 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31280 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__295__A
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__533__A
timestamp 1586364061
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_324
timestamp 1586364061
transform 1 0 30912 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_337
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_341
timestamp 1586364061
transform 1 0 32476 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_344
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _532_
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_nor2_4  _533_
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__530__A
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_364
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _301_
timestamp 1586364061
transform 1 0 36708 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__304__A
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__301__A
timestamp 1586364061
transform 1 0 36524 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_382
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_396
timestamp 1586364061
transform 1 0 37536 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_400
timestamp 1586364061
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 38640 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_419
timestamp 1586364061
transform 1 0 39652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_423
timestamp 1586364061
transform 1 0 40020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_428
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41400 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41216 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_434
timestamp 1586364061
transform 1 0 41032 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_447
timestamp 1586364061
transform 1 0 42228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_451
timestamp 1586364061
transform 1 0 42596 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _633_
timestamp 1586364061
transform 1 0 44160 0 1 8160
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43148 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_460
timestamp 1586364061
transform 1 0 43424 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_477
timestamp 1586364061
transform 1 0 44988 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_482
timestamp 1586364061
transform 1 0 45448 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _632_
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45632 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47196 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_486
timestamp 1586364061
transform 1 0 45816 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_498
timestamp 1586364061
transform 1 0 46920 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_503
timestamp 1586364061
transform 1 0 47380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 48852 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_515
timestamp 1586364061
transform 1 0 48484 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _620_
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_8  _627_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_236
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__565__B
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__598__B
timestamp 1586364061
transform 1 0 25760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__561__B
timestamp 1586364061
transform 1 0 27692 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28060 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_287
timestamp 1586364061
transform 1 0 27508 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_291
timestamp 1586364061
transform 1 0 27876 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_295
timestamp 1586364061
transform 1 0 28244 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _595_
timestamp 1586364061
transform 1 0 28888 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_301
timestamp 1586364061
transform 1 0 28796 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_311
timestamp 1586364061
transform 1 0 29716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_315
timestamp 1586364061
transform 1 0 30084 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_322
timestamp 1586364061
transform 1 0 30728 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _295_
timestamp 1586364061
transform 1 0 32568 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_334
timestamp 1586364061
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_341
timestamp 1586364061
transform 1 0 32476 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _530_
timestamp 1586364061
transform 1 0 34408 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__533__B
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__532__B
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_355
timestamp 1586364061
transform 1 0 33764 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_371
timestamp 1586364061
transform 1 0 35236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_375
timestamp 1586364061
transform 1 0 35604 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _304_
timestamp 1586364061
transform 1 0 36064 0 -1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_379
timestamp 1586364061
transform 1 0 35972 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 39468 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_409
timestamp 1586364061
transform 1 0 38732 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_428
timestamp 1586364061
transform 1 0 40480 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_436
timestamp 1586364061
transform 1 0 41216 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_450
timestamp 1586364061
transform 1 0 42504 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_454
timestamp 1586364061
transform 1 0 42872 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_468
timestamp 1586364061
transform 1 0 44160 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_472
timestamp 1586364061
transform 1 0 44528 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45632 0 -1 9248
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 47196 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_493
timestamp 1586364061
transform 1 0 46460 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_504
timestamp 1586364061
transform 1 0 47472 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 48852 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 314 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 2430 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_189
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__626__A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _626_
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_221
timestamp 1586364061
transform 1 0 21436 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__568__A
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _568_
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_231
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_228
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__568__B
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_242
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__597__B
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__597__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _597_
timestamp 1586364061
transform 1 0 23736 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _565_
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_255
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__598__A
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__565__A
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _598_
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_279
timestamp 1586364061
transform 1 0 26772 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_277
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_284
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_284
timestamp 1586364061
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__561__A
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 27416 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 27508 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _561_
timestamp 1586364061
transform 1 0 27600 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_298
timestamp 1586364061
transform 1 0 28520 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_13_297
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__596__A
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_308
timestamp 1586364061
transform 1 0 29440 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__596__B
timestamp 1586364061
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__556__B
timestamp 1586364061
transform 1 0 29992 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _596_
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_319
timestamp 1586364061
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_315
timestamp 1586364061
transform 1 0 30084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__559__B
timestamp 1586364061
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__559__A
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _559_
timestamp 1586364061
transform 1 0 30176 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_329
timestamp 1586364061
transform 1 0 31372 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_325
timestamp 1586364061
transform 1 0 31004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_326
timestamp 1586364061
transform 1 0 31096 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__580__A
timestamp 1586364061
transform 1 0 31280 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _580_
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_335
timestamp 1586364061
transform 1 0 31924 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_337
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _233_
timestamp 1586364061
transform 1 0 31832 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_341
timestamp 1586364061
transform 1 0 32476 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_341
timestamp 1586364061
transform 1 0 32476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 32660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 32292 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _256_
timestamp 1586364061
transform 1 0 32844 0 1 9248
box -38 -48 314 592
use scs8hd_or2_4  _242_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 32844 0 -1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_13_348
timestamp 1586364061
transform 1 0 33120 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_352
timestamp 1586364061
transform 1 0 33488 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_356
timestamp 1586364061
transform 1 0 33856 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_352
timestamp 1586364061
transform 1 0 33488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__B
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_364
timestamp 1586364061
transform 1 0 34592 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_371
timestamp 1586364061
transform 1 0 35236 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__531__B
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__531__A
timestamp 1586364061
transform 1 0 35052 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _531_
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 35604 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_387
timestamp 1586364061
transform 1 0 36708 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_382
timestamp 1586364061
transform 1 0 36248 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_376
timestamp 1586364061
transform 1 0 35696 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36064 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 35788 0 1 9248
box -38 -48 1050 592
use scs8hd_buf_1  _265_
timestamp 1586364061
transform 1 0 36432 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_395
timestamp 1586364061
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_399
timestamp 1586364061
transform 1 0 37812 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_392
timestamp 1586364061
transform 1 0 37168 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_388
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _280_
timestamp 1586364061
transform 1 0 37536 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_402
timestamp 1586364061
transform 1 0 38088 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37904 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 37996 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_410
timestamp 1586364061
transform 1 0 38824 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39008 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38548 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38548 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_416
timestamp 1586364061
transform 1 0 39376 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_13_418
timestamp 1586364061
transform 1 0 39560 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_414
timestamp 1586364061
transform 1 0 39192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39376 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_426
timestamp 1586364061
transform 1 0 40296 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__538__A
timestamp 1586364061
transform 1 0 40112 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _538_
timestamp 1586364061
transform 1 0 40112 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_437
timestamp 1586364061
transform 1 0 41308 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_433
timestamp 1586364061
transform 1 0 40940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_439
timestamp 1586364061
transform 1 0 41492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_435
timestamp 1586364061
transform 1 0 41124 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_431
timestamp 1586364061
transform 1 0 40756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41124 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__538__B
timestamp 1586364061
transform 1 0 40940 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_443
timestamp 1586364061
transform 1 0 41860 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42412 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_450
timestamp 1586364061
transform 1 0 42504 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_459
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_462
timestamp 1586364061
transform 1 0 43608 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_458
timestamp 1586364061
transform 1 0 43240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43424 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43976 0 1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_473
timestamp 1586364061
transform 1 0 44620 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_13_479
timestamp 1586364061
transform 1 0 45172 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_475
timestamp 1586364061
transform 1 0 44804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44988 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__635__A
timestamp 1586364061
transform 1 0 45448 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_485
timestamp 1586364061
transform 1 0 45724 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_484
timestamp 1586364061
transform 1 0 45632 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _635_
timestamp 1586364061
transform 1 0 45908 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_496
timestamp 1586364061
transform 1 0 46736 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_502
timestamp 1586364061
transform 1 0 47288 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_498
timestamp 1586364061
transform 1 0 46920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 47104 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_507
timestamp 1586364061
transform 1 0 47748 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_13_506
timestamp 1586364061
transform 1 0 47656 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 47472 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 47472 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 48852 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 48852 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_514
timestamp 1586364061
transform 1 0 48392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_515
timestamp 1586364061
transform 1 0 48484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 130 592
use scs8hd_clkbuf_1  clkbuf_1_0_0_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_212
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_216
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_251
timestamp 1586364061
transform 1 0 24196 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26312 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 27416 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_277
timestamp 1586364061
transform 1 0 26588 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_282
timestamp 1586364061
transform 1 0 27048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__560__B
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__560__A
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_buf_1  _243_
timestamp 1586364061
transform 1 0 29348 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_314
timestamp 1586364061
transform 1 0 29992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_310
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 29808 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 30176 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 32108 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 31924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__556__A
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_329
timestamp 1586364061
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_333
timestamp 1586364061
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_348
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_352
timestamp 1586364061
transform 1 0 33488 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__290__B
timestamp 1586364061
transform 1 0 33304 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_356
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__290__A
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__534__B
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__534__A
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_buf_1  _261_
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_370
timestamp 1586364061
transform 1 0 35144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 35328 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_374
timestamp 1586364061
transform 1 0 35512 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 37628 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__291__A
timestamp 1586364061
transform 1 0 37260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_395
timestamp 1586364061
transform 1 0 37444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_410
timestamp 1586364061
transform 1 0 38824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_414
timestamp 1586364061
transform 1 0 39192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39376 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_418
timestamp 1586364061
transform 1 0 39560 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_423
timestamp 1586364061
transform 1 0 40020 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_428
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42596 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 40848 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 40664 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_443
timestamp 1586364061
transform 1 0 41860 0 1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_15_454
timestamp 1586364061
transform 1 0 42872 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43884 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43700 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44896 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_458
timestamp 1586364061
transform 1 0 43240 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_461
timestamp 1586364061
transform 1 0 43516 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_474
timestamp 1586364061
transform 1 0 44712 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_478
timestamp 1586364061
transform 1 0 45080 0 1 10336
box -38 -48 406 592
use scs8hd_inv_8  _634_
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__634__A
timestamp 1586364061
transform 1 0 45816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_484
timestamp 1586364061
transform 1 0 45632 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_498
timestamp 1586364061
transform 1 0 46920 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 48852 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_510
timestamp 1586364061
transform 1 0 48024 0 1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21620 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_219
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_245
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28060 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_281
timestamp 1586364061
transform 1 0 26956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_291
timestamp 1586364061
transform 1 0 27876 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_295
timestamp 1586364061
transform 1 0 28244 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _556_
timestamp 1586364061
transform 1 0 30176 0 -1 11424
box -38 -48 866 592
use scs8hd_nor2_4  _560_
timestamp 1586364061
transform 1 0 28612 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29900 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_308
timestamp 1586364061
transform 1 0 29440 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_315
timestamp 1586364061
transform 1 0 30084 0 -1 11424
box -38 -48 130 592
use scs8hd_or2_4  _290_
timestamp 1586364061
transform 1 0 32844 0 -1 11424
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__255__B
timestamp 1586364061
transform 1 0 31556 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__B
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_325
timestamp 1586364061
transform 1 0 31004 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  FILLER_16_333
timestamp 1586364061
transform 1 0 31740 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_343
timestamp 1586364061
transform 1 0 32660 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _534_
timestamp 1586364061
transform 1 0 34960 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 33856 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_352
timestamp 1586364061
transform 1 0 33488 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_358
timestamp 1586364061
transform 1 0 34040 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_366
timestamp 1586364061
transform 1 0 34776 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _291_
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__542__B
timestamp 1586364061
transform 1 0 37168 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37904 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_4  FILLER_16_388
timestamp 1586364061
transform 1 0 36800 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_394
timestamp 1586364061
transform 1 0 37352 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_402
timestamp 1586364061
transform 1 0 38088 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38548 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__539__A
timestamp 1586364061
transform 1 0 40480 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_416
timestamp 1586364061
transform 1 0 39376 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_426
timestamp 1586364061
transform 1 0 40296 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 40664 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42136 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_441
timestamp 1586364061
transform 1 0 41676 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_445
timestamp 1586364061
transform 1 0 42044 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_448
timestamp 1586364061
transform 1 0 42320 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_456
timestamp 1586364061
transform 1 0 43056 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45448 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_459
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_463
timestamp 1586364061
transform 1 0 43700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_473
timestamp 1586364061
transform 1 0 44620 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_481
timestamp 1586364061
transform 1 0 45356 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_485
timestamp 1586364061
transform 1 0 45724 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_497
timestamp 1586364061
transform 1 0 46828 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_509
timestamp 1586364061
transform 1 0 47932 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 48852 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_515
timestamp 1586364061
transform 1 0 48484 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _567_
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__567__A
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__567__B
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_219
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__566__A
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27784 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__566__B
timestamp 1586364061
transform 1 0 26220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28152 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_271
timestamp 1586364061
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_288
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_292
timestamp 1586364061
transform 1 0 27968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_301
timestamp 1586364061
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_296
timestamp 1586364061
transform 1 0 28336 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_310
timestamp 1586364061
transform 1 0 29624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29716 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29900 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_322
timestamp 1586364061
transform 1 0 30728 0 1 11424
box -38 -48 222 592
use scs8hd_or2_4  _255_
timestamp 1586364061
transform 1 0 31556 0 1 11424
box -38 -48 682 592
use scs8hd_or2_4  _260_
timestamp 1586364061
transform 1 0 32936 0 1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 32476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 31372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_326
timestamp 1586364061
transform 1 0 31096 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_338
timestamp 1586364061
transform 1 0 32200 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_343
timestamp 1586364061
transform 1 0 32660 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _535_
timestamp 1586364061
transform 1 0 34960 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__279__B
timestamp 1586364061
transform 1 0 34132 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__535__A
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_353
timestamp 1586364061
transform 1 0 33580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_357
timestamp 1586364061
transform 1 0 33948 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_361
timestamp 1586364061
transform 1 0 34316 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _542_
timestamp 1586364061
transform 1 0 37168 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__288__A
timestamp 1586364061
transform 1 0 36616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__A
timestamp 1586364061
transform 1 0 36984 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__529__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_385
timestamp 1586364061
transform 1 0 36524 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_388
timestamp 1586364061
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_401
timestamp 1586364061
transform 1 0 37996 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_405
timestamp 1586364061
transform 1 0 38364 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__537__A
timestamp 1586364061
transform 1 0 38640 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _537_
timestamp 1586364061
transform 1 0 38824 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_419
timestamp 1586364061
transform 1 0 39652 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__539__B
timestamp 1586364061
transform 1 0 39836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_423
timestamp 1586364061
transform 1 0 40020 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _539_
timestamp 1586364061
transform 1 0 40480 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42136 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41952 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41584 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_437
timestamp 1586364061
transform 1 0 41308 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_442
timestamp 1586364061
transform 1 0 41768 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_455
timestamp 1586364061
transform 1 0 42964 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43700 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45264 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_459
timestamp 1586364061
transform 1 0 43332 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_472
timestamp 1586364061
transform 1 0 44528 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_482
timestamp 1586364061
transform 1 0 45448 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__608__A
timestamp 1586364061
transform 1 0 46828 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45632 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_486
timestamp 1586364061
transform 1 0 45816 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_489
timestamp 1586364061
transform 1 0 46092 0 1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_17_499
timestamp 1586364061
transform 1 0 47012 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 48852 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_511
timestamp 1586364061
transform 1 0 48116 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_515
timestamp 1586364061
transform 1 0 48484 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_clkbuf_16  clkbuf_0_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 1878 592
use scs8hd_decap_8  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _566_
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__572__B
timestamp 1586364061
transform 1 0 25944 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_280
timestamp 1586364061
transform 1 0 26864 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_291
timestamp 1586364061
transform 1 0 27876 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_295
timestamp 1586364061
transform 1 0 28244 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28612 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29900 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_298
timestamp 1586364061
transform 1 0 28520 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_302
timestamp 1586364061
transform 1 0 28888 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_308
timestamp 1586364061
transform 1 0 29440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_322
timestamp 1586364061
transform 1 0 30728 0 -1 12512
box -38 -48 1142 592
use scs8hd_or2_4  _264_
timestamp 1586364061
transform 1 0 32476 0 -1 12512
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_334
timestamp 1586364061
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_348
timestamp 1586364061
transform 1 0 33120 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_352
timestamp 1586364061
transform 1 0 33488 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__293__A
timestamp 1586364061
transform 1 0 33672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__B
timestamp 1586364061
transform 1 0 33304 0 -1 12512
box -38 -48 222 592
use scs8hd_or2_4  _279_
timestamp 1586364061
transform 1 0 33856 0 -1 12512
box -38 -48 682 592
use scs8hd_fill_2  FILLER_18_363
timestamp 1586364061
transform 1 0 34500 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_371
timestamp 1586364061
transform 1 0 35236 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_367
timestamp 1586364061
transform 1 0 34868 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__287__B
timestamp 1586364061
transform 1 0 35052 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__283__B
timestamp 1586364061
transform 1 0 34684 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__535__B
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _529_
timestamp 1586364061
transform 1 0 35604 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_1  _288_
timestamp 1586364061
transform 1 0 36616 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 37812 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__543__B
timestamp 1586364061
transform 1 0 36064 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__540__B
timestamp 1586364061
transform 1 0 37444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_378
timestamp 1586364061
transform 1 0 35880 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_382
timestamp 1586364061
transform 1 0 36248 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_18_389
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40388 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__537__B
timestamp 1586364061
transform 1 0 39008 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_410
timestamp 1586364061
transform 1 0 38824 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_414
timestamp 1586364061
transform 1 0 39192 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_422
timestamp 1586364061
transform 1 0 39928 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42596 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_438
timestamp 1586364061
transform 1 0 41400 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_449
timestamp 1586364061
transform 1 0 42412 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_453
timestamp 1586364061
transform 1 0 42780 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_466
timestamp 1586364061
transform 1 0 43976 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_462
timestamp 1586364061
transform 1 0 43608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_457
timestamp 1586364061
transform 1 0 43148 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43792 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_470
timestamp 1586364061
transform 1 0 44344 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44160 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45080 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45264 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_8  _608_
timestamp 1586364061
transform 1 0 46828 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_489
timestamp 1586364061
transform 1 0 46092 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_506
timestamp 1586364061
transform 1 0 47656 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 48852 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_514
timestamp 1586364061
transform 1 0 48392 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 2430 592
use scs8hd_fill_1  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 1050 592
use scs8hd_conb_1  _636_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__563__A
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__563__B
timestamp 1586364061
transform 1 0 21804 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_222
timestamp 1586364061
transform 1 0 21528 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _563_
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_240
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_255
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_252
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__562__A
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_1  _562_
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_267
timestamp 1586364061
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__572__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _572_
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_285
timestamp 1586364061
transform 1 0 27324 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_283
timestamp 1586364061
transform 1 0 27140 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_279
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__557__B
timestamp 1586364061
transform 1 0 27600 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__557__A
timestamp 1586364061
transform 1 0 27416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _557_
timestamp 1586364061
transform 1 0 27600 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_290
timestamp 1586364061
transform 1 0 27784 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_307
timestamp 1586364061
transform 1 0 29348 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_301
timestamp 1586364061
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_297
timestamp 1586364061
transform 1 0 28428 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 28336 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_315
timestamp 1586364061
transform 1 0 30084 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_315
timestamp 1586364061
transform 1 0 30084 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__555__A
timestamp 1586364061
transform 1 0 29532 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30176 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_319
timestamp 1586364061
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30636 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_329
timestamp 1586364061
transform 1 0 31372 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_325
timestamp 1586364061
transform 1 0 31004 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_326
timestamp 1586364061
transform 1 0 31096 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_337
timestamp 1586364061
transform 1 0 32108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_336
timestamp 1586364061
transform 1 0 32016 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__294__A
timestamp 1586364061
transform 1 0 32108 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_341
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 32752 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _294_
timestamp 1586364061
transform 1 0 32292 0 1 12512
box -38 -48 314 592
use scs8hd_or2_4  _275_
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 682 592
use scs8hd_fill_2  FILLER_19_346
timestamp 1586364061
transform 1 0 32936 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__B
timestamp 1586364061
transform 1 0 33120 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_353
timestamp 1586364061
transform 1 0 33580 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_349
timestamp 1586364061
transform 1 0 33212 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__303__A
timestamp 1586364061
transform 1 0 33764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__302__A
timestamp 1586364061
transform 1 0 33396 0 -1 13600
box -38 -48 222 592
use scs8hd_or2_4  _293_
timestamp 1586364061
transform 1 0 33304 0 1 12512
box -38 -48 682 592
use scs8hd_fill_1  FILLER_20_361
timestamp 1586364061
transform 1 0 34316 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_357
timestamp 1586364061
transform 1 0 33948 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_361
timestamp 1586364061
transform 1 0 34316 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_357
timestamp 1586364061
transform 1 0 33948 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__293__B
timestamp 1586364061
transform 1 0 34132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__D
timestamp 1586364061
transform 1 0 34408 0 -1 13600
box -38 -48 222 592
use scs8hd_or2_4  _283_
timestamp 1586364061
transform 1 0 34592 0 -1 13600
box -38 -48 682 592
use scs8hd_fill_2  FILLER_20_371
timestamp 1586364061
transform 1 0 35236 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_or2_4  _287_
timestamp 1586364061
transform 1 0 35052 0 1 12512
box -38 -48 682 592
use scs8hd_decap_4  FILLER_20_375
timestamp 1586364061
transform 1 0 35604 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__296__A
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_380
timestamp 1586364061
transform 1 0 36064 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_376
timestamp 1586364061
transform 1 0 35696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__A
timestamp 1586364061
transform 1 0 36248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 35880 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _543_
timestamp 1586364061
transform 1 0 35972 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_1  _284_
timestamp 1586364061
transform 1 0 36432 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_392
timestamp 1586364061
transform 1 0 37168 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_388
timestamp 1586364061
transform 1 0 36800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_387
timestamp 1586364061
transform 1 0 36708 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36984 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__536__A
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _536_
timestamp 1586364061
transform 1 0 37444 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_398
timestamp 1586364061
transform 1 0 37720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_396
timestamp 1586364061
transform 1 0 37536 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_402
timestamp 1586364061
transform 1 0 38088 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_398
timestamp 1586364061
transform 1 0 37720 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__540__A
timestamp 1586364061
transform 1 0 37904 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _540_
timestamp 1586364061
transform 1 0 37904 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_413
timestamp 1586364061
transform 1 0 39100 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_409
timestamp 1586364061
transform 1 0 38732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38916 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 38640 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_20_420
timestamp 1586364061
transform 1 0 39744 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_423
timestamp 1586364061
transform 1 0 40020 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_419
timestamp 1586364061
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__541__B
timestamp 1586364061
transform 1 0 40296 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 39836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _276_
timestamp 1586364061
transform 1 0 39468 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40480 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _541_
timestamp 1586364061
transform 1 0 40480 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_439
timestamp 1586364061
transform 1 0 41492 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_437
timestamp 1586364061
transform 1 0 41308 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__541__A
timestamp 1586364061
transform 1 0 41492 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_443
timestamp 1586364061
transform 1 0 41860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_441
timestamp 1586364061
transform 1 0 41676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41860 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_450
timestamp 1586364061
transform 1 0 42504 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_454
timestamp 1586364061
transform 1 0 42872 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43056 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_459
timestamp 1586364061
transform 1 0 43332 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_458
timestamp 1586364061
transform 1 0 43240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43424 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_471
timestamp 1586364061
transform 1 0 44436 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_475
timestamp 1586364061
transform 1 0 44804 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_471
timestamp 1586364061
transform 1 0 44436 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_481
timestamp 1586364061
transform 1 0 45356 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45172 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45172 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_492
timestamp 1586364061
transform 1 0 46368 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_488
timestamp 1586364061
transform 1 0 46000 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_485
timestamp 1586364061
transform 1 0 45724 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46184 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_505
timestamp 1586364061
transform 1 0 47564 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_502
timestamp 1586364061
transform 1 0 47288 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_498
timestamp 1586364061
transform 1 0 46920 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__609__A
timestamp 1586364061
transform 1 0 47104 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _609_
timestamp 1586364061
transform 1 0 46736 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 48852 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 48852 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_514
timestamp 1586364061
transform 1 0 48392 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_513
timestamp 1586364061
transform 1 0 48300 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use scs8hd_clkbuf_1  clkbuf_1_1_0_clk
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 2430 592
use scs8hd_decap_4  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_221
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_249
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27784 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_288
timestamp 1586364061
transform 1 0 27600 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_292
timestamp 1586364061
transform 1 0 27968 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_21_302
timestamp 1586364061
transform 1 0 28888 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_298
timestamp 1586364061
transform 1 0 28520 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__569__B
timestamp 1586364061
transform 1 0 28336 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__569__A
timestamp 1586364061
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use scs8hd_buf_1  _555_
timestamp 1586364061
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_316
timestamp 1586364061
transform 1 0 30176 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_313
timestamp 1586364061
transform 1 0 29900 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_309
timestamp 1586364061
transform 1 0 29532 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__558__A
timestamp 1586364061
transform 1 0 29992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 30360 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 30544 0 1 13600
box -38 -48 1050 592
use scs8hd_or2_4  _271_
timestamp 1586364061
transform 1 0 32292 0 1 13600
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 33120 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__271__B
timestamp 1586364061
transform 1 0 32108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__558__B
timestamp 1586364061
transform 1 0 31740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_331
timestamp 1586364061
transform 1 0 31556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_335
timestamp 1586364061
transform 1 0 31924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_346
timestamp 1586364061
transform 1 0 32936 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _296_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 34868 0 1 13600
box -38 -48 866 592
use scs8hd_buf_1  _303_
timestamp 1586364061
transform 1 0 33672 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__296__C
timestamp 1586364061
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__302__B
timestamp 1586364061
transform 1 0 33488 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_350
timestamp 1586364061
transform 1 0 33304 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_357
timestamp 1586364061
transform 1 0 33948 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_362
timestamp 1586364061
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 36984 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 36800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__B
timestamp 1586364061
transform 1 0 35880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 36248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_376
timestamp 1586364061
transform 1 0 35696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_380
timestamp 1586364061
transform 1 0 36064 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_384
timestamp 1586364061
transform 1 0 36432 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_401
timestamp 1586364061
transform 1 0 37996 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_405
timestamp 1586364061
transform 1 0 38364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 38180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38548 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _272_
timestamp 1586364061
transform 1 0 38732 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_412
timestamp 1586364061
transform 1 0 39008 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 39192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_416
timestamp 1586364061
transform 1 0 39376 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_420
timestamp 1586364061
transform 1 0 39744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39560 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_424
timestamp 1586364061
transform 1 0 40112 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39928 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__A
timestamp 1586364061
transform 1 0 43056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_431
timestamp 1586364061
transform 1 0 40756 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_435
timestamp 1586364061
transform 1 0 41124 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_449
timestamp 1586364061
transform 1 0 42412 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_453
timestamp 1586364061
transform 1 0 42780 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43424 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45080 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45448 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_458
timestamp 1586364061
transform 1 0 43240 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_471
timestamp 1586364061
transform 1 0 44436 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_475
timestamp 1586364061
transform 1 0 44804 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_480
timestamp 1586364061
transform 1 0 45264 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 46368 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 46828 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47196 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_484
timestamp 1586364061
transform 1 0 45632 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_21_489
timestamp 1586364061
transform 1 0 46092 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_495
timestamp 1586364061
transform 1 0 46644 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_499
timestamp 1586364061
transform 1 0 47012 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_503
timestamp 1586364061
transform 1 0 47380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 48852 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_515
timestamp 1586364061
transform 1 0 48484 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 2430 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24748 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_249
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_289
timestamp 1586364061
transform 1 0 27692 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_293
timestamp 1586364061
transform 1 0 28060 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _558_
timestamp 1586364061
transform 1 0 30268 0 -1 14688
box -38 -48 866 592
use scs8hd_nor2_4  _569_
timestamp 1586364061
transform 1 0 28704 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29716 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_296
timestamp 1586364061
transform 1 0 28336 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_309
timestamp 1586364061
transform 1 0 29532 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_313
timestamp 1586364061
transform 1 0 29900 0 -1 14688
box -38 -48 406 592
use scs8hd_or2_4  _302_
timestamp 1586364061
transform 1 0 32844 0 -1 14688
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_326
timestamp 1586364061
transform 1 0 31096 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_334
timestamp 1586364061
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_337
timestamp 1586364061
transform 1 0 32108 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_8  _235_
timestamp 1586364061
transform 1 0 34408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__246__B
timestamp 1586364061
transform 1 0 35420 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__C
timestamp 1586364061
transform 1 0 33672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__250__A
timestamp 1586364061
transform 1 0 34040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_352
timestamp 1586364061
transform 1 0 33488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_356
timestamp 1586364061
transform 1 0 33856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_360
timestamp 1586364061
transform 1 0 34224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_371
timestamp 1586364061
transform 1 0 35236 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_375
timestamp 1586364061
transform 1 0 35604 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _247_
timestamp 1586364061
transform 1 0 35972 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 37812 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__300__A
timestamp 1586364061
transform 1 0 36432 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__546__A
timestamp 1586364061
transform 1 0 36892 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_382
timestamp 1586364061
transform 1 0 36248 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_386
timestamp 1586364061
transform 1 0 36616 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_391
timestamp 1586364061
transform 1 0 37076 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_398
timestamp 1586364061
transform 1 0 37720 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39560 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40572 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_410
timestamp 1586364061
transform 1 0 38824 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_427
timestamp 1586364061
transform 1 0 40388 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_431
timestamp 1586364061
transform 1 0 40756 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_438
timestamp 1586364061
transform 1 0 41400 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_442
timestamp 1586364061
transform 1 0 41768 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41584 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_453
timestamp 1586364061
transform 1 0 42780 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_449
timestamp 1586364061
transform 1 0 42412 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42596 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _607_
timestamp 1586364061
transform 1 0 43424 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45080 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_459
timestamp 1586364061
transform 1 0 43332 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_469
timestamp 1586364061
transform 1 0 44252 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_477
timestamp 1586364061
transform 1 0 44988 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46644 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 46092 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46460 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_487
timestamp 1586364061
transform 1 0 45908 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_491
timestamp 1586364061
transform 1 0 46276 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_498
timestamp 1586364061
transform 1 0 46920 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 48852 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_510
timestamp 1586364061
transform 1 0 48024 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__312__A
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__312__B
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_200
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _564_
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__564__A
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__564__B
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__612__A
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__571__B
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__571__A
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_265
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__570__B
timestamp 1586364061
transform 1 0 27968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_270
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_285
timestamp 1586364061
transform 1 0 27324 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_289
timestamp 1586364061
transform 1 0 27692 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29256 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__570__A
timestamp 1586364061
transform 1 0 28612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_297
timestamp 1586364061
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_301
timestamp 1586364061
transform 1 0 28796 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_317
timestamp 1586364061
transform 1 0 30268 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30820 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_328
timestamp 1586364061
transform 1 0 31280 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 31464 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_332
timestamp 1586364061
transform 1 0 31648 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 32016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_341
timestamp 1586364061
transform 1 0 32476 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _236_
timestamp 1586364061
transform 1 0 32200 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_345
timestamp 1586364061
transform 1 0 32844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 32660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__D
timestamp 1586364061
transform 1 0 33028 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _246_
timestamp 1586364061
transform 1 0 34868 0 1 14688
box -38 -48 866 592
use scs8hd_or4_4  _249_
timestamp 1586364061
transform 1 0 33212 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__299__B
timestamp 1586364061
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__C
timestamp 1586364061
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_358
timestamp 1586364061
transform 1 0 34040 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_362
timestamp 1586364061
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_384
timestamp 1586364061
transform 1 0 36432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_380
timestamp 1586364061
transform 1 0 36064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_376
timestamp 1586364061
transform 1 0 35696 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__D
timestamp 1586364061
transform 1 0 36248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 35880 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_388
timestamp 1586364061
transform 1 0 36800 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__299__A
timestamp 1586364061
transform 1 0 36616 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _546_
timestamp 1586364061
transform 1 0 36892 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_402
timestamp 1586364061
transform 1 0 38088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_398
timestamp 1586364061
transform 1 0 37720 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__545__A
timestamp 1586364061
transform 1 0 37904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_409
timestamp 1586364061
transform 1 0 38732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__545__B
timestamp 1586364061
transform 1 0 38272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 38916 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _278_
timestamp 1586364061
transform 1 0 38456 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_419
timestamp 1586364061
transform 1 0 39652 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_413
timestamp 1586364061
transform 1 0 39100 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39468 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_423
timestamp 1586364061
transform 1 0 40020 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 14688
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42044 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__604__A
timestamp 1586364061
transform 1 0 41584 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_437
timestamp 1586364061
transform 1 0 41308 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_442
timestamp 1586364061
transform 1 0 41768 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_448
timestamp 1586364061
transform 1 0 42320 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_452
timestamp 1586364061
transform 1 0 42688 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_455
timestamp 1586364061
transform 1 0 42964 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43148 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44804 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_468
timestamp 1586364061
transform 1 0 44160 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_472
timestamp 1586364061
transform 1 0 44528 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_480
timestamp 1586364061
transform 1 0 45264 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45724 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 47288 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_484
timestamp 1586364061
transform 1 0 45632 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_487
timestamp 1586364061
transform 1 0 45908 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_498
timestamp 1586364061
transform 1 0 46920 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_504
timestamp 1586364061
transform 1 0 47472 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 48852 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _312_
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__310__B
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _612_
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_225
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_233
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _571_
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_260
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_264
timestamp 1586364061
transform 1 0 25392 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_272
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_285
timestamp 1586364061
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_289
timestamp 1586364061
transform 1 0 27692 0 -1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _570_
timestamp 1586364061
transform 1 0 28796 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_310
timestamp 1586364061
transform 1 0 29624 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_314
timestamp 1586364061
transform 1 0 29992 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_322
timestamp 1586364061
transform 1 0 30728 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_8  _238_
timestamp 1586364061
transform 1 0 32108 0 -1 15776
box -38 -48 866 592
use scs8hd_buf_1  _239_
timestamp 1586364061
transform 1 0 31004 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__241__C
timestamp 1586364061
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 31464 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_328
timestamp 1586364061
transform 1 0 31280 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_332
timestamp 1586364061
transform 1 0 31648 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_346
timestamp 1586364061
transform 1 0 32936 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_355
timestamp 1586364061
transform 1 0 33764 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_351
timestamp 1586364061
transform 1 0 33396 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__B
timestamp 1586364061
transform 1 0 33580 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__A
timestamp 1586364061
transform 1 0 33212 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _250_
timestamp 1586364061
transform 1 0 33856 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_363
timestamp 1586364061
transform 1 0 34500 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_359
timestamp 1586364061
transform 1 0 34132 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__D
timestamp 1586364061
transform 1 0 34316 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__C
timestamp 1586364061
transform 1 0 34684 0 -1 15776
box -38 -48 222 592
use scs8hd_or4_4  _299_
timestamp 1586364061
transform 1 0 34868 0 -1 15776
box -38 -48 866 592
use scs8hd_buf_1  _300_
timestamp 1586364061
transform 1 0 36432 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _545_
timestamp 1586364061
transform 1 0 37720 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__546__B
timestamp 1586364061
transform 1 0 36892 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_376
timestamp 1586364061
transform 1 0 35696 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_387
timestamp 1586364061
transform 1 0 36708 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_391
timestamp 1586364061
transform 1 0 37076 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39836 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38732 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_407
timestamp 1586364061
transform 1 0 38548 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_411
timestamp 1586364061
transform 1 0 38916 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_419
timestamp 1586364061
transform 1 0 39652 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _604_
timestamp 1586364061
transform 1 0 41584 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_430
timestamp 1586364061
transform 1 0 40664 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_434
timestamp 1586364061
transform 1 0 41032 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_437
timestamp 1586364061
transform 1 0 41308 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_449
timestamp 1586364061
transform 1 0 42412 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_457
timestamp 1586364061
transform 1 0 43148 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_468
timestamp 1586364061
transform 1 0 44160 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_480
timestamp 1586364061
transform 1 0 45264 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 47288 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45724 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46736 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_484
timestamp 1586364061
transform 1 0 45632 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_494
timestamp 1586364061
transform 1 0 46552 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_498
timestamp 1586364061
transform 1 0 46920 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_505
timestamp 1586364061
transform 1 0 47564 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 48852 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_513
timestamp 1586364061
transform 1 0 48300 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _311_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__311__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__310__A
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_167
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__A
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__B
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_235
timestamp 1586364061
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _639_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__614__A
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_248
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28244 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_271
timestamp 1586364061
transform 1 0 26036 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_287
timestamp 1586364061
transform 1 0 27508 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_291
timestamp 1586364061
transform 1 0 27876 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_301
timestamp 1586364061
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_297
timestamp 1586364061
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_306
timestamp 1586364061
transform 1 0 29256 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29348 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_320
timestamp 1586364061
transform 1 0 30544 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_316
timestamp 1586364061
transform 1 0 30176 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30360 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 30728 0 1 15776
box -38 -48 222 592
use scs8hd_or3_4  _259_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 32108 0 1 15776
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30912 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 33120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__B
timestamp 1586364061
transform 1 0 31924 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__B
timestamp 1586364061
transform 1 0 31556 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_327
timestamp 1586364061
transform 1 0 31188 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_333
timestamp 1586364061
transform 1 0 31740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_346
timestamp 1586364061
transform 1 0 32936 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_350
timestamp 1586364061
transform 1 0 33304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__C
timestamp 1586364061
transform 1 0 33488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_354
timestamp 1586364061
transform 1 0 33672 0 1 15776
box -38 -48 130 592
use scs8hd_buf_1  _297_
timestamp 1586364061
transform 1 0 33764 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_358
timestamp 1586364061
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_362
timestamp 1586364061
transform 1 0 34408 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__297__A
timestamp 1586364061
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_367
timestamp 1586364061
transform 1 0 34868 0 1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use scs8hd_buf_1  _327_
timestamp 1586364061
transform 1 0 34960 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_371
timestamp 1586364061
transform 1 0 35236 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_375
timestamp 1586364061
transform 1 0 35604 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 35420 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _544_
timestamp 1586364061
transform 1 0 36340 0 1 15776
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 37904 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 37352 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__327__A
timestamp 1586364061
transform 1 0 35788 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__A
timestamp 1586364061
transform 1 0 36156 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_379
timestamp 1586364061
transform 1 0 35972 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_392
timestamp 1586364061
transform 1 0 37168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_396
timestamp 1586364061
transform 1 0 37536 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__512__A
timestamp 1586364061
transform 1 0 39560 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__512__B
timestamp 1586364061
transform 1 0 39192 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_411
timestamp 1586364061
transform 1 0 38916 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_416
timestamp 1586364061
transform 1 0 39376 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_420
timestamp 1586364061
transform 1 0 39744 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_424
timestamp 1586364061
transform 1 0 40112 0 1 15776
box -38 -48 130 592
use scs8hd_inv_8  _605_
timestamp 1586364061
transform 1 0 42044 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41860 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__605__A
timestamp 1586364061
transform 1 0 41492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_437
timestamp 1586364061
transform 1 0 41308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_441
timestamp 1586364061
transform 1 0 41676 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_454
timestamp 1586364061
transform 1 0 42872 0 1 15776
box -38 -48 406 592
use scs8hd_inv_8  _606_
timestamp 1586364061
transform 1 0 43608 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 44620 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__610__A
timestamp 1586364061
transform 1 0 45448 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_458
timestamp 1586364061
transform 1 0 43240 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_461
timestamp 1586364061
transform 1 0 43516 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_471
timestamp 1586364061
transform 1 0 44436 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_475
timestamp 1586364061
transform 1 0 44804 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_481
timestamp 1586364061
transform 1 0 45356 0 1 15776
box -38 -48 130 592
use scs8hd_inv_8  _611_
timestamp 1586364061
transform 1 0 46092 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 47196 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__611__A
timestamp 1586364061
transform 1 0 45816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_484
timestamp 1586364061
transform 1 0 45632 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_498
timestamp 1586364061
transform 1 0 46920 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_503
timestamp 1586364061
transform 1 0 47380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 48852 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_515
timestamp 1586364061
transform 1 0 48484 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _310_
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_193
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__551__B
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__311__B
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__551__A
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _550_
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__309__A
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__A
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _309_
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__B
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_225
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _306_
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_240
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__306__A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_248
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__615__A
timestamp 1586364061
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__613__A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_inv_8  _615_
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _614_
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_273
timestamp 1586364061
transform 1 0 26220 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_277
timestamp 1586364061
transform 1 0 26588 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_287
timestamp 1586364061
transform 1 0 27508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_294
timestamp 1586364061
transform 1 0 28152 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_290
timestamp 1586364061
transform 1 0 27784 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_291
timestamp 1586364061
transform 1 0 27876 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__547__B
timestamp 1586364061
transform 1 0 28244 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_301
timestamp 1586364061
transform 1 0 28796 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_297
timestamp 1586364061
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_302
timestamp 1586364061
transform 1 0 28888 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_296
timestamp 1586364061
transform 1 0 28336 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__547__A
timestamp 1586364061
transform 1 0 28612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 28980 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_315
timestamp 1586364061
transform 1 0 30084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_314
timestamp 1586364061
transform 1 0 29992 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__305__A
timestamp 1586364061
transform 1 0 30268 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_319
timestamp 1586364061
transform 1 0 30452 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_322
timestamp 1586364061
transform 1 0 30728 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__305__B
timestamp 1586364061
transform 1 0 30636 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_331
timestamp 1586364061
transform 1 0 31556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_327
timestamp 1586364061
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_323
timestamp 1586364061
transform 1 0 30820 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_328
timestamp 1586364061
transform 1 0 31280 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 31464 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 31372 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _336_
timestamp 1586364061
transform 1 0 30912 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _253_
timestamp 1586364061
transform 1 0 31004 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_337
timestamp 1586364061
transform 1 0 32108 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_332
timestamp 1586364061
transform 1 0 31648 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__C
timestamp 1586364061
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__B
timestamp 1586364061
transform 1 0 31740 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use scs8hd_or3_4  _263_
timestamp 1586364061
transform 1 0 31924 0 1 16864
box -38 -48 866 592
use scs8hd_or3_4  _241_
timestamp 1586364061
transform 1 0 32384 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_348
timestamp 1586364061
transform 1 0 33120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_344
timestamp 1586364061
transform 1 0 32752 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__268__B
timestamp 1586364061
transform 1 0 32936 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_355
timestamp 1586364061
transform 1 0 33764 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_357
timestamp 1586364061
transform 1 0 33948 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_349
timestamp 1586364061
transform 1 0 33212 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__313__A
timestamp 1586364061
transform 1 0 33304 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__282__B
timestamp 1586364061
transform 1 0 34040 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _313_
timestamp 1586364061
transform 1 0 33488 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_364
timestamp 1586364061
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_360
timestamp 1586364061
transform 1 0 34224 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_366
timestamp 1586364061
transform 1 0 34776 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_362
timestamp 1586364061
transform 1 0 34408 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 34868 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 34408 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use scs8hd_or3_4  _282_
timestamp 1586364061
transform 1 0 34868 0 1 16864
box -38 -48 866 592
use scs8hd_buf_1  _245_
timestamp 1586364061
transform 1 0 34132 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_369
timestamp 1586364061
transform 1 0 35052 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_8  _240_
timestamp 1586364061
transform 1 0 35144 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_380
timestamp 1586364061
transform 1 0 36064 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_376
timestamp 1586364061
transform 1 0 35696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_386
timestamp 1586364061
transform 1 0 36616 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_383
timestamp 1586364061
transform 1 0 36340 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_379
timestamp 1586364061
transform 1 0 35972 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__282__C
timestamp 1586364061
transform 1 0 35880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 36432 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__286__C
timestamp 1586364061
transform 1 0 36248 0 1 16864
box -38 -48 222 592
use scs8hd_or3_4  _286_
timestamp 1586364061
transform 1 0 36432 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__324__A
timestamp 1586364061
transform 1 0 36800 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__B
timestamp 1586364061
transform 1 0 37168 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_390
timestamp 1586364061
transform 1 0 36984 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_393
timestamp 1586364061
transform 1 0 37260 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__528__A
timestamp 1586364061
transform 1 0 37720 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_394
timestamp 1586364061
transform 1 0 37352 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_398
timestamp 1586364061
transform 1 0 37720 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_397
timestamp 1586364061
transform 1 0 37628 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 37812 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_27_400
timestamp 1586364061
transform 1 0 37904 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_406
timestamp 1586364061
transform 1 0 38456 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_410
timestamp 1586364061
transform 1 0 38824 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__509__B
timestamp 1586364061
transform 1 0 39008 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__509__A
timestamp 1586364061
transform 1 0 38272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__508__A
timestamp 1586364061
transform 1 0 38640 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _509_
timestamp 1586364061
transform 1 0 38824 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_419
timestamp 1586364061
transform 1 0 39652 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_414
timestamp 1586364061
transform 1 0 39192 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__508__B
timestamp 1586364061
transform 1 0 39836 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _512_
timestamp 1586364061
transform 1 0 39560 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_423
timestamp 1586364061
transform 1 0 40020 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_427
timestamp 1586364061
transform 1 0 40388 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40572 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 40388 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 40940 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40940 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_431
timestamp 1586364061
transform 1 0 40756 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_431
timestamp 1586364061
transform 1 0 40756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_435
timestamp 1586364061
transform 1 0 41124 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41676 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_438
timestamp 1586364061
transform 1 0 41400 0 -1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 41676 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_452
timestamp 1586364061
transform 1 0 42688 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_449
timestamp 1586364061
transform 1 0 42412 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_443
timestamp 1586364061
transform 1 0 41860 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42136 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_456
timestamp 1586364061
transform 1 0 43056 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42872 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_466
timestamp 1586364061
transform 1 0 43976 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_462
timestamp 1586364061
transform 1 0 43608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_457
timestamp 1586364061
transform 1 0 43148 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43240 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__606__A
timestamp 1586364061
transform 1 0 43792 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43424 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_473
timestamp 1586364061
transform 1 0 44620 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_469
timestamp 1586364061
transform 1 0 44252 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_470
timestamp 1586364061
transform 1 0 44344 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44160 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44712 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 44620 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_480
timestamp 1586364061
transform 1 0 45264 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_476
timestamp 1586364061
transform 1 0 44896 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_480
timestamp 1586364061
transform 1 0 45264 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_476
timestamp 1586364061
transform 1 0 44896 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45080 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_492
timestamp 1586364061
transform 1 0 46368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_484
timestamp 1586364061
transform 1 0 45632 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_493
timestamp 1586364061
transform 1 0 46460 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 46000 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _610_
timestamp 1586364061
transform 1 0 45632 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_8  FILLER_27_508
timestamp 1586364061
transform 1 0 47840 0 1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_496
timestamp 1586364061
transform 1 0 46736 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_504
timestamp 1586364061
transform 1 0 47472 0 -1 16864
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 47196 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 48852 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 48852 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _551_
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_195
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _549_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_8  _613_
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_245
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_256
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_285
timestamp 1586364061
transform 1 0 27324 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_293
timestamp 1586364061
transform 1 0 28060 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_289
timestamp 1586364061
transform 1 0 27692 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 -1 17952
box -38 -48 314 592
use scs8hd_or2_4  _305_
timestamp 1586364061
transform 1 0 30636 0 -1 17952
box -38 -48 682 592
use scs8hd_or2_4  _547_
timestamp 1586364061
transform 1 0 29164 0 -1 17952
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__553__B
timestamp 1586364061
transform 1 0 30452 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29992 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_297
timestamp 1586364061
transform 1 0 28428 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_312
timestamp 1586364061
transform 1 0 29808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_316
timestamp 1586364061
transform 1 0 30176 0 -1 17952
box -38 -48 314 592
use scs8hd_or2_4  _268_
timestamp 1586364061
transform 1 0 32108 0 -1 17952
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 31832 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__336__A
timestamp 1586364061
transform 1 0 31464 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_328
timestamp 1586364061
transform 1 0 31280 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_332
timestamp 1586364061
transform 1 0 31648 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_344
timestamp 1586364061
transform 1 0 32752 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_8  _237_
timestamp 1586364061
transform 1 0 34408 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__254__B
timestamp 1586364061
transform 1 0 33304 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__498__B
timestamp 1586364061
transform 1 0 33948 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35512 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_352
timestamp 1586364061
transform 1 0 33488 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_356
timestamp 1586364061
transform 1 0 33856 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_359
timestamp 1586364061
transform 1 0 34132 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_371
timestamp 1586364061
transform 1 0 35236 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  _324_
timestamp 1586364061
transform 1 0 35972 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  _528_
timestamp 1586364061
transform 1 0 37720 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__286__B
timestamp 1586364061
transform 1 0 36432 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_376
timestamp 1586364061
transform 1 0 35696 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_382
timestamp 1586364061
transform 1 0 36248 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_386
timestamp 1586364061
transform 1 0 36616 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_394
timestamp 1586364061
transform 1 0 37352 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_401
timestamp 1586364061
transform 1 0 37996 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _508_
timestamp 1586364061
transform 1 0 38916 0 -1 17952
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40572 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39928 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_409
timestamp 1586364061
transform 1 0 38732 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_420
timestamp 1586364061
transform 1 0 39744 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_424
timestamp 1586364061
transform 1 0 40112 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_428
timestamp 1586364061
transform 1 0 40480 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_440
timestamp 1586364061
transform 1 0 41584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_452
timestamp 1586364061
transform 1 0 42688 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44712 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 43240 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 43792 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_462
timestamp 1586364061
transform 1 0 43608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_466
timestamp 1586364061
transform 1 0 43976 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_28_483
timestamp 1586364061
transform 1 0 45540 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 46092 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46460 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_491
timestamp 1586364061
transform 1 0 46276 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_495
timestamp 1586364061
transform 1 0 46644 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_507
timestamp 1586364061
transform 1 0 47748 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 48852 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_515
timestamp 1586364061
transform 1 0 48484 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _577_
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__577__A
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__577__B
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_216
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _548_
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__548__A
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__576__A
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__576__B
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_248
timestamp 1586364061
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_252
timestamp 1586364061
transform 1 0 24288 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__617__A
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25668 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 28244 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_280
timestamp 1586364061
transform 1 0 26864 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_293
timestamp 1586364061
transform 1 0 28060 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_301
timestamp 1586364061
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_297
timestamp 1586364061
transform 1 0 28428 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__554__A
timestamp 1586364061
transform 1 0 28612 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__308__A
timestamp 1586364061
transform 1 0 28980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_309
timestamp 1586364061
transform 1 0 29532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _554_
timestamp 1586364061
transform 1 0 29256 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_317
timestamp 1586364061
transform 1 0 30268 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_313
timestamp 1586364061
transform 1 0 29900 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__308__B
timestamp 1586364061
transform 1 0 29716 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__553__A
timestamp 1586364061
transform 1 0 30360 0 1 17952
box -38 -48 222 592
use scs8hd_or2_4  _252_
timestamp 1586364061
transform 1 0 30544 0 1 17952
box -38 -48 682 592
use scs8hd_or2_4  _274_
timestamp 1586364061
transform 1 0 31924 0 1 17952
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__252__B
timestamp 1586364061
transform 1 0 31372 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 32752 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 31740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__274__B
timestamp 1586364061
transform 1 0 33120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_327
timestamp 1586364061
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_331
timestamp 1586364061
transform 1 0 31556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_342
timestamp 1586364061
transform 1 0 32568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_346
timestamp 1586364061
transform 1 0 32936 0 1 17952
box -38 -48 222 592
use scs8hd_or2_4  _254_
timestamp 1586364061
transform 1 0 33304 0 1 17952
box -38 -48 682 592
use scs8hd_or2_4  _527_
timestamp 1586364061
transform 1 0 34868 0 1 17952
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 34132 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__498__A
timestamp 1586364061
transform 1 0 34500 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_357
timestamp 1586364061
transform 1 0 33948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_361
timestamp 1586364061
transform 1 0 34316 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_365
timestamp 1586364061
transform 1 0 34684 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_374
timestamp 1586364061
transform 1 0 35512 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _497_
timestamp 1586364061
transform 1 0 36340 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__527__A
timestamp 1586364061
transform 1 0 35696 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__497__A
timestamp 1586364061
transform 1 0 36156 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37352 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_378
timestamp 1586364061
transform 1 0 35880 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_392
timestamp 1586364061
transform 1 0 37168 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_396
timestamp 1586364061
transform 1 0 37536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_400
timestamp 1586364061
transform 1 0 37904 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_406
timestamp 1586364061
transform 1 0 38456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__B
timestamp 1586364061
transform 1 0 38272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__A
timestamp 1586364061
transform 1 0 38640 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _507_
timestamp 1586364061
transform 1 0 38824 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_423
timestamp 1586364061
transform 1 0 40020 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_419
timestamp 1586364061
transform 1 0 39652 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 40388 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 40480 0 1 17952
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42504 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42964 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41676 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_439
timestamp 1586364061
transform 1 0 41492 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_443
timestamp 1586364061
transform 1 0 41860 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_449
timestamp 1586364061
transform 1 0 42412 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_453
timestamp 1586364061
transform 1 0 42780 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 43516 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45172 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_457
timestamp 1586364061
transform 1 0 43148 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_472
timestamp 1586364061
transform 1 0 44528 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_477
timestamp 1586364061
transform 1 0 44988 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_481
timestamp 1586364061
transform 1 0 45356 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 46000 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45816 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 47104 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_485
timestamp 1586364061
transform 1 0 45724 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_498
timestamp 1586364061
transform 1 0 46920 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_502
timestamp 1586364061
transform 1 0 47288 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 48852 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_514
timestamp 1586364061
transform 1 0 48392 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__603__B
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_172
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_176
timestamp 1586364061
transform 1 0 17296 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__602__B
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _576_
timestamp 1586364061
transform 1 0 22632 0 -1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_225
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_233
timestamp 1586364061
transform 1 0 22540 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _617_
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_243
timestamp 1586364061
transform 1 0 23460 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_255
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_285
timestamp 1586364061
transform 1 0 27324 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_292
timestamp 1586364061
transform 1 0 27968 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_289
timestamp 1586364061
transform 1 0 27692 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__573__B
timestamp 1586364061
transform 1 0 27784 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_1  _269_
timestamp 1586364061
transform 1 0 28152 0 -1 19040
box -38 -48 314 592
use scs8hd_or2_4  _308_
timestamp 1586364061
transform 1 0 29164 0 -1 19040
box -38 -48 682 592
use scs8hd_or2_4  _553_
timestamp 1586364061
transform 1 0 30544 0 -1 19040
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__599__B
timestamp 1586364061
transform 1 0 28980 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_297
timestamp 1586364061
transform 1 0 28428 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_8  FILLER_30_312
timestamp 1586364061
transform 1 0 29808 0 -1 19040
box -38 -48 774 592
use scs8hd_or2_4  _232_
timestamp 1586364061
transform 1 0 32108 0 -1 19040
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 31372 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_327
timestamp 1586364061
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_331
timestamp 1586364061
transform 1 0 31556 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_335
timestamp 1586364061
transform 1 0 31924 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_344
timestamp 1586364061
transform 1 0 32752 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _498_
timestamp 1586364061
transform 1 0 33948 0 -1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35512 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__527__B
timestamp 1586364061
transform 1 0 34960 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_356
timestamp 1586364061
transform 1 0 33856 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_366
timestamp 1586364061
transform 1 0 34776 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_370
timestamp 1586364061
transform 1 0 35144 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__497__B
timestamp 1586364061
transform 1 0 36524 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37352 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_383
timestamp 1586364061
transform 1 0 36340 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_387
timestamp 1586364061
transform 1 0 36708 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_393
timestamp 1586364061
transform 1 0 37260 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_396
timestamp 1586364061
transform 1 0 37536 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39468 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_409
timestamp 1586364061
transform 1 0 38732 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_420
timestamp 1586364061
transform 1 0 39744 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 40756 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41952 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42872 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_430
timestamp 1586364061
transform 1 0 40664 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_442
timestamp 1586364061
transform 1 0 41768 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_446
timestamp 1586364061
transform 1 0 42136 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_456
timestamp 1586364061
transform 1 0 43056 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43792 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44804 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 43240 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 43516 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_459
timestamp 1586364061
transform 1 0 43332 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_463
timestamp 1586364061
transform 1 0 43700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_467
timestamp 1586364061
transform 1 0 44068 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46368 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_484
timestamp 1586364061
transform 1 0 45632 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_501
timestamp 1586364061
transform 1 0 47196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 48852 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_513
timestamp 1586364061
transform 1 0 48300 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _602_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_nor2_4  _603_
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__603__A
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__602__A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__601__A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__600__A
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_200
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _574_
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__574__A
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__616__A
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_256
timestamp 1586364061
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_260
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_or2_4  _573_
timestamp 1586364061
transform 1 0 27784 0 1 19040
box -38 -48 682 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__573__A
timestamp 1586364061
transform 1 0 27600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_281
timestamp 1586364061
transform 1 0 26956 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_285
timestamp 1586364061
transform 1 0 27324 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _307_
timestamp 1586364061
transform 1 0 29256 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__307__A
timestamp 1586364061
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__599__A
timestamp 1586364061
transform 1 0 28612 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__A
timestamp 1586364061
transform 1 0 30452 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_297
timestamp 1586364061
transform 1 0 28428 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_301
timestamp 1586364061
transform 1 0 28796 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_315
timestamp 1586364061
transform 1 0 30084 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_321
timestamp 1586364061
transform 1 0 30636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_329
timestamp 1586364061
transform 1 0 31372 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_325
timestamp 1586364061
transform 1 0 31004 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__486__B
timestamp 1586364061
transform 1 0 30820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__270__B
timestamp 1586364061
transform 1 0 31464 0 1 19040
box -38 -48 222 592
use scs8hd_or2_4  _270_
timestamp 1586364061
transform 1 0 31648 0 1 19040
box -38 -48 682 592
use scs8hd_fill_2  FILLER_31_343
timestamp 1586364061
transform 1 0 32660 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_339
timestamp 1586364061
transform 1 0 32292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__339__A
timestamp 1586364061
transform 1 0 32844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 32476 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _330_
timestamp 1586364061
transform 1 0 33028 0 1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 34868 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 34408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__330__A
timestamp 1586364061
transform 1 0 33488 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__A
timestamp 1586364061
transform 1 0 33856 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_350
timestamp 1586364061
transform 1 0 33304 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_354
timestamp 1586364061
transform 1 0 33672 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_358
timestamp 1586364061
transform 1 0 34040 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_364
timestamp 1586364061
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37352 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__505__A
timestamp 1586364061
transform 1 0 36064 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37168 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_378
timestamp 1586364061
transform 1 0 35880 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_382
timestamp 1586364061
transform 1 0 36248 0 1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_31_388
timestamp 1586364061
transform 1 0 36800 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_31_407
timestamp 1586364061
transform 1 0 38548 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_403
timestamp 1586364061
transform 1 0 38180 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__506__A
timestamp 1586364061
transform 1 0 38364 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_412
timestamp 1586364061
transform 1 0 39008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__510__B
timestamp 1586364061
transform 1 0 38824 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__510__A
timestamp 1586364061
transform 1 0 39192 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_423
timestamp 1586364061
transform 1 0 40020 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_419
timestamp 1586364061
transform 1 0 39652 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_428
timestamp 1586364061
transform 1 0 40480 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 40388 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41308 0 1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42872 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42320 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41124 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42688 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_434
timestamp 1586364061
transform 1 0 41032 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_446
timestamp 1586364061
transform 1 0 42136 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_450
timestamp 1586364061
transform 1 0 42504 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _641_
timestamp 1586364061
transform 1 0 44988 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43884 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44252 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_463
timestamp 1586364061
transform 1 0 43700 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_467
timestamp 1586364061
transform 1 0 44068 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_471
timestamp 1586364061
transform 1 0 44436 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_480
timestamp 1586364061
transform 1 0 45264 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 46000 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46276 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_484
timestamp 1586364061
transform 1 0 45632 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_489
timestamp 1586364061
transform 1 0 46092 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_493
timestamp 1586364061
transform 1 0 46460 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_505
timestamp 1586364061
transform 1 0 47564 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 48852 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_513
timestamp 1586364061
transform 1 0 48300 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _601_
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__601__B
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_173
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 590 592
use scs8hd_buf_1  _600_
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__575__B
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_207
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_226
timestamp 1586364061
transform 1 0 21896 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_234
timestamp 1586364061
transform 1 0 22632 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_8  _616_
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_248
timestamp 1586364061
transform 1 0 23920 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_256
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__619__A
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__618__A
timestamp 1586364061
transform 1 0 27600 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_273
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_285
timestamp 1586364061
transform 1 0 27324 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_290
timestamp 1586364061
transform 1 0 27784 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _486_
timestamp 1586364061
transform 1 0 30452 0 -1 20128
box -38 -48 866 592
use scs8hd_or2_4  _599_
timestamp 1586364061
transform 1 0 28980 0 -1 20128
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_302
timestamp 1586364061
transform 1 0 28888 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_310
timestamp 1586364061
transform 1 0 29624 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_314
timestamp 1586364061
transform 1 0 29992 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_318
timestamp 1586364061
transform 1 0 30360 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_1  _333_
timestamp 1586364061
transform 1 0 33120 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_1  _339_
timestamp 1586364061
transform 1 0 32108 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_328
timestamp 1586364061
transform 1 0 31280 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_340
timestamp 1586364061
transform 1 0 32384 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _258_
timestamp 1586364061
transform 1 0 34408 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_1  _505_
timestamp 1586364061
transform 1 0 35604 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 34868 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_351
timestamp 1586364061
transform 1 0 33396 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_359
timestamp 1586364061
transform 1 0 34132 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_365
timestamp 1586364061
transform 1 0 34684 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_369
timestamp 1586364061
transform 1 0 35052 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_373
timestamp 1586364061
transform 1 0 35420 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_378
timestamp 1586364061
transform 1 0 35880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_382
timestamp 1586364061
transform 1 0 36248 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_389
timestamp 1586364061
transform 1 0 36892 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_6  FILLER_32_398
timestamp 1586364061
transform 1 0 37720 0 -1 20128
box -38 -48 590 592
use scs8hd_buf_1  _506_
timestamp 1586364061
transform 1 0 38272 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _510_
timestamp 1586364061
transform 1 0 39284 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__513__B
timestamp 1586364061
transform 1 0 39100 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_407
timestamp 1586364061
transform 1 0 38548 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_4  FILLER_32_424
timestamp 1586364061
transform 1 0 40112 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_430
timestamp 1586364061
transform 1 0 40664 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_436
timestamp 1586364061
transform 1 0 41216 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_439
timestamp 1586364061
transform 1 0 41492 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_450
timestamp 1586364061
transform 1 0 42504 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_454
timestamp 1586364061
transform 1 0 42872 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 43240 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_457
timestamp 1586364061
transform 1 0 43148 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_468
timestamp 1586364061
transform 1 0 44160 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_32_479
timestamp 1586364061
transform 1 0 45172 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_483
timestamp 1586364061
transform 1 0 45540 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45908 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45632 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46368 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_486
timestamp 1586364061
transform 1 0 45816 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_490
timestamp 1586364061
transform 1 0 46184 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_494
timestamp 1586364061
transform 1 0 46552 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_506
timestamp 1586364061
transform 1 0 47656 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 48852 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_514
timestamp 1586364061
transform 1 0 48392 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_168
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_175
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_192
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__575__A
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 314 592
use scs8hd_nor2_4  _575_
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_222
timestamp 1586364061
transform 1 0 21528 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 866 592
use scs8hd_conb_1  _638_
timestamp 1586364061
transform 1 0 21252 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_233
timestamp 1586364061
transform 1 0 22540 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_237
timestamp 1586364061
transform 1 0 22908 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_8  FILLER_33_235
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _645_
timestamp 1586364061
transform 1 0 23552 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_248
timestamp 1586364061
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_252
timestamp 1586364061
transform 1 0 24288 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_252
timestamp 1586364061
transform 1 0 24288 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_267
timestamp 1586364061
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 25392 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_8  _619_
timestamp 1586364061
transform 1 0 26036 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_287
timestamp 1586364061
transform 1 0 27508 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_279
timestamp 1586364061
transform 1 0 26772 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_284
timestamp 1586364061
transform 1 0 27232 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_280
timestamp 1586364061
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__488__B
timestamp 1586364061
transform 1 0 27416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__487__A
timestamp 1586364061
transform 1 0 27600 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_8  _618_
timestamp 1586364061
transform 1 0 27600 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_290
timestamp 1586364061
transform 1 0 27784 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _488_
timestamp 1586364061
transform 1 0 27876 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_304
timestamp 1586364061
transform 1 0 29072 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_300
timestamp 1586364061
transform 1 0 28704 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_301
timestamp 1586364061
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_297
timestamp 1586364061
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28888 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__B
timestamp 1586364061
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__488__A
timestamp 1586364061
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_308
timestamp 1586364061
transform 1 0 29440 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_313
timestamp 1586364061
transform 1 0 29900 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29256 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29624 0 -1 21216
box -38 -48 866 592
use scs8hd_or2_4  _579_
timestamp 1586364061
transform 1 0 29256 0 1 20128
box -38 -48 682 592
use scs8hd_decap_6  FILLER_34_319
timestamp 1586364061
transform 1 0 30452 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_321
timestamp 1586364061
transform 1 0 30636 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_317
timestamp 1586364061
transform 1 0 30268 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__A
timestamp 1586364061
transform 1 0 30084 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_333
timestamp 1586364061
transform 1 0 31740 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_327
timestamp 1586364061
transform 1 0 31188 0 -1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31004 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 31004 0 1 20128
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_33_340
timestamp 1586364061
transform 1 0 32384 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_336
timestamp 1586364061
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__B
timestamp 1586364061
transform 1 0 32568 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__A
timestamp 1586364061
transform 1 0 32200 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _485_
timestamp 1586364061
transform 1 0 32108 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_1  _342_
timestamp 1586364061
transform 1 0 32752 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_346
timestamp 1586364061
transform 1 0 32936 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_347
timestamp 1586364061
transform 1 0 33028 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__342__A
timestamp 1586364061
transform 1 0 33212 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__B
timestamp 1586364061
transform 1 0 33212 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__496__B
timestamp 1586364061
transform 1 0 33672 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_351
timestamp 1586364061
transform 1 0 33396 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__496__A
timestamp 1586364061
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_356
timestamp 1586364061
transform 1 0 33856 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_360
timestamp 1586364061
transform 1 0 34224 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_357
timestamp 1586364061
transform 1 0 33948 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _496_
timestamp 1586364061
transform 1 0 34040 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_6  FILLER_34_351
timestamp 1586364061
transform 1 0 33396 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_6  FILLER_34_371
timestamp 1586364061
transform 1 0 35236 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_367
timestamp 1586364061
transform 1 0 34868 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35052 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 34868 0 1 20128
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_33_382
timestamp 1586364061
transform 1 0 36248 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_378
timestamp 1586364061
transform 1 0 35880 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__B
timestamp 1586364061
transform 1 0 36064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__A
timestamp 1586364061
transform 1 0 36432 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35788 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_394
timestamp 1586364061
transform 1 0 37352 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_386
timestamp 1586364061
transform 1 0 36616 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_395
timestamp 1586364061
transform 1 0 37444 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37444 0 -1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _499_
timestamp 1586364061
transform 1 0 36616 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_400
timestamp 1586364061
transform 1 0 37904 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38088 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_412
timestamp 1586364061
transform 1 0 39008 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_407
timestamp 1586364061
transform 1 0 38548 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_404
timestamp 1586364061
transform 1 0 38272 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__511__B
timestamp 1586364061
transform 1 0 38824 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__511__A
timestamp 1586364061
transform 1 0 38640 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _511_
timestamp 1586364061
transform 1 0 38824 0 1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_424
timestamp 1586364061
transform 1 0 40112 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_423
timestamp 1586364061
transform 1 0 40020 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_419
timestamp 1586364061
transform 1 0 39652 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__513__A
timestamp 1586364061
transform 1 0 39836 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _513_
timestamp 1586364061
transform 1 0 39284 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 40388 0 1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 40480 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_34_430
timestamp 1586364061
transform 1 0 40664 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_439
timestamp 1586364061
transform 1 0 41492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41032 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_449
timestamp 1586364061
transform 1 0 42412 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_445
timestamp 1586364061
transform 1 0 42044 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_447
timestamp 1586364061
transform 1 0 42228 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_443
timestamp 1586364061
transform 1 0 41860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42228 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 20128
box -38 -48 866 592
use scs8hd_decap_6  FILLER_34_459
timestamp 1586364061
transform 1 0 43332 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_457
timestamp 1586364061
transform 1 0 43148 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_468
timestamp 1586364061
transform 1 0 44160 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_464
timestamp 1586364061
transform 1 0 43792 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 43976 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 43240 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 43884 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_476
timestamp 1586364061
transform 1 0 44896 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_472
timestamp 1586364061
transform 1 0 44528 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44804 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 44344 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_480
timestamp 1586364061
transform 1 0 45264 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45632 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 46000 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_484
timestamp 1586364061
transform 1 0 45632 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_498
timestamp 1586364061
transform 1 0 46920 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_493
timestamp 1586364061
transform 1 0 46460 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_505
timestamp 1586364061
transform 1 0 47564 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 48852 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 48852 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_510
timestamp 1586364061
transform 1 0 48024 0 1 20128
box -38 -48 590 592
use scs8hd_decap_3  FILLER_34_513
timestamp 1586364061
transform 1 0 48300 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_164
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_conb_1  _637_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_195
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_216
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_224
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_231
timestamp 1586364061
transform 1 0 22356 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_235
timestamp 1586364061
transform 1 0 22724 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_255
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _487_
timestamp 1586364061
transform 1 0 27600 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__487__B
timestamp 1586364061
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_272
timestamp 1586364061
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_278
timestamp 1586364061
transform 1 0 26680 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_284
timestamp 1586364061
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29256 0 1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_297
timestamp 1586364061
transform 1 0 28428 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_301
timestamp 1586364061
transform 1 0 28796 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_317
timestamp 1586364061
transform 1 0 30268 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_321
timestamp 1586364061
transform 1 0 30636 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31556 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__A
timestamp 1586364061
transform 1 0 33028 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31372 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_325
timestamp 1586364061
transform 1 0 31004 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_340
timestamp 1586364061
transform 1 0 32384 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_344
timestamp 1586364061
transform 1 0 32752 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_358
timestamp 1586364061
transform 1 0 34040 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _501_
timestamp 1586364061
transform 1 0 33212 0 1 21216
box -38 -48 866 592
use scs8hd_fill_1  FILLER_35_367
timestamp 1586364061
transform 1 0 34868 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_362
timestamp 1586364061
transform 1 0 34408 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34592 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use scs8hd_conb_1  _642_
timestamp 1586364061
transform 1 0 34960 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_371
timestamp 1586364061
transform 1 0 35236 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35604 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 36616 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 36432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__B
timestamp 1586364061
transform 1 0 37996 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_377
timestamp 1586364061
transform 1 0 35788 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_381
timestamp 1586364061
transform 1 0 36156 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_397
timestamp 1586364061
transform 1 0 37628 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_403
timestamp 1586364061
transform 1 0 38180 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__A
timestamp 1586364061
transform 1 0 38364 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _514_
timestamp 1586364061
transform 1 0 38548 0 1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_35_423
timestamp 1586364061
transform 1 0 40020 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_420
timestamp 1586364061
transform 1 0 39744 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_416
timestamp 1586364061
transform 1 0 39376 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 40388 0 1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 40480 0 1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_439
timestamp 1586364061
transform 1 0 41492 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_443
timestamp 1586364061
transform 1 0 41860 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_456
timestamp 1586364061
transform 1 0 43056 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45448 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44252 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_461
timestamp 1586364061
transform 1 0 43516 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_465
timestamp 1586364061
transform 1 0 43884 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_480
timestamp 1586364061
transform 1 0 45264 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_484
timestamp 1586364061
transform 1 0 45632 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45816 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 46000 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_496
timestamp 1586364061
transform 1 0 46736 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_492
timestamp 1586364061
transform 1 0 46368 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46920 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 47104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_507
timestamp 1586364061
transform 1 0 47748 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_503
timestamp 1586364061
transform 1 0 47380 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47564 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 48852 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_515
timestamp 1586364061
transform 1 0 48484 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_36_157
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_161
timestamp 1586364061
transform 1 0 15916 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_165
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_174
timestamp 1586364061
transform 1 0 17112 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_185
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_189
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_210
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_221
timestamp 1586364061
transform 1 0 21436 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_225
timestamp 1586364061
transform 1 0 21804 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_242
timestamp 1586364061
transform 1 0 23368 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_248
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_259
timestamp 1586364061
transform 1 0 24932 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_265
timestamp 1586364061
transform 1 0 25484 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27508 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27324 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_269
timestamp 1586364061
transform 1 0 25852 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_279
timestamp 1586364061
transform 1 0 26772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_283
timestamp 1586364061
transform 1 0 27140 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_290
timestamp 1586364061
transform 1 0 27784 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28612 0 -1 22304
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_298
timestamp 1586364061
transform 1 0 28520 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_310
timestamp 1586364061
transform 1 0 29624 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_314
timestamp 1586364061
transform 1 0 29992 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_327
timestamp 1586364061
transform 1 0 31188 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  FILLER_36_333
timestamp 1586364061
transform 1 0 31740 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_348
timestamp 1586364061
transform 1 0 33120 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 33856 0 -1 22304
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35604 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35052 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_367
timestamp 1586364061
transform 1 0 34868 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_371
timestamp 1586364061
transform 1 0 35236 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36616 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_384
timestamp 1586364061
transform 1 0 36432 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_388
timestamp 1586364061
transform 1 0 36800 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_393
timestamp 1586364061
transform 1 0 37260 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40204 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_407
timestamp 1586364061
transform 1 0 38548 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_419
timestamp 1586364061
transform 1 0 39652 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_4  FILLER_36_428
timestamp 1586364061
transform 1 0 40480 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__523__B
timestamp 1586364061
transform 1 0 40848 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_434
timestamp 1586364061
transform 1 0 41032 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_445
timestamp 1586364061
transform 1 0 42044 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_453
timestamp 1586364061
transform 1 0 42780 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45172 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 43240 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44436 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_457
timestamp 1586364061
transform 1 0 43148 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_468
timestamp 1586364061
transform 1 0 44160 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_473
timestamp 1586364061
transform 1 0 44620 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46736 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_488
timestamp 1586364061
transform 1 0 46000 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_499
timestamp 1586364061
transform 1 0 47012 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 48852 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_511
timestamp 1586364061
transform 1 0 48116 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_515
timestamp 1586364061
transform 1 0 48484 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_151
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_155
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_214
timestamp 1586364061
transform 1 0 20792 0 1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__415__A
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_222
timestamp 1586364061
transform 1 0 21528 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_255
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_272
timestamp 1586364061
transform 1 0 26128 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_289
timestamp 1586364061
transform 1 0 27692 0 1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28428 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30636 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_299
timestamp 1586364061
transform 1 0 28612 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_315
timestamp 1586364061
transform 1 0 30084 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_319
timestamp 1586364061
transform 1 0 30452 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32108 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31740 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_326
timestamp 1586364061
transform 1 0 31096 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_330
timestamp 1586364061
transform 1 0 31464 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_335
timestamp 1586364061
transform 1 0 31924 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_339
timestamp 1586364061
transform 1 0 32292 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_357
timestamp 1586364061
transform 1 0 33948 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_353
timestamp 1586364061
transform 1 0 33580 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_349
timestamp 1586364061
transform 1 0 33212 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33396 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__A
timestamp 1586364061
transform 1 0 33764 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_361
timestamp 1586364061
transform 1 0 34316 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__B
timestamp 1586364061
transform 1 0 34132 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 22304
box -38 -48 866 592
use scs8hd_fill_1  FILLER_37_384
timestamp 1586364061
transform 1 0 36432 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_380
timestamp 1586364061
transform 1 0 36064 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_376
timestamp 1586364061
transform 1 0 35696 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36524 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_387
timestamp 1586364061
transform 1 0 36708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36892 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37076 0 1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_37_400
timestamp 1586364061
transform 1 0 37904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38088 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_404
timestamp 1586364061
transform 1 0 38272 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_412
timestamp 1586364061
transform 1 0 39008 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__B
timestamp 1586364061
transform 1 0 38824 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__A
timestamp 1586364061
transform 1 0 39192 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_423
timestamp 1586364061
transform 1 0 40020 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_419
timestamp 1586364061
transform 1 0 39652 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_428
timestamp 1586364061
transform 1 0 40480 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 40388 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41308 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41768 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__523__A
timestamp 1586364061
transform 1 0 40848 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_434
timestamp 1586364061
transform 1 0 41032 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_440
timestamp 1586364061
transform 1 0 41584 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_444
timestamp 1586364061
transform 1 0 41952 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_452
timestamp 1586364061
transform 1 0 42688 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44528 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45356 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43976 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_464
timestamp 1586364061
transform 1 0 43792 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_468
timestamp 1586364061
transform 1 0 44160 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_475
timestamp 1586364061
transform 1 0 44804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_479
timestamp 1586364061
transform 1 0 45172 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_483
timestamp 1586364061
transform 1 0 45540 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 46000 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_487
timestamp 1586364061
transform 1 0 45908 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_492
timestamp 1586364061
transform 1 0 46368 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_496
timestamp 1586364061
transform 1 0 46736 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_508
timestamp 1586364061
transform 1 0 47840 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 48852 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_171
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_183
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_198
timestamp 1586364061
transform 1 0 19320 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_204
timestamp 1586364061
transform 1 0 19872 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_208
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 590 592
use scs8hd_buf_1  _415_
timestamp 1586364061
transform 1 0 21344 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_219
timestamp 1586364061
transform 1 0 21252 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_223
timestamp 1586364061
transform 1 0 21620 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_240
timestamp 1586364061
transform 1 0 23184 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_244
timestamp 1586364061
transform 1 0 23552 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_260
timestamp 1586364061
transform 1 0 25024 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_257
timestamp 1586364061
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_268
timestamp 1586364061
transform 1 0 25760 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_264
timestamp 1586364061
transform 1 0 25392 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__490__B
timestamp 1586364061
transform 1 0 27600 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28152 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_285
timestamp 1586364061
transform 1 0 27324 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_290
timestamp 1586364061
transform 1 0 27784 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28428 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29440 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_296
timestamp 1586364061
transform 1 0 28336 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_300
timestamp 1586364061
transform 1 0 28704 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_38_317
timestamp 1586364061
transform 1 0 30268 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _643_
timestamp 1586364061
transform 1 0 31004 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_328
timestamp 1586364061
transform 1 0 31280 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_346
timestamp 1586364061
transform 1 0 32936 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _500_
timestamp 1586364061
transform 1 0 33764 0 -1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35328 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_350
timestamp 1586364061
transform 1 0 33304 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_354
timestamp 1586364061
transform 1 0 33672 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_364
timestamp 1586364061
transform 1 0 34592 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_369
timestamp 1586364061
transform 1 0 35052 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_375
timestamp 1586364061
transform 1 0 35604 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_382
timestamp 1586364061
transform 1 0 36248 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_379
timestamp 1586364061
transform 1 0 35972 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36064 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_392
timestamp 1586364061
transform 1 0 37168 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_388
timestamp 1586364061
transform 1 0 36800 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36984 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_401
timestamp 1586364061
transform 1 0 37996 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_396
timestamp 1586364061
transform 1 0 37536 0 -1 23392
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 23392
box -38 -48 314 592
use scs8hd_nor2_4  _521_
timestamp 1586364061
transform 1 0 39284 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__518__B
timestamp 1586364061
transform 1 0 38824 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40296 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_409
timestamp 1586364061
transform 1 0 38732 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_412
timestamp 1586364061
transform 1 0 39008 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_424
timestamp 1586364061
transform 1 0 40112 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_428
timestamp 1586364061
transform 1 0 40480 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _523_
timestamp 1586364061
transform 1 0 40848 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40664 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_441
timestamp 1586364061
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_453
timestamp 1586364061
transform 1 0 42780 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44528 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 43240 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 44252 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_457
timestamp 1586364061
transform 1 0 43148 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_462
timestamp 1586364061
transform 1 0 43608 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_468
timestamp 1586364061
transform 1 0 44160 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_471
timestamp 1586364061
transform 1 0 44436 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_475
timestamp 1586364061
transform 1 0 44804 0 -1 23392
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46000 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_487
timestamp 1586364061
transform 1 0 45908 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_490
timestamp 1586364061
transform 1 0 46184 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_502
timestamp 1586364061
transform 1 0 47288 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 48852 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_514
timestamp 1586364061
transform 1 0 48392 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_171
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_192
timestamp 1586364061
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_205
timestamp 1586364061
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_198
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_209
timestamp 1586364061
transform 1 0 20332 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_223
timestamp 1586364061
transform 1 0 21620 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_233
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_237
timestamp 1586364061
transform 1 0 22908 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_6  FILLER_40_250
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_248
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_256
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_252
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_267
timestamp 1586364061
transform 1 0 25668 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_277
timestamp 1586364061
transform 1 0 26588 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_273
timestamp 1586364061
transform 1 0 26220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25944 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_289
timestamp 1586364061
transform 1 0 27692 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_285
timestamp 1586364061
transform 1 0 27324 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_285
timestamp 1586364061
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_281
timestamp 1586364061
transform 1 0 26956 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__490__A
timestamp 1586364061
transform 1 0 27416 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _490_
timestamp 1586364061
transform 1 0 27600 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_293
timestamp 1586364061
transform 1 0 28060 0 -1 24480
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 28152 0 -1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_40_305
timestamp 1586364061
transform 1 0 29164 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_301
timestamp 1586364061
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_297
timestamp 1586364061
transform 1 0 28428 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_313
timestamp 1586364061
transform 1 0 29900 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_309
timestamp 1586364061
transform 1 0 29532 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29348 0 -1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_321
timestamp 1586364061
transform 1 0 30636 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_317
timestamp 1586364061
transform 1 0 30268 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_319
timestamp 1586364061
transform 1 0 30452 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_315
timestamp 1586364061
transform 1 0 30084 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30452 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30268 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_328
timestamp 1586364061
transform 1 0 31280 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_330
timestamp 1586364061
transform 1 0 31464 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_326
timestamp 1586364061
transform 1 0 31096 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_333
timestamp 1586364061
transform 1 0 31740 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_339
timestamp 1586364061
transform 1 0 32292 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_334
timestamp 1586364061
transform 1 0 31832 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32476 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31648 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_346
timestamp 1586364061
transform 1 0 32936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_347
timestamp 1586364061
transform 1 0 33028 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_343
timestamp 1586364061
transform 1 0 32660 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32752 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_358
timestamp 1586364061
transform 1 0 34040 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_350
timestamp 1586364061
transform 1 0 33304 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_358
timestamp 1586364061
transform 1 0 34040 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_351
timestamp 1586364061
transform 1 0 33396 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34132 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33212 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_372
timestamp 1586364061
transform 1 0 35328 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_363
timestamp 1586364061
transform 1 0 34500 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 34316 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 23392
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 34316 0 -1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35512 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_376
timestamp 1586364061
transform 1 0 35696 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_382
timestamp 1586364061
transform 1 0 36248 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_376
timestamp 1586364061
transform 1 0 35696 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_393
timestamp 1586364061
transform 1 0 37260 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_389
timestamp 1586364061
transform 1 0 36892 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36800 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_398
timestamp 1586364061
transform 1 0 37720 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_402
timestamp 1586364061
transform 1 0 38088 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_397
timestamp 1586364061
transform 1 0 37628 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__519__A
timestamp 1586364061
transform 1 0 37904 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _519_
timestamp 1586364061
transform 1 0 37904 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_409
timestamp 1586364061
transform 1 0 38732 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_406
timestamp 1586364061
transform 1 0 38456 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__519__B
timestamp 1586364061
transform 1 0 38272 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__518__A
timestamp 1586364061
transform 1 0 38640 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _518_
timestamp 1586364061
transform 1 0 38824 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_423
timestamp 1586364061
transform 1 0 40020 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_419
timestamp 1586364061
transform 1 0 39652 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 39468 0 -1 24480
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_40_428
timestamp 1586364061
transform 1 0 40480 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_428
timestamp 1586364061
transform 1 0 40480 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 40388 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_433
timestamp 1586364061
transform 1 0 40940 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_441
timestamp 1586364061
transform 1 0 41676 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 -1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40664 0 1 23392
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 41216 0 -1 24480
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_40_451
timestamp 1586364061
transform 1 0 42596 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_447
timestamp 1586364061
transform 1 0 42228 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_453
timestamp 1586364061
transform 1 0 42780 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_449
timestamp 1586364061
transform 1 0 42412 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_445
timestamp 1586364061
transform 1 0 42044 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42412 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42228 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 41860 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_467
timestamp 1586364061
transform 1 0 44068 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_459
timestamp 1586364061
transform 1 0 43332 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_457
timestamp 1586364061
transform 1 0 43148 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_466
timestamp 1586364061
transform 1 0 43976 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 43240 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43148 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_477
timestamp 1586364061
transform 1 0 44988 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_471
timestamp 1586364061
transform 1 0 44436 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 44252 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45172 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44712 0 1 23392
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 44252 0 -1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_40_480
timestamp 1586364061
transform 1 0 45264 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_481
timestamp 1586364061
transform 1 0 45356 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45448 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_484
timestamp 1586364061
transform 1 0 45632 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_492
timestamp 1586364061
transform 1 0 46368 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_485
timestamp 1586364061
transform 1 0 45724 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 46000 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46000 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_497
timestamp 1586364061
transform 1 0 46828 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_508
timestamp 1586364061
transform 1 0 47840 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_39_496
timestamp 1586364061
transform 1 0 46736 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_509
timestamp 1586364061
transform 1 0 47932 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 48852 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 48852 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_515
timestamp 1586364061
transform 1 0 48484 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_154
timestamp 1586364061
transform 1 0 15272 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_158
timestamp 1586364061
transform 1 0 15640 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_200
timestamp 1586364061
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_213
timestamp 1586364061
transform 1 0 20700 0 1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_217
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_224
timestamp 1586364061
transform 1 0 21712 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_254
timestamp 1586364061
transform 1 0 24472 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26864 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28060 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_274
timestamp 1586364061
transform 1 0 26312 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_278
timestamp 1586364061
transform 1 0 26680 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_291
timestamp 1586364061
transform 1 0 27876 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_295
timestamp 1586364061
transform 1 0 28244 0 1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29808 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28704 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_299
timestamp 1586364061
transform 1 0 28612 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_302
timestamp 1586364061
transform 1 0 28888 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_306
timestamp 1586364061
transform 1 0 29256 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_310
timestamp 1586364061
transform 1 0 29624 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_327
timestamp 1586364061
transform 1 0 31188 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_323
timestamp 1586364061
transform 1 0 30820 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31372 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31556 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_340
timestamp 1586364061
transform 1 0 32384 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_344
timestamp 1586364061
transform 1 0 32752 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32568 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32936 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33120 0 1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34132 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_357
timestamp 1586364061
transform 1 0 33948 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_361
timestamp 1586364061
transform 1 0 34316 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_385
timestamp 1586364061
transform 1 0 36524 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_380
timestamp 1586364061
transform 1 0 36064 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_376
timestamp 1586364061
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36340 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36708 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_400
timestamp 1586364061
transform 1 0 37904 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_396
timestamp 1586364061
transform 1 0 37536 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38088 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38272 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 40388 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__520__A
timestamp 1586364061
transform 1 0 39284 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__520__B
timestamp 1586364061
transform 1 0 39652 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_413
timestamp 1586364061
transform 1 0 39100 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_417
timestamp 1586364061
transform 1 0 39468 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_421
timestamp 1586364061
transform 1 0 39836 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_41_428
timestamp 1586364061
transform 1 0 40480 0 1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 42320 0 1 24480
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40756 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 42136 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_440
timestamp 1586364061
transform 1 0 41584 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_444
timestamp 1586364061
transform 1 0 41952 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44252 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45448 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43884 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_459
timestamp 1586364061
transform 1 0 43332 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_463
timestamp 1586364061
transform 1 0 43700 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_467
timestamp 1586364061
transform 1 0 44068 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_480
timestamp 1586364061
transform 1 0 45264 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 46000 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45816 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_484
timestamp 1586364061
transform 1 0 45632 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_498
timestamp 1586364061
transform 1 0 46920 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 48852 0 1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_41_510
timestamp 1586364061
transform 1 0 48024 0 1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_151
timestamp 1586364061
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_169
timestamp 1586364061
transform 1 0 16652 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_182
timestamp 1586364061
transform 1 0 17848 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_186
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_189
timestamp 1586364061
transform 1 0 18492 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_207
timestamp 1586364061
transform 1 0 20148 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_215
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_221
timestamp 1586364061
transform 1 0 21436 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_225
timestamp 1586364061
transform 1 0 21804 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_229
timestamp 1586364061
transform 1 0 22172 0 -1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__465__B
timestamp 1586364061
transform 1 0 24656 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_247
timestamp 1586364061
transform 1 0 23828 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_255
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_267
timestamp 1586364061
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_271
timestamp 1586364061
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_287
timestamp 1586364061
transform 1 0 27508 0 -1 25568
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28704 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29716 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_299
timestamp 1586364061
transform 1 0 28612 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_309
timestamp 1586364061
transform 1 0 29532 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_313
timestamp 1586364061
transform 1 0 29900 0 -1 25568
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_328
timestamp 1586364061
transform 1 0 31280 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_346
timestamp 1586364061
transform 1 0 32936 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34776 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34224 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_354
timestamp 1586364061
transform 1 0 33672 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_358
timestamp 1586364061
transform 1 0 34040 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_362
timestamp 1586364061
transform 1 0 34408 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_375
timestamp 1586364061
transform 1 0 35604 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_381
timestamp 1586364061
transform 1 0 36156 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35972 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_386
timestamp 1586364061
transform 1 0 36616 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36800 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36340 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_396
timestamp 1586364061
transform 1 0 37536 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_390
timestamp 1586364061
transform 1 0 36984 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_401
timestamp 1586364061
transform 1 0 37996 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 25568
box -38 -48 314 592
use scs8hd_nor2_4  _520_
timestamp 1586364061
transform 1 0 39192 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__525__A
timestamp 1586364061
transform 1 0 38180 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38548 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_405
timestamp 1586364061
transform 1 0 38364 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_409
timestamp 1586364061
transform 1 0 38732 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_413
timestamp 1586364061
transform 1 0 39100 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_423
timestamp 1586364061
transform 1 0 40020 0 -1 25568
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40940 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41400 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_431
timestamp 1586364061
transform 1 0 40756 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_435
timestamp 1586364061
transform 1 0 41124 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_449
timestamp 1586364061
transform 1 0 42412 0 -1 25568
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45172 0 -1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 43240 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44436 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_457
timestamp 1586364061
transform 1 0 43148 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_468
timestamp 1586364061
transform 1 0 44160 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_473
timestamp 1586364061
transform 1 0 44620 0 -1 25568
box -38 -48 590 592
use scs8hd_conb_1  _640_
timestamp 1586364061
transform 1 0 46736 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 46184 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_488
timestamp 1586364061
transform 1 0 46000 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_492
timestamp 1586364061
transform 1 0 46368 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_499
timestamp 1586364061
transform 1 0 47012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 48852 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_511
timestamp 1586364061
transform 1 0 48116 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_515
timestamp 1586364061
transform 1 0 48484 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 14812 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_43_160
timestamp 1586364061
transform 1 0 15824 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_168
timestamp 1586364061
transform 1 0 16560 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_164
timestamp 1586364061
transform 1 0 16192 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 25568
box -38 -48 222 592
use scs8hd_conb_1  _646_
timestamp 1586364061
transform 1 0 16928 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_179
timestamp 1586364061
transform 1 0 17572 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_175
timestamp 1586364061
transform 1 0 17204 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 25568
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_195
timestamp 1586364061
transform 1 0 19044 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_199
timestamp 1586364061
transform 1 0 19412 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_214
timestamp 1586364061
transform 1 0 20792 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 22540 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22908 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_218
timestamp 1586364061
transform 1 0 21160 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_231
timestamp 1586364061
transform 1 0 22356 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_235
timestamp 1586364061
transform 1 0 22724 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_239
timestamp 1586364061
transform 1 0 23092 0 1 25568
box -38 -48 406 592
use scs8hd_decap_4  FILLER_43_252
timestamp 1586364061
transform 1 0 24288 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_248
timestamp 1586364061
transform 1 0 23920 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_243
timestamp 1586364061
transform 1 0 23460 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_43_263
timestamp 1586364061
transform 1 0 25300 0 1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_43_259
timestamp 1586364061
transform 1 0 24932 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_256
timestamp 1586364061
transform 1 0 24656 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__465__A
timestamp 1586364061
transform 1 0 24748 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 25392 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 25576 0 1 25568
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26956 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_277
timestamp 1586364061
transform 1 0 26588 0 1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_43_283
timestamp 1586364061
transform 1 0 27140 0 1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_43_291
timestamp 1586364061
transform 1 0 27876 0 1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30268 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_297
timestamp 1586364061
transform 1 0 28428 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_301
timestamp 1586364061
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_315
timestamp 1586364061
transform 1 0 30084 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_319
timestamp 1586364061
transform 1 0 30452 0 1 25568
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_330
timestamp 1586364061
transform 1 0 31464 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31188 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_334
timestamp 1586364061
transform 1 0 31832 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__495__A
timestamp 1586364061
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31648 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_341
timestamp 1586364061
transform 1 0 32476 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_345
timestamp 1586364061
transform 1 0 32844 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_351
timestamp 1586364061
transform 1 0 33396 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__494__A
timestamp 1586364061
transform 1 0 33212 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_358
timestamp 1586364061
transform 1 0 34040 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_362
timestamp 1586364061
transform 1 0 34408 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_370
timestamp 1586364061
transform 1 0 35144 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_374
timestamp 1586364061
transform 1 0 35512 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_381
timestamp 1586364061
transform 1 0 36156 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_378
timestamp 1586364061
transform 1 0 35880 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_386
timestamp 1586364061
transform 1 0 36616 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36800 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36340 0 1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_43_390
timestamp 1586364061
transform 1 0 36984 0 1 25568
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__525__B
timestamp 1586364061
transform 1 0 37536 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_402
timestamp 1586364061
transform 1 0 38088 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_398
timestamp 1586364061
transform 1 0 37720 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 25568
box -38 -48 222 592
use scs8hd_nor2_4  _525_
timestamp 1586364061
transform 1 0 38180 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 40388 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__522__A
timestamp 1586364061
transform 1 0 39192 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__B
timestamp 1586364061
transform 1 0 39560 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_412
timestamp 1586364061
transform 1 0 39008 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_416
timestamp 1586364061
transform 1 0 39376 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_420
timestamp 1586364061
transform 1 0 39744 0 1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_43_426
timestamp 1586364061
transform 1 0 40296 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_428
timestamp 1586364061
transform 1 0 40480 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_432
timestamp 1586364061
transform 1 0 40848 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40664 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 1 25568
box -38 -48 866 592
use scs8hd_decap_3  FILLER_43_446
timestamp 1586364061
transform 1 0 42136 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_442
timestamp 1586364061
transform 1 0 41768 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41952 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_455
timestamp 1586364061
transform 1 0 42964 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_451
timestamp 1586364061
transform 1 0 42596 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43148 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_472
timestamp 1586364061
transform 1 0 44528 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_468
timestamp 1586364061
transform 1 0 44160 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44712 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_483
timestamp 1586364061
transform 1 0 45540 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_479
timestamp 1586364061
transform 1 0 45172 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45356 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_43_487
timestamp 1586364061
transform 1 0 45908 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45724 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_492
timestamp 1586364061
transform 1 0 46368 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 46000 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_496
timestamp 1586364061
transform 1 0 46736 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 47104 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_507
timestamp 1586364061
transform 1 0 47748 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_503
timestamp 1586364061
transform 1 0 47380 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47564 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 47932 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 48852 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_511
timestamp 1586364061
transform 1 0 48116 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_515
timestamp 1586364061
transform 1 0 48484 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__453__A
timestamp 1586364061
transform 1 0 14260 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__B
timestamp 1586364061
transform 1 0 14996 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_6  FILLER_44_169
timestamp 1586364061
transform 1 0 16652 0 -1 26656
box -38 -48 590 592
use scs8hd_fill_2  FILLER_44_165
timestamp 1586364061
transform 1 0 16284 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__455__B
timestamp 1586364061
transform 1 0 16468 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_179
timestamp 1586364061
transform 1 0 17572 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_175
timestamp 1586364061
transform 1 0 17204 0 -1 26656
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_186
timestamp 1586364061
transform 1 0 18216 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_183
timestamp 1586364061
transform 1 0 17940 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19320 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_196
timestamp 1586364061
transform 1 0 19136 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_200
timestamp 1586364061
transform 1 0 19504 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_205
timestamp 1586364061
transform 1 0 19964 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_213
timestamp 1586364061
transform 1 0 20700 0 -1 26656
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 26656
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__468__B
timestamp 1586364061
transform 1 0 21344 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_218
timestamp 1586364061
transform 1 0 21160 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_222
timestamp 1586364061
transform 1 0 21528 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_227
timestamp 1586364061
transform 1 0 21988 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _465_
timestamp 1586364061
transform 1 0 24748 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__464__B
timestamp 1586364061
transform 1 0 25760 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_242
timestamp 1586364061
transform 1 0 23368 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_44_254
timestamp 1586364061
transform 1 0 24472 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_266
timestamp 1586364061
transform 1 0 25576 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_270
timestamp 1586364061
transform 1 0 25944 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_276
timestamp 1586364061
transform 1 0 26496 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_274
timestamp 1586364061
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__466__B
timestamp 1586364061
transform 1 0 26680 0 -1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_280
timestamp 1586364061
transform 1 0 26864 0 -1 26656
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26956 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_284
timestamp 1586364061
transform 1 0 27232 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_290
timestamp 1586364061
transform 1 0 27784 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__489__B
timestamp 1586364061
transform 1 0 27600 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27968 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_295
timestamp 1586364061
transform 1 0 28244 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_299
timestamp 1586364061
transform 1 0 28612 0 -1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28428 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28980 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_306
timestamp 1586364061
transform 1 0 29256 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_310
timestamp 1586364061
transform 1 0 29624 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_317
timestamp 1586364061
transform 1 0 30268 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30452 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_321
timestamp 1586364061
transform 1 0 30636 0 -1 26656
box -38 -48 222 592
use scs8hd_buf_1  _495_
timestamp 1586364061
transform 1 0 32200 0 -1 26656
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_328
timestamp 1586364061
transform 1 0 31280 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_337
timestamp 1586364061
transform 1 0 32108 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_341
timestamp 1586364061
transform 1 0 32476 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_345
timestamp 1586364061
transform 1 0 32844 0 -1 26656
box -38 -48 406 592
use scs8hd_buf_1  _494_
timestamp 1586364061
transform 1 0 33212 0 -1 26656
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 34224 0 -1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__502__B
timestamp 1586364061
transform 1 0 33856 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35604 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_352
timestamp 1586364061
transform 1 0 33488 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_358
timestamp 1586364061
transform 1 0 34040 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_371
timestamp 1586364061
transform 1 0 35236 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37904 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_377
timestamp 1586364061
transform 1 0 35788 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_388
timestamp 1586364061
transform 1 0 36800 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_396
timestamp 1586364061
transform 1 0 37536 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_398
timestamp 1586364061
transform 1 0 37720 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _522_
timestamp 1586364061
transform 1 0 38916 0 -1 26656
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38364 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_403
timestamp 1586364061
transform 1 0 38180 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_407
timestamp 1586364061
transform 1 0 38548 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_8  FILLER_44_420
timestamp 1586364061
transform 1 0 39744 0 -1 26656
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40940 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_431
timestamp 1586364061
transform 1 0 40756 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_435
timestamp 1586364061
transform 1 0 41124 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_8  FILLER_44_450
timestamp 1586364061
transform 1 0 42504 0 -1 26656
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 43240 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 44528 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_468
timestamp 1586364061
transform 1 0 44160 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_8  FILLER_44_474
timestamp 1586364061
transform 1 0 44712 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_482
timestamp 1586364061
transform 1 0 45448 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 47196 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45632 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46644 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_493
timestamp 1586364061
transform 1 0 46460 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_497
timestamp 1586364061
transform 1 0 46828 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_504
timestamp 1586364061
transform 1 0 47472 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 48852 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_45_139
timestamp 1586364061
transform 1 0 13892 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__453__B
timestamp 1586364061
transform 1 0 13708 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__413__A
timestamp 1586364061
transform 1 0 14076 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _453_
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_152
timestamp 1586364061
transform 1 0 15088 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_156
timestamp 1586364061
transform 1 0 15456 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__455__A
timestamp 1586364061
transform 1 0 15640 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__A
timestamp 1586364061
transform 1 0 15272 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _455_
timestamp 1586364061
transform 1 0 15824 0 1 26656
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18032 0 1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__452__A
timestamp 1586364061
transform 1 0 17020 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__452__B
timestamp 1586364061
transform 1 0 17388 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_169
timestamp 1586364061
transform 1 0 16652 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_175
timestamp 1586364061
transform 1 0 17204 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_179
timestamp 1586364061
transform 1 0 17572 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19780 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_195
timestamp 1586364061
transform 1 0 19044 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_199
timestamp 1586364061
transform 1 0 19412 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_214
timestamp 1586364061
transform 1 0 20792 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21804 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__468__A
timestamp 1586364061
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_218
timestamp 1586364061
transform 1 0 21160 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_222
timestamp 1586364061
transform 1 0 21528 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_236
timestamp 1586364061
transform 1 0 22816 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_240
timestamp 1586364061
transform 1 0 23184 0 1 26656
box -38 -48 222 592
use scs8hd_buf_1  _419_
timestamp 1586364061
transform 1 0 24012 0 1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _464_
timestamp 1586364061
transform 1 0 25024 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__419__A
timestamp 1586364061
transform 1 0 24472 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__463__A
timestamp 1586364061
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_245
timestamp 1586364061
transform 1 0 23644 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_252
timestamp 1586364061
transform 1 0 24288 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_256
timestamp 1586364061
transform 1 0 24656 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_273
timestamp 1586364061
transform 1 0 26220 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_269
timestamp 1586364061
transform 1 0 25852 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__466__A
timestamp 1586364061
transform 1 0 26404 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__464__A
timestamp 1586364061
transform 1 0 26036 0 1 26656
box -38 -48 222 592
use scs8hd_buf_1  _417_
timestamp 1586364061
transform 1 0 26588 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_284
timestamp 1586364061
transform 1 0 27232 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_280
timestamp 1586364061
transform 1 0 26864 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__489__A
timestamp 1586364061
transform 1 0 27416 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__417__A
timestamp 1586364061
transform 1 0 27048 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _489_
timestamp 1586364061
transform 1 0 27600 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_301
timestamp 1586364061
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_297
timestamp 1586364061
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_319
timestamp 1586364061
transform 1 0 30452 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_315
timestamp 1586364061
transform 1 0 30084 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30636 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__503__A
timestamp 1586364061
transform 1 0 33028 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__503__B
timestamp 1586364061
transform 1 0 32660 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_332
timestamp 1586364061
transform 1 0 31648 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_336
timestamp 1586364061
transform 1 0 32016 0 1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_45_339
timestamp 1586364061
transform 1 0 32292 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_345
timestamp 1586364061
transform 1 0 32844 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _503_
timestamp 1586364061
transform 1 0 33212 0 1 26656
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 34868 0 1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__502__A
timestamp 1586364061
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_358
timestamp 1586364061
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_362
timestamp 1586364061
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36616 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__517__A
timestamp 1586364061
transform 1 0 37996 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37628 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_378
timestamp 1586364061
transform 1 0 35880 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_382
timestamp 1586364061
transform 1 0 36248 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_395
timestamp 1586364061
transform 1 0 37444 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_399
timestamp 1586364061
transform 1 0 37812 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_412
timestamp 1586364061
transform 1 0 39008 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 39192 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38180 0 1 26656
box -38 -48 866 592
use scs8hd_fill_1  FILLER_45_424
timestamp 1586364061
transform 1 0 40112 0 1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_45_420
timestamp 1586364061
transform 1 0 39744 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_416
timestamp 1586364061
transform 1 0 39376 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39560 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 40388 0 1 26656
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 40480 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_439
timestamp 1586364061
transform 1 0 41492 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_443
timestamp 1586364061
transform 1 0 41860 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_447
timestamp 1586364061
transform 1 0 42228 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_453
timestamp 1586364061
transform 1 0 42780 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43148 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 44528 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45448 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44160 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_466
timestamp 1586364061
transform 1 0 43976 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_470
timestamp 1586364061
transform 1 0 44344 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_474
timestamp 1586364061
transform 1 0 44712 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_480
timestamp 1586364061
transform 1 0 45264 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 46000 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 47104 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 47472 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_484
timestamp 1586364061
transform 1 0 45632 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_498
timestamp 1586364061
transform 1 0 46920 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_502
timestamp 1586364061
transform 1 0 47288 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_506
timestamp 1586364061
transform 1 0 47656 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 48852 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_514
timestamp 1586364061
transform 1 0 48392 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__456__B
timestamp 1586364061
transform 1 0 13248 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 774 592
use scs8hd_fill_1  FILLER_47_131
timestamp 1586364061
transform 1 0 13156 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_134
timestamp 1586364061
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_138
timestamp 1586364061
transform 1 0 13800 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__456__A
timestamp 1586364061
transform 1 0 13616 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__407__A
timestamp 1586364061
transform 1 0 13984 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _456_
timestamp 1586364061
transform 1 0 14168 0 1 27744
box -38 -48 866 592
use scs8hd_buf_1  _413_
timestamp 1586364061
transform 1 0 14168 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_47_151
timestamp 1586364061
transform 1 0 14996 0 1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_161
timestamp 1586364061
transform 1 0 15916 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_157
timestamp 1586364061
transform 1 0 15548 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _454_
timestamp 1586364061
transform 1 0 15272 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_46_168
timestamp 1586364061
transform 1 0 16560 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_3  FILLER_46_163
timestamp 1586364061
transform 1 0 16100 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__457__B
timestamp 1586364061
transform 1 0 16376 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__457__A
timestamp 1586364061
transform 1 0 16192 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _457_
timestamp 1586364061
transform 1 0 16376 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_179
timestamp 1586364061
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_175
timestamp 1586364061
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_172
timestamp 1586364061
transform 1 0 16928 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__441__A
timestamp 1586364061
transform 1 0 17388 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _452_
timestamp 1586364061
transform 1 0 17020 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_187
timestamp 1586364061
transform 1 0 18308 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_186
timestamp 1586364061
transform 1 0 18216 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_182
timestamp 1586364061
transform 1 0 17848 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__441__B
timestamp 1586364061
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use scs8hd_buf_1  _451_
timestamp 1586364061
transform 1 0 18032 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_47_199
timestamp 1586364061
transform 1 0 19412 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_195
timestamp 1586364061
transform 1 0 19044 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_191
timestamp 1586364061
transform 1 0 18676 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_194
timestamp 1586364061
transform 1 0 18952 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__451__A
timestamp 1586364061
transform 1 0 18492 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__459__B
timestamp 1586364061
transform 1 0 19228 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__459__A
timestamp 1586364061
transform 1 0 18860 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 27744
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_46_206
timestamp 1586364061
transform 1 0 20056 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__458__A
timestamp 1586364061
transform 1 0 19688 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _458_
timestamp 1586364061
transform 1 0 19872 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_213
timestamp 1586364061
transform 1 0 20700 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_6  FILLER_47_217
timestamp 1586364061
transform 1 0 21068 0 1 27744
box -38 -48 590 592
use scs8hd_decap_4  FILLER_46_225
timestamp 1586364061
transform 1 0 21804 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_215
timestamp 1586364061
transform 1 0 20884 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__450__A
timestamp 1586364061
transform 1 0 20884 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__467__A
timestamp 1586364061
transform 1 0 21620 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _468_
timestamp 1586364061
transform 1 0 20976 0 -1 27744
box -38 -48 866 592
use scs8hd_nor2_4  _467_
timestamp 1586364061
transform 1 0 21804 0 1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_47_238
timestamp 1586364061
transform 1 0 23000 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_234
timestamp 1586364061
transform 1 0 22632 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_232
timestamp 1586364061
transform 1 0 22448 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_229
timestamp 1586364061
transform 1 0 22172 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__469__B
timestamp 1586364061
transform 1 0 22264 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__469__A
timestamp 1586364061
transform 1 0 22816 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22540 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_47_245
timestamp 1586364061
transform 1 0 23644 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_248
timestamp 1586364061
transform 1 0 23920 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_244
timestamp 1586364061
transform 1 0 23552 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__B
timestamp 1586364061
transform 1 0 23736 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__A
timestamp 1586364061
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use scs8hd_nor2_4  _470_
timestamp 1586364061
transform 1 0 23736 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_263
timestamp 1586364061
transform 1 0 25300 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_259
timestamp 1586364061
transform 1 0 24932 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_255
timestamp 1586364061
transform 1 0 24564 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25116 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__463__B
timestamp 1586364061
transform 1 0 24656 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24748 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 25484 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _463_
timestamp 1586364061
transform 1 0 24840 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_46_267
timestamp 1586364061
transform 1 0 25668 0 -1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 25668 0 1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_278
timestamp 1586364061
transform 1 0 26680 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_271
timestamp 1586364061
transform 1 0 26036 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26864 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use scs8hd_nor2_4  _466_
timestamp 1586364061
transform 1 0 26496 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_290
timestamp 1586364061
transform 1 0 27784 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_47_282
timestamp 1586364061
transform 1 0 27048 0 1 27744
box -38 -48 774 592
use scs8hd_decap_8  FILLER_46_285
timestamp 1586364061
transform 1 0 27324 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__475__B
timestamp 1586364061
transform 1 0 27968 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_293
timestamp 1586364061
transform 1 0 28060 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 27744
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 28152 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_301
timestamp 1586364061
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_297
timestamp 1586364061
transform 1 0 28428 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_305
timestamp 1586364061
transform 1 0 29164 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__475__A
timestamp 1586364061
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_313
timestamp 1586364061
transform 1 0 29900 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_309
timestamp 1586364061
transform 1 0 29532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_309
timestamp 1586364061
transform 1 0 29532 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29348 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_322
timestamp 1586364061
transform 1 0 30728 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_317
timestamp 1586364061
transform 1 0 30268 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_317
timestamp 1586364061
transform 1 0 30268 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__472__A
timestamp 1586364061
transform 1 0 30084 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 27744
box -38 -48 866 592
use scs8hd_buf_1  _484_
timestamp 1586364061
transform 1 0 30452 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_326
timestamp 1586364061
transform 1 0 31096 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_332
timestamp 1586364061
transform 1 0 31648 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_327
timestamp 1586364061
transform 1 0 31188 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31464 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__461__A
timestamp 1586364061
transform 1 0 30912 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 31280 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 31464 0 1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_345
timestamp 1586364061
transform 1 0 32844 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_341
timestamp 1586364061
transform 1 0 32476 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__B
timestamp 1586364061
transform 1 0 31832 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__A
timestamp 1586364061
transform 1 0 32660 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_46_348
timestamp 1586364061
transform 1 0 33120 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__A
timestamp 1586364061
transform 1 0 33028 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_356
timestamp 1586364061
transform 1 0 33856 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_352
timestamp 1586364061
transform 1 0 33488 0 1 27744
box -38 -48 406 592
use scs8hd_decap_4  FILLER_46_352
timestamp 1586364061
transform 1 0 33488 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__483__A
timestamp 1586364061
transform 1 0 33304 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__A
timestamp 1586364061
transform 1 0 33948 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _502_
timestamp 1586364061
transform 1 0 33856 0 -1 27744
box -38 -48 866 592
use scs8hd_buf_1  _483_
timestamp 1586364061
transform 1 0 33212 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_367
timestamp 1586364061
transform 1 0 34868 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_363
timestamp 1586364061
transform 1 0 34500 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_359
timestamp 1586364061
transform 1 0 34132 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_365
timestamp 1586364061
transform 1 0 34684 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__D
timestamp 1586364061
transform 1 0 34868 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__B
timestamp 1586364061
transform 1 0 34316 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_374
timestamp 1586364061
transform 1 0 35512 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_373
timestamp 1586364061
transform 1 0 35420 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_369
timestamp 1586364061
transform 1 0 35052 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__C
timestamp 1586364061
transform 1 0 35052 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35604 0 -1 27744
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35236 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_378
timestamp 1586364061
transform 1 0 35880 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_384
timestamp 1586364061
transform 1 0 36432 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__515__A
timestamp 1586364061
transform 1 0 36064 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35696 0 1 27744
box -38 -48 222 592
use scs8hd_buf_1  _328_
timestamp 1586364061
transform 1 0 36248 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_389
timestamp 1586364061
transform 1 0 36892 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_385
timestamp 1586364061
transform 1 0 36524 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_388
timestamp 1586364061
transform 1 0 36800 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__331__A
timestamp 1586364061
transform 1 0 37076 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__328__A
timestamp 1586364061
transform 1 0 36708 0 1 27744
box -38 -48 222 592
use scs8hd_buf_1  _337_
timestamp 1586364061
transform 1 0 37260 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_400
timestamp 1586364061
transform 1 0 37904 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_396
timestamp 1586364061
transform 1 0 37536 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_402
timestamp 1586364061
transform 1 0 38088 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_398
timestamp 1586364061
transform 1 0 37720 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_396
timestamp 1586364061
transform 1 0 37536 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__337__A
timestamp 1586364061
transform 1 0 38088 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__A
timestamp 1586364061
transform 1 0 37720 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_414
timestamp 1586364061
transform 1 0 39192 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_404
timestamp 1586364061
transform 1 0 38272 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_410
timestamp 1586364061
transform 1 0 38824 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_406
timestamp 1586364061
transform 1 0 38456 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__524__B
timestamp 1586364061
transform 1 0 38640 0 -1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 39192 0 -1 27744
box -38 -48 1050 592
use scs8hd_nor2_4  _524_
timestamp 1586364061
transform 1 0 38364 0 1 27744
box -38 -48 866 592
use scs8hd_buf_1  _517_
timestamp 1586364061
transform 1 0 38180 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_426
timestamp 1586364061
transform 1 0 40296 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_422
timestamp 1586364061
transform 1 0 39928 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_418
timestamp 1586364061
transform 1 0 39560 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_425
timestamp 1586364061
transform 1 0 40204 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__364__B
timestamp 1586364061
transform 1 0 39744 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__364__A
timestamp 1586364061
transform 1 0 39376 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_428
timestamp 1586364061
transform 1 0 40480 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 40388 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_432
timestamp 1586364061
transform 1 0 40848 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_436
timestamp 1586364061
transform 1 0 41216 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_4  FILLER_46_430
timestamp 1586364061
transform 1 0 40664 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40664 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41032 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_447
timestamp 1586364061
transform 1 0 42228 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_443
timestamp 1586364061
transform 1 0 41860 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_440
timestamp 1586364061
transform 1 0 41584 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_454
timestamp 1586364061
transform 1 0 42872 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_450
timestamp 1586364061
transform 1 0 42504 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43056 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42596 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_466
timestamp 1586364061
transform 1 0 43976 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_462
timestamp 1586364061
transform 1 0 43608 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_458
timestamp 1586364061
transform 1 0 43240 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_462
timestamp 1586364061
transform 1 0 43608 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43424 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44068 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_47_474
timestamp 1586364061
transform 1 0 44712 0 1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_470
timestamp 1586364061
transform 1 0 44344 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_470
timestamp 1586364061
transform 1 0 44344 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44528 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 44528 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_47_482
timestamp 1586364061
transform 1 0 45448 0 1 27744
box -38 -48 130 592
use scs8hd_decap_6  FILLER_46_483
timestamp 1586364061
transform 1 0 45540 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45540 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46276 0 -1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 46000 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__425__A
timestamp 1586364061
transform 1 0 47104 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 46092 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_500
timestamp 1586364061
transform 1 0 47104 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_47_485
timestamp 1586364061
transform 1 0 45724 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_498
timestamp 1586364061
transform 1 0 46920 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_502
timestamp 1586364061
transform 1 0 47288 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 48852 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 48852 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_512
timestamp 1586364061
transform 1 0 48208 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_514
timestamp 1586364061
transform 1 0 48392 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__442__B
timestamp 1586364061
transform 1 0 13248 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_134
timestamp 1586364061
transform 1 0 13432 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_138
timestamp 1586364061
transform 1 0 13800 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__443__B
timestamp 1586364061
transform 1 0 13616 0 -1 28832
box -38 -48 222 592
use scs8hd_buf_1  _407_
timestamp 1586364061
transform 1 0 14168 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_151
timestamp 1586364061
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_48_158
timestamp 1586364061
transform 1 0 15640 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_154
timestamp 1586364061
transform 1 0 15272 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 28832
box -38 -48 866 592
use scs8hd_nor2_4  _441_
timestamp 1586364061
transform 1 0 17296 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_168
timestamp 1586364061
transform 1 0 16560 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_185
timestamp 1586364061
transform 1 0 18124 0 -1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _459_
timestamp 1586364061
transform 1 0 18860 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__458__B
timestamp 1586364061
transform 1 0 19872 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_189
timestamp 1586364061
transform 1 0 18492 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_202
timestamp 1586364061
transform 1 0 19688 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_206
timestamp 1586364061
transform 1 0 20056 0 -1 28832
box -38 -48 774 592
use scs8hd_buf_1  _450_
timestamp 1586364061
transform 1 0 20884 0 -1 28832
box -38 -48 314 592
use scs8hd_nor2_4  _469_
timestamp 1586364061
transform 1 0 22264 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__467__B
timestamp 1586364061
transform 1 0 21804 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_218
timestamp 1586364061
transform 1 0 21160 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_222
timestamp 1586364061
transform 1 0 21528 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_227
timestamp 1586364061
transform 1 0 21988 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_239
timestamp 1586364061
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24472 0 -1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__477__B
timestamp 1586364061
transform 1 0 25760 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_251
timestamp 1586364061
transform 1 0 24196 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_265
timestamp 1586364061
transform 1 0 25484 0 -1 28832
box -38 -48 314 592
use scs8hd_nor2_4  _475_
timestamp 1586364061
transform 1 0 28152 0 -1 28832
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_270
timestamp 1586364061
transform 1 0 25944 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_274
timestamp 1586364061
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_279
timestamp 1586364061
transform 1 0 26772 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_48_291
timestamp 1586364061
transform 1 0 27876 0 -1 28832
box -38 -48 314 592
use scs8hd_buf_1  _472_
timestamp 1586364061
transform 1 0 29992 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__484__A
timestamp 1586364061
transform 1 0 30452 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29256 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29624 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_303
timestamp 1586364061
transform 1 0 28980 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_308
timestamp 1586364061
transform 1 0 29440 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_312
timestamp 1586364061
transform 1 0 29808 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_317
timestamp 1586364061
transform 1 0 30268 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_321
timestamp 1586364061
transform 1 0 30636 0 -1 28832
box -38 -48 406 592
use scs8hd_buf_1  _461_
timestamp 1586364061
transform 1 0 31004 0 -1 28832
box -38 -48 314 592
use scs8hd_nor2_4  _492_
timestamp 1586364061
transform 1 0 32108 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__491__B
timestamp 1586364061
transform 1 0 31464 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_328
timestamp 1586364061
transform 1 0 31280 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_332
timestamp 1586364061
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_3  FILLER_48_346
timestamp 1586364061
transform 1 0 32936 0 -1 28832
box -38 -48 314 592
use scs8hd_or4_4  _526_
timestamp 1586364061
transform 1 0 34316 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 33212 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__C
timestamp 1586364061
transform 1 0 33580 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__A
timestamp 1586364061
transform 1 0 35328 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__B
timestamp 1586364061
transform 1 0 34132 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_351
timestamp 1586364061
transform 1 0 33396 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_355
timestamp 1586364061
transform 1 0 33764 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_48_370
timestamp 1586364061
transform 1 0 35144 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_374
timestamp 1586364061
transform 1 0 35512 0 -1 28832
box -38 -48 406 592
use scs8hd_buf_1  _331_
timestamp 1586364061
transform 1 0 36432 0 -1 28832
box -38 -48 314 592
use scs8hd_buf_1  _334_
timestamp 1586364061
transform 1 0 37720 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__515__D
timestamp 1586364061
transform 1 0 35972 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_378
timestamp 1586364061
transform 1 0 35880 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  FILLER_48_381
timestamp 1586364061
transform 1 0 36156 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_387
timestamp 1586364061
transform 1 0 36708 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_395
timestamp 1586364061
transform 1 0 37444 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_401
timestamp 1586364061
transform 1 0 37996 0 -1 28832
box -38 -48 406 592
use scs8hd_nor2_4  _364_
timestamp 1586364061
transform 1 0 39008 0 -1 28832
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__524__A
timestamp 1586364061
transform 1 0 38364 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38732 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_407
timestamp 1586364061
transform 1 0 38548 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_411
timestamp 1586364061
transform 1 0 38916 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_421
timestamp 1586364061
transform 1 0 39836 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41400 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41032 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_432
timestamp 1586364061
transform 1 0 40848 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_436
timestamp 1586364061
transform 1 0 41216 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_449
timestamp 1586364061
transform 1 0 42412 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_453
timestamp 1586364061
transform 1 0 42780 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_462
timestamp 1586364061
transform 1 0 43608 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_457
timestamp 1586364061
transform 1 0 43148 0 -1 28832
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 43240 0 -1 28832
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_470
timestamp 1586364061
transform 1 0 44344 0 -1 28832
box -38 -48 222 592
use scs8hd_conb_1  _653_
timestamp 1586364061
transform 1 0 44528 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_479
timestamp 1586364061
transform 1 0 45172 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_475
timestamp 1586364061
transform 1 0 44804 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45356 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44988 0 -1 28832
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45540 0 -1 28832
box -38 -48 314 592
use scs8hd_buf_1  _425_
timestamp 1586364061
transform 1 0 46552 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__318__A
timestamp 1586364061
transform 1 0 47012 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46092 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_486
timestamp 1586364061
transform 1 0 45816 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_491
timestamp 1586364061
transform 1 0 46276 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_497
timestamp 1586364061
transform 1 0 46828 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_501
timestamp 1586364061
transform 1 0 47196 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 48852 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_513
timestamp 1586364061
transform 1 0 48300 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_nor2_4  _442_
timestamp 1586364061
transform 1 0 13248 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__442__A
timestamp 1586364061
transform 1 0 13064 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_129
timestamp 1586364061
transform 1 0 12972 0 1 28832
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14812 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__443__A
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_141
timestamp 1586364061
transform 1 0 14076 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_145
timestamp 1586364061
transform 1 0 14444 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_160
timestamp 1586364061
transform 1 0 15824 0 1 28832
box -38 -48 222 592
use scs8hd_buf_1  _421_
timestamp 1586364061
transform 1 0 16928 0 1 28832
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18032 0 1 28832
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__421__A
timestamp 1586364061
transform 1 0 17388 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_164
timestamp 1586364061
transform 1 0 16192 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_175
timestamp 1586364061
transform 1 0 17204 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_179
timestamp 1586364061
transform 1 0 17572 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_195
timestamp 1586364061
transform 1 0 19044 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_199
timestamp 1586364061
transform 1 0 19412 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_205
timestamp 1586364061
transform 1 0 19964 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_209
timestamp 1586364061
transform 1 0 20332 0 1 28832
box -38 -48 222 592
use scs8hd_buf_1  _462_
timestamp 1586364061
transform 1 0 22540 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__478__A
timestamp 1586364061
transform 1 0 23000 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__B
timestamp 1586364061
transform 1 0 22356 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_222
timestamp 1586364061
transform 1 0 21528 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_226
timestamp 1586364061
transform 1 0 21896 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_230
timestamp 1586364061
transform 1 0 22264 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_236
timestamp 1586364061
transform 1 0 22816 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_240
timestamp 1586364061
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_250
timestamp 1586364061
transform 1 0 24104 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_245
timestamp 1586364061
transform 1 0 23644 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__462__A
timestamp 1586364061
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_258
timestamp 1586364061
transform 1 0 24840 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_254
timestamp 1586364061
transform 1 0 24472 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_262
timestamp 1586364061
transform 1 0 25208 0 1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__477__A
timestamp 1586364061
transform 1 0 25576 0 1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _477_
timestamp 1586364061
transform 1 0 25760 0 1 28832
box -38 -48 866 592
use scs8hd_buf_1  _473_
timestamp 1586364061
transform 1 0 28152 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27968 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27140 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_277
timestamp 1586364061
transform 1 0 26588 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_281
timestamp 1586364061
transform 1 0 26956 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_285
timestamp 1586364061
transform 1 0 27324 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_291
timestamp 1586364061
transform 1 0 27876 0 1 28832
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__A
timestamp 1586364061
transform 1 0 30636 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__473__A
timestamp 1586364061
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_297
timestamp 1586364061
transform 1 0 28428 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_301
timestamp 1586364061
transform 1 0 28796 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_315
timestamp 1586364061
transform 1 0 30084 0 1 28832
box -38 -48 590 592
use scs8hd_nor2_4  _491_
timestamp 1586364061
transform 1 0 31188 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 33028 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__C
timestamp 1586364061
transform 1 0 32660 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__D
timestamp 1586364061
transform 1 0 32292 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__491__A
timestamp 1586364061
transform 1 0 31004 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_323
timestamp 1586364061
transform 1 0 30820 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_336
timestamp 1586364061
transform 1 0 32016 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_341
timestamp 1586364061
transform 1 0 32476 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_345
timestamp 1586364061
transform 1 0 32844 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_358
timestamp 1586364061
transform 1 0 34040 0 1 28832
box -38 -48 222 592
use scs8hd_or4_4  _231_
timestamp 1586364061
transform 1 0 33212 0 1 28832
box -38 -48 866 592
use scs8hd_fill_1  FILLER_49_367
timestamp 1586364061
transform 1 0 34868 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_362
timestamp 1586364061
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__314__A
timestamp 1586364061
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__C
timestamp 1586364061
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use scs8hd_buf_1  _314_
timestamp 1586364061
transform 1 0 34960 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_375
timestamp 1586364061
transform 1 0 35604 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_371
timestamp 1586364061
transform 1 0 35236 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__D
timestamp 1586364061
transform 1 0 35420 0 1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _362_
timestamp 1586364061
transform 1 0 37628 0 1 28832
box -38 -48 866 592
use scs8hd_or4_4  _515_
timestamp 1586364061
transform 1 0 35972 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__515__C
timestamp 1586364061
transform 1 0 35788 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__325__A
timestamp 1586364061
transform 1 0 36984 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__362__A
timestamp 1586364061
transform 1 0 37444 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_388
timestamp 1586364061
transform 1 0 36800 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_392
timestamp 1586364061
transform 1 0 37168 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_410
timestamp 1586364061
transform 1 0 38824 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_406
timestamp 1586364061
transform 1 0 38456 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__516__A
timestamp 1586364061
transform 1 0 39008 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38640 0 1 28832
box -38 -48 222 592
use scs8hd_buf_1  _516_
timestamp 1586364061
transform 1 0 39192 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_423
timestamp 1586364061
transform 1 0 40020 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_417
timestamp 1586364061
transform 1 0 39468 0 1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__423__A
timestamp 1586364061
transform 1 0 39836 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 40388 0 1 28832
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40480 0 1 28832
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 41676 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_439
timestamp 1586364061
transform 1 0 41492 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_443
timestamp 1586364061
transform 1 0 41860 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_456
timestamp 1586364061
transform 1 0 43056 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 43332 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44252 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45448 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 43700 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_461
timestamp 1586364061
transform 1 0 43516 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_465
timestamp 1586364061
transform 1 0 43884 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_480
timestamp 1586364061
transform 1 0 45264 0 1 28832
box -38 -48 222 592
use scs8hd_inv_8  _229_
timestamp 1586364061
transform 1 0 46736 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 46000 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__318__B
timestamp 1586364061
transform 1 0 46552 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 45816 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_484
timestamp 1586364061
transform 1 0 45632 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_489
timestamp 1586364061
transform 1 0 46092 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_493
timestamp 1586364061
transform 1 0 46460 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_505
timestamp 1586364061
transform 1 0 47564 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 48852 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_513
timestamp 1586364061
transform 1 0 48300 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _443_
timestamp 1586364061
transform 1 0 13616 0 -1 29920
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_50_135
timestamp 1586364061
transform 1 0 13524 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_6  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 590 592
use scs8hd_conb_1  _647_
timestamp 1586364061
transform 1 0 17204 0 -1 29920
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_165
timestamp 1586364061
transform 1 0 16284 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_173
timestamp 1586364061
transform 1 0 17020 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_178
timestamp 1586364061
transform 1 0 17480 0 -1 29920
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_195
timestamp 1586364061
transform 1 0 19044 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_206
timestamp 1586364061
transform 1 0 20056 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_210
timestamp 1586364061
transform 1 0 20424 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _478_
timestamp 1586364061
transform 1 0 22632 0 -1 29920
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_8  FILLER_50_224
timestamp 1586364061
transform 1 0 21712 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_232
timestamp 1586364061
transform 1 0 22448 0 -1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 23644 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24012 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_243
timestamp 1586364061
transform 1 0 23460 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_247
timestamp 1586364061
transform 1 0 23828 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_260
timestamp 1586364061
transform 1 0 25024 0 -1 29920
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_50_272
timestamp 1586364061
transform 1 0 26128 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_50_276
timestamp 1586364061
transform 1 0 26496 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_287
timestamp 1586364061
transform 1 0 27508 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_295
timestamp 1586364061
transform 1 0 28244 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 28428 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__460__A
timestamp 1586364061
transform 1 0 30452 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29624 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29992 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_308
timestamp 1586364061
transform 1 0 29440 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_312
timestamp 1586364061
transform 1 0 29808 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_316
timestamp 1586364061
transform 1 0 30176 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_321
timestamp 1586364061
transform 1 0 30636 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_328
timestamp 1586364061
transform 1 0 31280 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__C
timestamp 1586364061
transform 1 0 30820 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__D
timestamp 1586364061
transform 1 0 31464 0 -1 29920
box -38 -48 222 592
use scs8hd_buf_1  _340_
timestamp 1586364061
transform 1 0 31004 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_341
timestamp 1586364061
transform 1 0 32476 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_337
timestamp 1586364061
transform 1 0 32108 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_332
timestamp 1586364061
transform 1 0 31648 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__A
timestamp 1586364061
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__D
timestamp 1586364061
transform 1 0 32292 0 -1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__482__D
timestamp 1586364061
transform 1 0 32844 0 -1 29920
box -38 -48 222 592
use scs8hd_or4_4  _482_
timestamp 1586364061
transform 1 0 33028 0 -1 29920
box -38 -48 866 592
use scs8hd_or4_4  _493_
timestamp 1586364061
transform 1 0 34592 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__578__D
timestamp 1586364061
transform 1 0 34408 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__482__B
timestamp 1586364061
transform 1 0 34040 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_356
timestamp 1586364061
transform 1 0 33856 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_360
timestamp 1586364061
transform 1 0 34224 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_373
timestamp 1586364061
transform 1 0 35420 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_378
timestamp 1586364061
transform 1 0 35880 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__515__B
timestamp 1586364061
transform 1 0 35696 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_382
timestamp 1586364061
transform 1 0 36248 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 36064 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__C
timestamp 1586364061
transform 1 0 36432 0 -1 29920
box -38 -48 222 592
use scs8hd_buf_1  _325_
timestamp 1586364061
transform 1 0 36616 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_389
timestamp 1586364061
transform 1 0 36892 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__A
timestamp 1586364061
transform 1 0 37076 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_393
timestamp 1586364061
transform 1 0 37260 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_398
timestamp 1586364061
transform 1 0 37720 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__382__A
timestamp 1586364061
transform 1 0 37444 0 -1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_50_402
timestamp 1586364061
transform 1 0 38088 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__362__B
timestamp 1586364061
transform 1 0 37904 0 -1 29920
box -38 -48 222 592
use scs8hd_buf_1  _423_
timestamp 1586364061
transform 1 0 40112 0 -1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 38364 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__363__B
timestamp 1586364061
transform 1 0 39560 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40572 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_416
timestamp 1586364061
transform 1 0 39376 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_420
timestamp 1586364061
transform 1 0 39744 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_50_427
timestamp 1586364061
transform 1 0 40388 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 41492 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_431
timestamp 1586364061
transform 1 0 40756 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_450
timestamp 1586364061
transform 1 0 42504 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_454
timestamp 1586364061
transform 1 0 42872 0 -1 29920
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 43332 0 -1 29920
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45080 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 43240 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44528 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44896 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_470
timestamp 1586364061
transform 1 0 44344 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_474
timestamp 1586364061
transform 1 0 44712 0 -1 29920
box -38 -48 222 592
use scs8hd_nand2_4  _318_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 46736 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_8  FILLER_50_487
timestamp 1586364061
transform 1 0 45908 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_50_495
timestamp 1586364061
transform 1 0 46644 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_505
timestamp 1586364061
transform 1 0 47564 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 48852 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_513
timestamp 1586364061
transform 1 0 48300 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__444__A
timestamp 1586364061
transform 1 0 13340 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__444__B
timestamp 1586364061
transform 1 0 12972 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_127
timestamp 1586364061
transform 1 0 12788 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_131
timestamp 1586364061
transform 1 0 13156 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_142
timestamp 1586364061
transform 1 0 14168 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_138
timestamp 1586364061
transform 1 0 13800 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_51_153
timestamp 1586364061
transform 1 0 15180 0 1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_51_149
timestamp 1586364061
transform 1 0 14812 0 1 29920
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_51_156
timestamp 1586364061
transform 1 0 15456 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_51_170
timestamp 1586364061
transform 1 0 16744 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_166
timestamp 1586364061
transform 1 0 16376 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_179
timestamp 1586364061
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_174
timestamp 1586364061
transform 1 0 17112 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 29920
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 29920
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_193
timestamp 1586364061
transform 1 0 18860 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_197
timestamp 1586364061
transform 1 0 19228 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_204
timestamp 1586364061
transform 1 0 19872 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_208
timestamp 1586364061
transform 1 0 20240 0 1 29920
box -38 -48 222 592
use scs8hd_buf_1  _439_
timestamp 1586364061
transform 1 0 22172 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__439__A
timestamp 1586364061
transform 1 0 22632 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_221
timestamp 1586364061
transform 1 0 21436 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_225
timestamp 1586364061
transform 1 0 21804 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_232
timestamp 1586364061
transform 1 0 22448 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_236
timestamp 1586364061
transform 1 0 22816 0 1 29920
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 23644 0 1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_242
timestamp 1586364061
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_256
timestamp 1586364061
transform 1 0 24656 0 1 29920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_51_261
timestamp 1586364061
transform 1 0 25116 0 1 29920
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 26220 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27968 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 26036 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27416 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_269
timestamp 1586364061
transform 1 0 25852 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_284
timestamp 1586364061
transform 1 0 27232 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_288
timestamp 1586364061
transform 1 0 27600 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_295
timestamp 1586364061
transform 1 0 28244 0 1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 29256 0 1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__C
timestamp 1586364061
transform 1 0 30544 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_299
timestamp 1586364061
transform 1 0 28612 0 1 29920
box -38 -48 406 592
use scs8hd_decap_3  FILLER_51_317
timestamp 1586364061
transform 1 0 30268 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_322
timestamp 1586364061
transform 1 0 30728 0 1 29920
box -38 -48 222 592
use scs8hd_or4_4  _460_
timestamp 1586364061
transform 1 0 31464 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__552__B
timestamp 1586364061
transform 1 0 33028 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__B
timestamp 1586364061
transform 1 0 31280 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__B
timestamp 1586364061
transform 1 0 32476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__343__A
timestamp 1586364061
transform 1 0 30912 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_326
timestamp 1586364061
transform 1 0 31096 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_339
timestamp 1586364061
transform 1 0 32292 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_343
timestamp 1586364061
transform 1 0 32660 0 1 29920
box -38 -48 406 592
use scs8hd_decap_4  FILLER_51_358
timestamp 1586364061
transform 1 0 34040 0 1 29920
box -38 -48 406 592
use scs8hd_or4_4  _552_
timestamp 1586364061
transform 1 0 33212 0 1 29920
box -38 -48 866 592
use scs8hd_fill_1  FILLER_51_365
timestamp 1586364061
transform 1 0 34684 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_362
timestamp 1586364061
transform 1 0 34408 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__578__A
timestamp 1586364061
transform 1 0 34500 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use scs8hd_buf_1  _319_
timestamp 1586364061
transform 1 0 34868 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_374
timestamp 1586364061
transform 1 0 35512 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_370
timestamp 1586364061
transform 1 0 35144 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__B
timestamp 1586364061
transform 1 0 35328 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_378
timestamp 1586364061
transform 1 0 35880 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__578__C
timestamp 1586364061
transform 1 0 35696 0 1 29920
box -38 -48 222 592
use scs8hd_or4_4  _504_
timestamp 1586364061
transform 1 0 35972 0 1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_51_392
timestamp 1586364061
transform 1 0 37168 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_388
timestamp 1586364061
transform 1 0 36800 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__B
timestamp 1586364061
transform 1 0 37352 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__D
timestamp 1586364061
transform 1 0 36984 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_399
timestamp 1586364061
transform 1 0 37812 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__360__A
timestamp 1586364061
transform 1 0 37996 0 1 29920
box -38 -48 222 592
use scs8hd_buf_1  _382_
timestamp 1586364061
transform 1 0 37536 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_403
timestamp 1586364061
transform 1 0 38180 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__A
timestamp 1586364061
transform 1 0 38364 0 1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _361_
timestamp 1586364061
transform 1 0 38548 0 1 29920
box -38 -48 866 592
use scs8hd_fill_1  FILLER_51_424
timestamp 1586364061
transform 1 0 40112 0 1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_51_420
timestamp 1586364061
transform 1 0 39744 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_416
timestamp 1586364061
transform 1 0 39376 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__363__A
timestamp 1586364061
transform 1 0 39560 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 40388 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 40480 0 1 29920
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42688 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42504 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_439
timestamp 1586364061
transform 1 0 41492 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_443
timestamp 1586364061
transform 1 0 41860 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_447
timestamp 1586364061
transform 1 0 42228 0 1 29920
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44252 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45448 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_461
timestamp 1586364061
transform 1 0 43516 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_465
timestamp 1586364061
transform 1 0 43884 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_480
timestamp 1586364061
transform 1 0 45264 0 1 29920
box -38 -48 222 592
use scs8hd_or2_4  _230_
timestamp 1586364061
transform 1 0 46644 0 1 29920
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 46000 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 47472 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46276 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_484
timestamp 1586364061
transform 1 0 45632 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_489
timestamp 1586364061
transform 1 0 46092 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_493
timestamp 1586364061
transform 1 0 46460 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_502
timestamp 1586364061
transform 1 0 47288 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_506
timestamp 1586364061
transform 1 0 47656 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 48852 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_514
timestamp 1586364061
transform 1 0 48392 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_8  FILLER_52_128
timestamp 1586364061
transform 1 0 12880 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_131
timestamp 1586364061
transform 1 0 13156 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_142
timestamp 1586364061
transform 1 0 14168 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_138
timestamp 1586364061
transform 1 0 13800 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 31008
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _444_
timestamp 1586364061
transform 1 0 13616 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_153
timestamp 1586364061
transform 1 0 15180 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_149
timestamp 1586364061
transform 1 0 14812 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 31008
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 31008
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_53_173
timestamp 1586364061
transform 1 0 17020 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_170
timestamp 1586364061
transform 1 0 16744 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_166
timestamp 1586364061
transform 1 0 16376 0 1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_165
timestamp 1586364061
transform 1 0 16284 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_179
timestamp 1586364061
transform 1 0 17572 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_177
timestamp 1586364061
transform 1 0 17388 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 31008
box -38 -48 866 592
use scs8hd_decap_3  FILLER_53_197
timestamp 1586364061
transform 1 0 19228 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_193
timestamp 1586364061
transform 1 0 18860 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_191
timestamp 1586364061
transform 1 0 18676 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_206
timestamp 1586364061
transform 1 0 20056 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_202
timestamp 1586364061
transform 1 0 19688 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_52_211
timestamp 1586364061
transform 1 0 20516 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_206
timestamp 1586364061
transform 1 0 20056 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_226
timestamp 1586364061
transform 1 0 21896 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_222
timestamp 1586364061
transform 1 0 21528 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_218
timestamp 1586364061
transform 1 0 21160 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_224
timestamp 1586364061
transform 1 0 21712 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_240
timestamp 1586364061
transform 1 0 23184 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_236
timestamp 1586364061
transform 1 0 22816 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_230
timestamp 1586364061
transform 1 0 22264 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_236
timestamp 1586364061
transform 1 0 22816 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23000 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__476__B
timestamp 1586364061
transform 1 0 22356 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 31008
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 31008
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_53_250
timestamp 1586364061
transform 1 0 24104 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_245
timestamp 1586364061
transform 1 0 23644 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_251
timestamp 1586364061
transform 1 0 24196 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__476__A
timestamp 1586364061
transform 1 0 23368 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_52_256
timestamp 1586364061
transform 1 0 24656 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_53_267
timestamp 1586364061
transform 1 0 25668 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_263
timestamp 1586364061
transform 1 0 25300 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_262
timestamp 1586364061
transform 1 0 25208 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_53_281
timestamp 1586364061
transform 1 0 26956 0 1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_52_274
timestamp 1586364061
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_270
timestamp 1586364061
transform 1 0 25944 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26128 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_292
timestamp 1586364061
transform 1 0 27968 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_285
timestamp 1586364061
transform 1 0 27324 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_301
timestamp 1586364061
transform 1 0 28796 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_296
timestamp 1586364061
transform 1 0 28336 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_52_297
timestamp 1586364061
transform 1 0 28428 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28796 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__480__A
timestamp 1586364061
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__474__A
timestamp 1586364061
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28980 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_312
timestamp 1586364061
transform 1 0 29808 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__480__B
timestamp 1586364061
transform 1 0 29992 0 -1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _474_
timestamp 1586364061
transform 1 0 29256 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_320
timestamp 1586364061
transform 1 0 30544 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_315
timestamp 1586364061
transform 1 0 30084 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_322
timestamp 1586364061
transform 1 0 30728 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_6  FILLER_52_316
timestamp 1586364061
transform 1 0 30176 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__438__C
timestamp 1586364061
transform 1 0 30360 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_328
timestamp 1586364061
transform 1 0 31280 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_324
timestamp 1586364061
transform 1 0 30912 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_52_328
timestamp 1586364061
transform 1 0 31280 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__471__A
timestamp 1586364061
transform 1 0 30820 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__D
timestamp 1586364061
transform 1 0 31556 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__B
timestamp 1586364061
transform 1 0 31372 0 1 31008
box -38 -48 222 592
use scs8hd_or4_4  _438_
timestamp 1586364061
transform 1 0 31556 0 1 31008
box -38 -48 866 592
use scs8hd_buf_1  _343_
timestamp 1586364061
transform 1 0 31004 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_340
timestamp 1586364061
transform 1 0 32384 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_333
timestamp 1586364061
transform 1 0 31740 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use scs8hd_or4_4  _449_
timestamp 1586364061
transform 1 0 32108 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_3  FILLER_53_344
timestamp 1586364061
transform 1 0 32752 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_346
timestamp 1586364061
transform 1 0 32936 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__381__A
timestamp 1586364061
transform 1 0 33028 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__B
timestamp 1586364061
transform 1 0 32568 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_358
timestamp 1586364061
transform 1 0 34040 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_355
timestamp 1586364061
transform 1 0 33764 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_351
timestamp 1586364061
transform 1 0 33396 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__A
timestamp 1586364061
transform 1 0 33948 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__D
timestamp 1586364061
transform 1 0 33580 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__C
timestamp 1586364061
transform 1 0 33212 0 -1 31008
box -38 -48 222 592
use scs8hd_inv_8  _381_
timestamp 1586364061
transform 1 0 33212 0 1 31008
box -38 -48 866 592
use scs8hd_fill_1  FILLER_53_365
timestamp 1586364061
transform 1 0 34684 0 1 31008
box -38 -48 130 592
use scs8hd_fill_1  FILLER_53_362
timestamp 1586364061
transform 1 0 34408 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_359
timestamp 1586364061
transform 1 0 34132 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__316__A
timestamp 1586364061
transform 1 0 34500 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use scs8hd_or4_4  _578_
timestamp 1586364061
transform 1 0 34500 0 -1 31008
box -38 -48 866 592
use scs8hd_buf_1  _345_
timestamp 1586364061
transform 1 0 34868 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_374
timestamp 1586364061
transform 1 0 35512 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_370
timestamp 1586364061
transform 1 0 35144 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_372
timestamp 1586364061
transform 1 0 35328 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__319__A
timestamp 1586364061
transform 1 0 35512 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__345__A
timestamp 1586364061
transform 1 0 35328 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_384
timestamp 1586364061
transform 1 0 36432 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_378
timestamp 1586364061
transform 1 0 35880 0 1 31008
box -38 -48 406 592
use scs8hd_decap_4  FILLER_52_383
timestamp 1586364061
transform 1 0 36340 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_376
timestamp 1586364061
transform 1 0 35696 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__B
timestamp 1586364061
transform 1 0 35880 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__A
timestamp 1586364061
transform 1 0 35696 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__359__A
timestamp 1586364061
transform 1 0 36248 0 1 31008
box -38 -48 222 592
use scs8hd_buf_1  _228_
timestamp 1586364061
transform 1 0 36064 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_6  FILLER_52_390
timestamp 1586364061
transform 1 0 36984 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_52_387
timestamp 1586364061
transform 1 0 36708 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__366__B
timestamp 1586364061
transform 1 0 36800 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__366__A
timestamp 1586364061
transform 1 0 36616 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _366_
timestamp 1586364061
transform 1 0 36800 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_397
timestamp 1586364061
transform 1 0 37628 0 1 31008
box -38 -48 406 592
use scs8hd_decap_4  FILLER_52_401
timestamp 1586364061
transform 1 0 37996 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_396
timestamp 1586364061
transform 1 0 37536 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 37996 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use scs8hd_buf_1  _360_
timestamp 1586364061
transform 1 0 37720 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_403
timestamp 1586364061
transform 1 0 38180 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_407
timestamp 1586364061
transform 1 0 38548 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__365__B
timestamp 1586364061
transform 1 0 38732 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__365__A
timestamp 1586364061
transform 1 0 38364 0 -1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _365_
timestamp 1586364061
transform 1 0 38364 0 1 31008
box -38 -48 866 592
use scs8hd_nor2_4  _363_
timestamp 1586364061
transform 1 0 38916 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_422
timestamp 1586364061
transform 1 0 39928 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_418
timestamp 1586364061
transform 1 0 39560 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_414
timestamp 1586364061
transform 1 0 39192 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_420
timestamp 1586364061
transform 1 0 39744 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39376 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 39744 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_428
timestamp 1586364061
transform 1 0 40480 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_426
timestamp 1586364061
transform 1 0 40296 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 40388 0 1 31008
box -38 -48 130 592
use scs8hd_fill_1  FILLER_52_436
timestamp 1586364061
transform 1 0 41216 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_430
timestamp 1586364061
transform 1 0 40664 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41032 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40848 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41308 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41032 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_447
timestamp 1586364061
transform 1 0 42228 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_443
timestamp 1586364061
transform 1 0 41860 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_446
timestamp 1586364061
transform 1 0 42136 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42320 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_451
timestamp 1586364061
transform 1 0 42596 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_454
timestamp 1586364061
transform 1 0 42872 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_450
timestamp 1586364061
transform 1 0 42504 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_464
timestamp 1586364061
transform 1 0 43792 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_462
timestamp 1586364061
transform 1 0 43608 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_52_457
timestamp 1586364061
transform 1 0 43148 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43976 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 43240 0 -1 31008
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_475
timestamp 1586364061
transform 1 0 44804 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_468
timestamp 1586364061
transform 1 0 44160 0 1 31008
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44344 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44528 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_483
timestamp 1586364061
transform 1 0 45540 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_479
timestamp 1586364061
transform 1 0 45172 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_479
timestamp 1586364061
transform 1 0 45172 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45356 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45908 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45724 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_487
timestamp 1586364061
transform 1 0 45908 0 1 31008
box -38 -48 130 592
use scs8hd_buf_1  _408_
timestamp 1586364061
transform 1 0 46092 0 1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 46000 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_490
timestamp 1586364061
transform 1 0 46184 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_492
timestamp 1586364061
transform 1 0 46368 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__408__A
timestamp 1586364061
transform 1 0 46552 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 46644 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_494
timestamp 1586364061
transform 1 0 46552 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_500
timestamp 1586364061
transform 1 0 47104 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_496
timestamp 1586364061
transform 1 0 46736 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_497
timestamp 1586364061
transform 1 0 46828 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46920 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_509
timestamp 1586364061
transform 1 0 47932 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 48852 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 48852 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_515
timestamp 1586364061
transform 1 0 48484 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_512
timestamp 1586364061
transform 1 0 48208 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_135
timestamp 1586364061
transform 1 0 13524 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_149
timestamp 1586364061
transform 1 0 14812 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_163
timestamp 1586364061
transform 1 0 16100 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_167
timestamp 1586364061
transform 1 0 16468 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_8  FILLER_54_174
timestamp 1586364061
transform 1 0 17112 0 -1 32096
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_191
timestamp 1586364061
transform 1 0 18676 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_199
timestamp 1586364061
transform 1 0 19412 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_203
timestamp 1586364061
transform 1 0 19780 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_54_211
timestamp 1586364061
transform 1 0 20516 0 -1 32096
box -38 -48 314 592
use scs8hd_nor2_4  _476_
timestamp 1586364061
transform 1 0 22724 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_224
timestamp 1586364061
transform 1 0 21712 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_228
timestamp 1586364061
transform 1 0 22080 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_54_234
timestamp 1586364061
transform 1 0 22632 0 -1 32096
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_244
timestamp 1586364061
transform 1 0 23552 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_252
timestamp 1586364061
transform 1 0 24288 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_255
timestamp 1586364061
transform 1 0 24564 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_54_267
timestamp 1586364061
transform 1 0 25668 0 -1 32096
box -38 -48 774 592
use scs8hd_conb_1  _644_
timestamp 1586364061
transform 1 0 27232 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_276
timestamp 1586364061
transform 1 0 26496 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_54_287
timestamp 1586364061
transform 1 0 27508 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_291
timestamp 1586364061
transform 1 0 27876 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_301
timestamp 1586364061
transform 1 0 28796 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_297
timestamp 1586364061
transform 1 0 28428 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28612 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__474__B
timestamp 1586364061
transform 1 0 28980 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _480_
timestamp 1586364061
transform 1 0 29164 0 -1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_54_314
timestamp 1586364061
transform 1 0 29992 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_318
timestamp 1586364061
transform 1 0 30360 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__481__B
timestamp 1586364061
transform 1 0 30544 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__481__A
timestamp 1586364061
transform 1 0 30176 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30728 0 -1 32096
box -38 -48 314 592
use scs8hd_or4_4  _471_
timestamp 1586364061
transform 1 0 32108 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__471__D
timestamp 1586364061
transform 1 0 31832 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__A
timestamp 1586364061
transform 1 0 31464 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__C
timestamp 1586364061
transform 1 0 33120 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_325
timestamp 1586364061
transform 1 0 31004 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_329
timestamp 1586364061
transform 1 0 31372 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_332
timestamp 1586364061
transform 1 0 31648 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_346
timestamp 1586364061
transform 1 0 32936 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_8  _316_
timestamp 1586364061
transform 1 0 34500 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__383__B
timestamp 1586364061
transform 1 0 33672 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__D
timestamp 1586364061
transform 1 0 35512 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__D
timestamp 1586364061
transform 1 0 34316 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_350
timestamp 1586364061
transform 1 0 33304 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_4  FILLER_54_356
timestamp 1586364061
transform 1 0 33856 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_360
timestamp 1586364061
transform 1 0 34224 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_372
timestamp 1586364061
transform 1 0 35328 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_387
timestamp 1586364061
transform 1 0 36708 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_380
timestamp 1586364061
transform 1 0 36064 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_376
timestamp 1586364061
transform 1 0 35696 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__B
timestamp 1586364061
transform 1 0 36248 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__C
timestamp 1586364061
transform 1 0 35880 0 -1 32096
box -38 -48 222 592
use scs8hd_buf_1  _359_
timestamp 1586364061
transform 1 0 36432 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_54_398
timestamp 1586364061
transform 1 0 37720 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_395
timestamp 1586364061
transform 1 0 37444 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_391
timestamp 1586364061
transform 1 0 37076 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__C
timestamp 1586364061
transform 1 0 37260 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__B
timestamp 1586364061
transform 1 0 36892 0 -1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 37996 0 -1 32096
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 39744 0 -1 32096
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_54_412
timestamp 1586364061
transform 1 0 39008 0 -1 32096
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41492 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42780 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_431
timestamp 1586364061
transform 1 0 40756 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_54_436
timestamp 1586364061
transform 1 0 41216 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_448
timestamp 1586364061
transform 1 0 42320 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_452
timestamp 1586364061
transform 1 0 42688 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_455
timestamp 1586364061
transform 1 0 42964 0 -1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44896 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 43240 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_468
timestamp 1586364061
transform 1 0 44160 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_472
timestamp 1586364061
transform 1 0 44528 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_54_475
timestamp 1586364061
transform 1 0 44804 0 -1 32096
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46460 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 46092 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_485
timestamp 1586364061
transform 1 0 45724 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_491
timestamp 1586364061
transform 1 0 46276 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_54_496
timestamp 1586364061
transform 1 0 46736 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_508
timestamp 1586364061
transform 1 0 47840 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 48852 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__445__A
timestamp 1586364061
transform 1 0 13156 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__445__B
timestamp 1586364061
transform 1 0 12788 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_129
timestamp 1586364061
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14352 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_136
timestamp 1586364061
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_140
timestamp 1586364061
transform 1 0 13984 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_155
timestamp 1586364061
transform 1 0 15364 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_159
timestamp 1586364061
transform 1 0 15732 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_168
timestamp 1586364061
transform 1 0 16560 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_163
timestamp 1586364061
transform 1 0 16100 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__446__B
timestamp 1586364061
transform 1 0 16376 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__440__A
timestamp 1586364061
transform 1 0 16744 0 1 32096
box -38 -48 222 592
use scs8hd_buf_1  _440_
timestamp 1586364061
transform 1 0 16928 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_179
timestamp 1586364061
transform 1 0 17572 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_175
timestamp 1586364061
transform 1 0 17204 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__446__A
timestamp 1586364061
transform 1 0 17388 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 32096
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_195
timestamp 1586364061
transform 1 0 19044 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_199
timestamp 1586364061
transform 1 0 19412 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_203
timestamp 1586364061
transform 1 0 19780 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_209
timestamp 1586364061
transform 1 0 20332 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_213
timestamp 1586364061
transform 1 0 20700 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21068 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_228
timestamp 1586364061
transform 1 0 22080 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_232
timestamp 1586364061
transform 1 0 22448 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_236
timestamp 1586364061
transform 1 0 22816 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_249
timestamp 1586364061
transform 1 0 24012 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_245
timestamp 1586364061
transform 1 0 23644 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_242
timestamp 1586364061
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23828 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 1 32096
box -38 -48 866 592
use scs8hd_decap_6  FILLER_55_266
timestamp 1586364061
transform 1 0 25576 0 1 32096
box -38 -48 590 592
use scs8hd_fill_2  FILLER_55_262
timestamp 1586364061
transform 1 0 25208 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26312 0 1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_277
timestamp 1586364061
transform 1 0 26588 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_281
timestamp 1586364061
transform 1 0 26956 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_294
timestamp 1586364061
transform 1 0 28152 0 1 32096
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 29256 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__A
timestamp 1586364061
transform 1 0 30544 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28428 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_299
timestamp 1586364061
transform 1 0 28612 0 1 32096
box -38 -48 406 592
use scs8hd_decap_3  FILLER_55_317
timestamp 1586364061
transform 1 0 30268 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_322
timestamp 1586364061
transform 1 0 30728 0 1 32096
box -38 -48 222 592
use scs8hd_or4_4  _385_
timestamp 1586364061
transform 1 0 31832 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__409__D
timestamp 1586364061
transform 1 0 32844 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__D
timestamp 1586364061
transform 1 0 31648 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__B
timestamp 1586364061
transform 1 0 31280 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__B
timestamp 1586364061
transform 1 0 30912 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_326
timestamp 1586364061
transform 1 0 31096 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_330
timestamp 1586364061
transform 1 0 31464 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_343
timestamp 1586364061
transform 1 0 32660 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_347
timestamp 1586364061
transform 1 0 33028 0 1 32096
box -38 -48 222 592
use scs8hd_or2_4  _317_
timestamp 1586364061
transform 1 0 33396 0 1 32096
box -38 -48 682 592
use scs8hd_or4_4  _396_
timestamp 1586364061
transform 1 0 34868 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__317__B
timestamp 1586364061
transform 1 0 34224 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__383__A
timestamp 1586364061
transform 1 0 33212 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__B
timestamp 1586364061
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_358
timestamp 1586364061
transform 1 0 34040 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_362
timestamp 1586364061
transform 1 0 34408 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_380
timestamp 1586364061
transform 1 0 36064 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_376
timestamp 1586364061
transform 1 0 35696 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__A
timestamp 1586364061
transform 1 0 36248 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__A
timestamp 1586364061
transform 1 0 35880 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _367_
timestamp 1586364061
transform 1 0 36432 0 1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_55_397
timestamp 1586364061
transform 1 0 37628 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_393
timestamp 1586364061
transform 1 0 37260 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__368__A
timestamp 1586364061
transform 1 0 37444 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 37812 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 37996 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 40388 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__368__B
timestamp 1586364061
transform 1 0 39192 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_412
timestamp 1586364061
transform 1 0 39008 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_416
timestamp 1586364061
transform 1 0 39376 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_420
timestamp 1586364061
transform 1 0 39744 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_423
timestamp 1586364061
transform 1 0 40020 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_428
timestamp 1586364061
transform 1 0 40480 0 1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42780 0 1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41032 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42596 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40848 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_443
timestamp 1586364061
transform 1 0 41860 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_447
timestamp 1586364061
transform 1 0 42228 0 1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44344 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43792 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45356 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44160 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_462
timestamp 1586364061
transform 1 0 43608 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_466
timestamp 1586364061
transform 1 0 43976 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_479
timestamp 1586364061
transform 1 0 45172 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_483
timestamp 1586364061
transform 1 0 45540 0 1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 46092 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 46000 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45816 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 47104 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_498
timestamp 1586364061
transform 1 0 46920 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_502
timestamp 1586364061
transform 1 0 47288 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 48852 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_514
timestamp 1586364061
transform 1 0 48392 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 590 592
use scs8hd_nor2_4  _445_
timestamp 1586364061
transform 1 0 13616 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_135
timestamp 1586364061
transform 1 0 13524 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _446_
timestamp 1586364061
transform 1 0 16836 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__448__A
timestamp 1586364061
transform 1 0 18308 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17848 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_163
timestamp 1586364061
transform 1 0 16100 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_180
timestamp 1586364061
transform 1 0 17664 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_184
timestamp 1586364061
transform 1 0 18032 0 -1 33184
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_189
timestamp 1586364061
transform 1 0 18492 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_193
timestamp 1586364061
transform 1 0 18860 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_206
timestamp 1586364061
transform 1 0 20056 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_210
timestamp 1586364061
transform 1 0 20424 0 -1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 33184
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_12  FILLER_56_224
timestamp 1586364061
transform 1 0 21712 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_236
timestamp 1586364061
transform 1 0 22816 0 -1 33184
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_251
timestamp 1586364061
transform 1 0 24196 0 -1 33184
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_56_263
timestamp 1586364061
transform 1 0 25300 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_6  FILLER_56_267
timestamp 1586364061
transform 1 0 25668 0 -1 33184
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_285
timestamp 1586364061
transform 1 0 27324 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_289
timestamp 1586364061
transform 1 0 27692 0 -1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _481_
timestamp 1586364061
transform 1 0 29992 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28428 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29624 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_306
timestamp 1586364061
transform 1 0 29256 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_56_312
timestamp 1586364061
transform 1 0 29808 0 -1 33184
box -38 -48 222 592
use scs8hd_or4_4  _409_
timestamp 1586364061
transform 1 0 32108 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__385__A
timestamp 1586364061
transform 1 0 31832 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__C
timestamp 1586364061
transform 1 0 31464 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__C
timestamp 1586364061
transform 1 0 31096 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_323
timestamp 1586364061
transform 1 0 30820 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_328
timestamp 1586364061
transform 1 0 31280 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_332
timestamp 1586364061
transform 1 0 31648 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_346
timestamp 1586364061
transform 1 0 32936 0 -1 33184
box -38 -48 406 592
use scs8hd_or4_4  _358_
timestamp 1586364061
transform 1 0 35236 0 -1 33184
box -38 -48 866 592
use scs8hd_nand2_4  _383_
timestamp 1586364061
transform 1 0 33672 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__346__A
timestamp 1586364061
transform 1 0 34960 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__317__A
timestamp 1586364061
transform 1 0 33396 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_350
timestamp 1586364061
transform 1 0 33304 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_353
timestamp 1586364061
transform 1 0 33580 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_363
timestamp 1586364061
transform 1 0 34500 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_367
timestamp 1586364061
transform 1 0 34868 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_370
timestamp 1586364061
transform 1 0 35144 0 -1 33184
box -38 -48 130 592
use scs8hd_nor2_4  _368_
timestamp 1586364061
transform 1 0 37720 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__369__B
timestamp 1586364061
transform 1 0 36432 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__D
timestamp 1586364061
transform 1 0 36800 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__C
timestamp 1586364061
transform 1 0 37168 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_380
timestamp 1586364061
transform 1 0 36064 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_56_386
timestamp 1586364061
transform 1 0 36616 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_390
timestamp 1586364061
transform 1 0 36984 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_394
timestamp 1586364061
transform 1 0 37352 0 -1 33184
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39836 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38732 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_407
timestamp 1586364061
transform 1 0 38548 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_411
timestamp 1586364061
transform 1 0 38916 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_419
timestamp 1586364061
transform 1 0 39652 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_424
timestamp 1586364061
transform 1 0 40112 0 -1 33184
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40848 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_12  FILLER_56_441
timestamp 1586364061
transform 1 0 41676 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_453
timestamp 1586364061
transform 1 0 42780 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_4  FILLER_56_465
timestamp 1586364061
transform 1 0 43884 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_3  FILLER_56_459
timestamp 1586364061
transform 1 0 43332 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_457
timestamp 1586364061
transform 1 0 43148 0 -1 33184
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 43240 0 -1 33184
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43608 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_472
timestamp 1586364061
transform 1 0 44528 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_469
timestamp 1586364061
transform 1 0 44252 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44620 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_8  FILLER_56_482
timestamp 1586364061
transform 1 0 45448 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46184 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_493
timestamp 1586364061
transform 1 0 46460 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_56_505
timestamp 1586364061
transform 1 0 47564 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 48852 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_513
timestamp 1586364061
transform 1 0 48300 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_nor2_4  _416_
timestamp 1586364061
transform 1 0 15272 0 1 33184
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__B
timestamp 1586364061
transform 1 0 15088 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_146
timestamp 1586364061
transform 1 0 14536 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_150
timestamp 1586364061
transform 1 0 14904 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_167
timestamp 1586364061
transform 1 0 16468 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_163
timestamp 1586364061
transform 1 0 16100 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16284 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_179
timestamp 1586364061
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_175
timestamp 1586364061
transform 1 0 17204 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_171
timestamp 1586364061
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_184
timestamp 1586364061
transform 1 0 18032 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__448__B
timestamp 1586364061
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use scs8hd_nor2_4  _448_
timestamp 1586364061
transform 1 0 18308 0 1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_196
timestamp 1586364061
transform 1 0 19136 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_200
timestamp 1586364061
transform 1 0 19504 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_213
timestamp 1586364061
transform 1 0 20700 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_217
timestamp 1586364061
transform 1 0 21068 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__447__A
timestamp 1586364061
transform 1 0 21252 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _447_
timestamp 1586364061
transform 1 0 21436 0 1 33184
box -38 -48 866 592
use scs8hd_fill_1  FILLER_57_234
timestamp 1586364061
transform 1 0 22632 0 1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_57_230
timestamp 1586364061
transform 1 0 22264 0 1 33184
box -38 -48 406 592
use scs8hd_decap_3  FILLER_57_241
timestamp 1586364061
transform 1 0 23276 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_237
timestamp 1586364061
transform 1 0 22908 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__479__B
timestamp 1586364061
transform 1 0 23092 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__479__A
timestamp 1586364061
transform 1 0 22724 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 33184
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_245
timestamp 1586364061
transform 1 0 23644 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_258
timestamp 1586364061
transform 1 0 24840 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_262
timestamp 1586364061
transform 1 0 25208 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_273
timestamp 1586364061
transform 1 0 26220 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_269
timestamp 1586364061
transform 1 0 25852 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_57_287
timestamp 1586364061
transform 1 0 27508 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_295
timestamp 1586364061
transform 1 0 28244 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_291
timestamp 1586364061
transform 1 0 27876 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 29716 0 1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 29532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28428 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_299
timestamp 1586364061
transform 1 0 28612 0 1 33184
box -38 -48 406 592
use scs8hd_decap_3  FILLER_57_306
timestamp 1586364061
transform 1 0 29256 0 1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_57_322
timestamp 1586364061
transform 1 0 30728 0 1 33184
box -38 -48 406 592
use scs8hd_or4_4  _427_
timestamp 1586364061
transform 1 0 31740 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__406__A
timestamp 1586364061
transform 1 0 32752 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__D
timestamp 1586364061
transform 1 0 31556 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__C
timestamp 1586364061
transform 1 0 31188 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_326
timestamp 1586364061
transform 1 0 31096 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_329
timestamp 1586364061
transform 1 0 31372 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_342
timestamp 1586364061
transform 1 0 32568 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_346
timestamp 1586364061
transform 1 0 32936 0 1 33184
box -38 -48 314 592
use scs8hd_or4_4  _320_
timestamp 1586364061
transform 1 0 34868 0 1 33184
box -38 -48 866 592
use scs8hd_or2_4  _357_
timestamp 1586364061
transform 1 0 33396 0 1 33184
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__357__A
timestamp 1586364061
transform 1 0 34224 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__357__B
timestamp 1586364061
transform 1 0 33212 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_358
timestamp 1586364061
transform 1 0 34040 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_362
timestamp 1586364061
transform 1 0 34408 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_380
timestamp 1586364061
transform 1 0 36064 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_376
timestamp 1586364061
transform 1 0 35696 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__320__A
timestamp 1586364061
transform 1 0 35880 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__A
timestamp 1586364061
transform 1 0 36248 0 1 33184
box -38 -48 222 592
use scs8hd_or4_4  _369_
timestamp 1586364061
transform 1 0 36432 0 1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_57_393
timestamp 1586364061
transform 1 0 37260 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__C
timestamp 1586364061
transform 1 0 37444 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_397
timestamp 1586364061
transform 1 0 37628 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__349__B
timestamp 1586364061
transform 1 0 37812 0 1 33184
box -38 -48 222 592
use scs8hd_buf_1  _380_
timestamp 1586364061
transform 1 0 37996 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_404
timestamp 1586364061
transform 1 0 38272 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__349__A
timestamp 1586364061
transform 1 0 38456 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_412
timestamp 1586364061
transform 1 0 39008 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_408
timestamp 1586364061
transform 1 0 38640 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__380__A
timestamp 1586364061
transform 1 0 38824 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_419
timestamp 1586364061
transform 1 0 39652 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_423
timestamp 1586364061
transform 1 0 40020 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_428
timestamp 1586364061
transform 1 0 40480 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 40388 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_433
timestamp 1586364061
transform 1 0 40940 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40664 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_437
timestamp 1586364061
transform 1 0 41308 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_441
timestamp 1586364061
transform 1 0 41676 0 1 33184
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41768 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_445
timestamp 1586364061
transform 1 0 42044 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_449
timestamp 1586364061
transform 1 0 42412 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_456
timestamp 1586364061
transform 1 0 43056 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42780 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_460
timestamp 1586364061
transform 1 0 43424 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43240 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_464
timestamp 1586364061
transform 1 0 43792 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_468
timestamp 1586364061
transform 1 0 44160 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43976 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_474
timestamp 1586364061
transform 1 0 44712 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44436 0 1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_57_478
timestamp 1586364061
transform 1 0 45080 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44896 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_482
timestamp 1586364061
transform 1 0 45448 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45540 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 46000 0 1 33184
box -38 -48 130 592
use scs8hd_decap_3  FILLER_57_485
timestamp 1586364061
transform 1 0 45724 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_489
timestamp 1586364061
transform 1 0 46092 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_501
timestamp 1586364061
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 48852 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_513
timestamp 1586364061
transform 1 0 48300 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__414__A
timestamp 1586364061
transform 1 0 13248 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_134
timestamp 1586364061
transform 1 0 13432 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__416__A
timestamp 1586364061
transform 1 0 15456 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_146
timestamp 1586364061
transform 1 0 14536 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_151
timestamp 1586364061
transform 1 0 14996 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_154
timestamp 1586364061
transform 1 0 15272 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_158
timestamp 1586364061
transform 1 0 15640 0 -1 34272
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 34272
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_173
timestamp 1586364061
transform 1 0 17020 0 -1 34272
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_190
timestamp 1586364061
transform 1 0 18584 0 -1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_58_198
timestamp 1586364061
transform 1 0 19320 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_202
timestamp 1586364061
transform 1 0 19688 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_206
timestamp 1586364061
transform 1 0 20056 0 -1 34272
box -38 -48 774 592
use scs8hd_nor2_4  _479_
timestamp 1586364061
transform 1 0 22724 0 -1 34272
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__447__B
timestamp 1586364061
transform 1 0 21436 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_218
timestamp 1586364061
transform 1 0 21160 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_223
timestamp 1586364061
transform 1 0 21620 0 -1 34272
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_244
timestamp 1586364061
transform 1 0 23552 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_248
timestamp 1586364061
transform 1 0 23920 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_251
timestamp 1586364061
transform 1 0 24196 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_264
timestamp 1586364061
transform 1 0 25392 0 -1 34272
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_272
timestamp 1586364061
transform 1 0 26128 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_285
timestamp 1586364061
transform 1 0 27324 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_289
timestamp 1586364061
transform 1 0 27692 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29624 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_302
timestamp 1586364061
transform 1 0 28888 0 -1 34272
box -38 -48 590 592
use scs8hd_decap_6  FILLER_58_319
timestamp 1586364061
transform 1 0 30452 0 -1 34272
box -38 -48 590 592
use scs8hd_nor2_4  _406_
timestamp 1586364061
transform 1 0 32108 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__427__B
timestamp 1586364061
transform 1 0 31740 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__406__B
timestamp 1586364061
transform 1 0 31372 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__A
timestamp 1586364061
transform 1 0 31004 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_327
timestamp 1586364061
transform 1 0 31188 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_331
timestamp 1586364061
transform 1 0 31556 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_335
timestamp 1586364061
transform 1 0 31924 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_346
timestamp 1586364061
transform 1 0 32936 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_353
timestamp 1586364061
transform 1 0 33580 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_350
timestamp 1586364061
transform 1 0 33304 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__320__D
timestamp 1586364061
transform 1 0 33396 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__320__C
timestamp 1586364061
transform 1 0 33764 0 -1 34272
box -38 -48 222 592
use scs8hd_buf_1  _226_
timestamp 1586364061
transform 1 0 33948 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_367
timestamp 1586364061
transform 1 0 34868 0 -1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_58_364
timestamp 1586364061
transform 1 0 34592 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_360
timestamp 1586364061
transform 1 0 34224 0 -1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 34684 0 -1 34272
box -38 -48 222 592
use scs8hd_or4_4  _346_
timestamp 1586364061
transform 1 0 34960 0 -1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_58_381
timestamp 1586364061
transform 1 0 36156 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_377
timestamp 1586364061
transform 1 0 35788 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__320__B
timestamp 1586364061
transform 1 0 36340 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__B
timestamp 1586364061
transform 1 0 35972 0 -1 34272
box -38 -48 222 592
use scs8hd_buf_1  _347_
timestamp 1586364061
transform 1 0 36524 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_392
timestamp 1586364061
transform 1 0 37168 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_388
timestamp 1586364061
transform 1 0 36800 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__A
timestamp 1586364061
transform 1 0 36984 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_398
timestamp 1586364061
transform 1 0 37720 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_58_396
timestamp 1586364061
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37904 0 -1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use scs8hd_nor2_4  _349_
timestamp 1586364061
transform 1 0 38088 0 -1 34272
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39928 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 40572 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39100 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_411
timestamp 1586364061
transform 1 0 38916 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_415
timestamp 1586364061
transform 1 0 39284 0 -1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_58_421
timestamp 1586364061
transform 1 0 39836 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_425
timestamp 1586364061
transform 1 0 40204 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_431
timestamp 1586364061
transform 1 0 40756 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_442
timestamp 1586364061
transform 1 0 41768 0 -1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_58_448
timestamp 1586364061
transform 1 0 42320 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_451
timestamp 1586364061
transform 1 0 42596 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_455
timestamp 1586364061
transform 1 0 42964 0 -1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45540 0 -1 34272
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 43240 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44620 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_459
timestamp 1586364061
transform 1 0 43332 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_471
timestamp 1586364061
transform 1 0 44436 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_475
timestamp 1586364061
transform 1 0 44804 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_58_486
timestamp 1586364061
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_498
timestamp 1586364061
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 48852 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_6  FILLER_58_510
timestamp 1586364061
transform 1 0 48024 0 -1 34272
box -38 -48 590 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_60_133
timestamp 1586364061
transform 1 0 13340 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_129
timestamp 1586364061
transform 1 0 12972 0 1 34272
box -38 -48 130 592
use scs8hd_decap_6  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__418__A
timestamp 1586364061
transform 1 0 13156 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__414__B
timestamp 1586364061
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_nor2_4  _414_
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_146
timestamp 1586364061
transform 1 0 14536 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_138
timestamp 1586364061
transform 1 0 13800 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_6  FILLER_59_141
timestamp 1586364061
transform 1 0 14076 0 1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__420__A
timestamp 1586364061
transform 1 0 13616 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_157
timestamp 1586364061
transform 1 0 15548 0 -1 35360
box -38 -48 590 592
use scs8hd_decap_3  FILLER_60_150
timestamp 1586364061
transform 1 0 14904 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 14812 0 1 34272
box -38 -48 1050 592
use scs8hd_buf_1  _411_
timestamp 1586364061
transform 1 0 15272 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_160
timestamp 1586364061
transform 1 0 15824 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_168
timestamp 1586364061
transform 1 0 16560 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_164
timestamp 1586364061
transform 1 0 16192 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__411__A
timestamp 1586364061
transform 1 0 16008 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_174
timestamp 1586364061
transform 1 0 17112 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_179
timestamp 1586364061
transform 1 0 17572 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_175
timestamp 1586364061
transform 1 0 17204 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_184
timestamp 1586364061
transform 1 0 18032 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_184
timestamp 1586364061
transform 1 0 18032 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__A
timestamp 1586364061
transform 1 0 17848 0 -1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_200
timestamp 1586364061
transform 1 0 19504 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_60_188
timestamp 1586364061
transform 1 0 18400 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_192
timestamp 1586364061
transform 1 0 18768 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_188
timestamp 1586364061
transform 1 0 18400 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 34272
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_60_212
timestamp 1586364061
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_209
timestamp 1586364061
transform 1 0 20332 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_205
timestamp 1586364061
transform 1 0 19964 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_219
timestamp 1586364061
transform 1 0 21252 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_60_215
timestamp 1586364061
transform 1 0 20884 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  FILLER_59_222
timestamp 1586364061
transform 1 0 21528 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 1 34272
box -38 -48 222 592
use scs8hd_conb_1  _649_
timestamp 1586364061
transform 1 0 20976 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_227
timestamp 1586364061
transform 1 0 21988 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_236
timestamp 1586364061
transform 1 0 22816 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_231
timestamp 1586364061
transform 1 0 22356 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_227
timestamp 1586364061
transform 1 0 21988 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 22172 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 34272
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 35360
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_60_240
timestamp 1586364061
transform 1 0 23184 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_240
timestamp 1586364061
transform 1 0 23184 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_248
timestamp 1586364061
transform 1 0 23920 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 35360
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_60_257
timestamp 1586364061
transform 1 0 24748 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_6  FILLER_59_256
timestamp 1586364061
transform 1 0 24656 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_252
timestamp 1586364061
transform 1 0 24288 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_267
timestamp 1586364061
transform 1 0 25668 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_262
timestamp 1586364061
transform 1 0 25208 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25484 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_276
timestamp 1586364061
transform 1 0 26496 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_271
timestamp 1586364061
transform 1 0 26036 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_8  FILLER_59_274
timestamp 1586364061
transform 1 0 26312 0 1 34272
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_287
timestamp 1586364061
transform 1 0 27508 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_60_280
timestamp 1586364061
transform 1 0 26864 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_4  FILLER_59_286
timestamp 1586364061
transform 1 0 27416 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_282
timestamp 1586364061
transform 1 0 27048 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27232 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27232 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_295
timestamp 1586364061
transform 1 0 28244 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27784 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 35360
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27968 0 1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_304
timestamp 1586364061
transform 1 0 29072 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_303
timestamp 1586364061
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_299
timestamp 1586364061
transform 1 0 28612 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28796 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28428 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_318
timestamp 1586364061
transform 1 0 30360 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_320
timestamp 1586364061
transform 1 0 30544 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_313
timestamp 1586364061
transform 1 0 29900 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_309
timestamp 1586364061
transform 1 0 29532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30176 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__B
timestamp 1586364061
transform 1 0 30084 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30268 0 1 34272
box -38 -48 314 592
use scs8hd_nor2_4  _404_
timestamp 1586364061
transform 1 0 30452 0 -1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_328
timestamp 1586364061
transform 1 0 31280 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_331
timestamp 1586364061
transform 1 0 31556 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_324
timestamp 1586364061
transform 1 0 30912 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__A
timestamp 1586364061
transform 1 0 31096 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_345
timestamp 1586364061
transform 1 0 32844 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_341
timestamp 1586364061
transform 1 0 32476 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_337
timestamp 1586364061
transform 1 0 32108 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_335
timestamp 1586364061
transform 1 0 31924 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__405__B
timestamp 1586364061
transform 1 0 32292 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__405__A
timestamp 1586364061
transform 1 0 32108 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use scs8hd_nor2_4  _405_
timestamp 1586364061
transform 1 0 32292 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_59_348
timestamp 1586364061
transform 1 0 33120 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32936 0 -1 35360
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_60_357
timestamp 1586364061
transform 1 0 33948 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_356
timestamp 1586364061
transform 1 0 33856 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_352
timestamp 1586364061
transform 1 0 33488 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 33304 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_367
timestamp 1586364061
transform 1 0 34868 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_362
timestamp 1586364061
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__315__A
timestamp 1586364061
transform 1 0 34224 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use scs8hd_inv_8  _315_
timestamp 1586364061
transform 1 0 34960 0 1 34272
box -38 -48 866 592
use scs8hd_or2_4  _227_
timestamp 1586364061
transform 1 0 34684 0 -1 35360
box -38 -48 682 592
use scs8hd_fill_2  FILLER_60_372
timestamp 1586364061
transform 1 0 35328 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__D
timestamp 1586364061
transform 1 0 35512 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_376
timestamp 1586364061
transform 1 0 35696 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  FILLER_59_386
timestamp 1586364061
transform 1 0 36616 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_382
timestamp 1586364061
transform 1 0 36248 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_377
timestamp 1586364061
transform 1 0 35788 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__356__B
timestamp 1586364061
transform 1 0 36432 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__356__A
timestamp 1586364061
transform 1 0 36064 0 1 34272
box -38 -48 222 592
use scs8hd_nor2_4  _356_
timestamp 1586364061
transform 1 0 36064 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_3  FILLER_60_398
timestamp 1586364061
transform 1 0 37720 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_393
timestamp 1586364061
transform 1 0 37260 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_389
timestamp 1586364061
transform 1 0 36892 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__B
timestamp 1586364061
transform 1 0 37076 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__A
timestamp 1586364061
transform 1 0 36892 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use scs8hd_nor2_4  _350_
timestamp 1586364061
transform 1 0 37076 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_59_400
timestamp 1586364061
transform 1 0 37904 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38088 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 37996 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_60_412
timestamp 1586364061
transform 1 0 39008 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_404
timestamp 1586364061
transform 1 0 38272 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__B
timestamp 1586364061
transform 1 0 39192 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 38640 0 1 34272
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_60_428
timestamp 1586364061
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_416
timestamp 1586364061
transform 1 0 39376 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_428
timestamp 1586364061
transform 1 0 40480 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_423
timestamp 1586364061
transform 1 0 40020 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_419
timestamp 1586364061
transform 1 0 39652 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 40572 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_60_440
timestamp 1586364061
transform 1 0 41584 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_441
timestamp 1586364061
transform 1 0 41676 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 -1 35360
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40664 0 1 34272
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_60_444
timestamp 1586364061
transform 1 0 41952 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_445
timestamp 1586364061
transform 1 0 42044 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41860 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42412 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_456
timestamp 1586364061
transform 1 0 43056 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_462
timestamp 1586364061
transform 1 0 43608 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_458
timestamp 1586364061
transform 1 0 43240 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43424 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43976 0 1 34272
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_472
timestamp 1586364061
transform 1 0 44528 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_468
timestamp 1586364061
transform 1 0 44160 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_475
timestamp 1586364061
transform 1 0 44804 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_483
timestamp 1586364061
transform 1 0 45540 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_479
timestamp 1586364061
transform 1 0 45172 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45356 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44988 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44896 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_485
timestamp 1586364061
transform 1 0 45724 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_492
timestamp 1586364061
transform 1 0 46368 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_487
timestamp 1586364061
transform 1 0 45908 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46460 0 -1 35360
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_60_508
timestamp 1586364061
transform 1 0 47840 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_496
timestamp 1586364061
transform 1 0 46736 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_500
timestamp 1586364061
transform 1 0 47104 0 1 34272
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_496
timestamp 1586364061
transform 1 0 46736 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46920 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 48852 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 48852 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_59_512
timestamp 1586364061
transform 1 0 48208 0 1 34272
box -38 -48 406 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_nor2_4  _418_
timestamp 1586364061
transform 1 0 13156 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__418__B
timestamp 1586364061
transform 1 0 12972 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14720 0 1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__420__B
timestamp 1586364061
transform 1 0 14168 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_140
timestamp 1586364061
transform 1 0 13984 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_144
timestamp 1586364061
transform 1 0 14352 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_159
timestamp 1586364061
transform 1 0 15732 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_163
timestamp 1586364061
transform 1 0 16100 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_167
timestamp 1586364061
transform 1 0 16468 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_171
timestamp 1586364061
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_175
timestamp 1586364061
transform 1 0 17204 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_179
timestamp 1586364061
transform 1 0 17572 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_184
timestamp 1586364061
transform 1 0 18032 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__422__B
timestamp 1586364061
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_192
timestamp 1586364061
transform 1 0 18768 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_188
timestamp 1586364061
transform 1 0 18400 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 35360
box -38 -48 866 592
use scs8hd_fill_2  FILLER_61_205
timestamp 1586364061
transform 1 0 19964 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_214
timestamp 1586364061
transform 1 0 20792 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_209
timestamp 1586364061
transform 1 0 20332 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__412__A
timestamp 1586364061
transform 1 0 22172 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__B
timestamp 1586364061
transform 1 0 20976 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_227
timestamp 1586364061
transform 1 0 21988 0 1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_61_231
timestamp 1586364061
transform 1 0 22356 0 1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_61_237
timestamp 1586364061
transform 1 0 22908 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_240
timestamp 1586364061
transform 1 0 23184 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_248
timestamp 1586364061
transform 1 0 23920 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_260
timestamp 1586364061
transform 1 0 25024 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_252
timestamp 1586364061
transform 1 0 24288 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_264
timestamp 1586364061
transform 1 0 25392 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25576 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25760 0 1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_277
timestamp 1586364061
transform 1 0 26588 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_281
timestamp 1586364061
transform 1 0 26956 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_285
timestamp 1586364061
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_297
timestamp 1586364061
transform 1 0 28428 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_301
timestamp 1586364061
transform 1 0 28796 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_309
timestamp 1586364061
transform 1 0 29532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_313
timestamp 1586364061
transform 1 0 29900 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_318
timestamp 1586364061
transform 1 0 30360 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30176 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_322
timestamp 1586364061
transform 1 0 30728 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30544 0 1 35360
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32844 0 1 35360
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 31096 0 1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30912 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32660 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32292 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_337
timestamp 1586364061
transform 1 0 32108 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_341
timestamp 1586364061
transform 1 0 32476 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__355__B
timestamp 1586364061
transform 1 0 35604 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34040 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34408 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_356
timestamp 1586364061
transform 1 0 33856 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_360
timestamp 1586364061
transform 1 0 34224 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_364
timestamp 1586364061
transform 1 0 34592 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_367
timestamp 1586364061
transform 1 0 34868 0 1 35360
box -38 -48 774 592
use scs8hd_buf_1  _348_
timestamp 1586364061
transform 1 0 35788 0 1 35360
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 36800 0 1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 36616 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__355__A
timestamp 1586364061
transform 1 0 36248 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_380
timestamp 1586364061
transform 1 0 36064 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_384
timestamp 1586364061
transform 1 0 36432 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_399
timestamp 1586364061
transform 1 0 37812 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_406
timestamp 1586364061
transform 1 0 38456 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_403
timestamp 1586364061
transform 1 0 38180 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__351__B
timestamp 1586364061
transform 1 0 38272 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__351__A
timestamp 1586364061
transform 1 0 38640 0 1 35360
box -38 -48 222 592
use scs8hd_nor2_4  _351_
timestamp 1586364061
transform 1 0 38824 0 1 35360
box -38 -48 866 592
use scs8hd_fill_2  FILLER_61_419
timestamp 1586364061
transform 1 0 39652 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__A
timestamp 1586364061
transform 1 0 39836 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_423
timestamp 1586364061
transform 1 0 40020 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41584 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41308 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_431
timestamp 1586364061
transform 1 0 40756 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_435
timestamp 1586364061
transform 1 0 41124 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_439
timestamp 1586364061
transform 1 0 41492 0 1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_61_449
timestamp 1586364061
transform 1 0 42412 0 1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_61_464
timestamp 1586364061
transform 1 0 43792 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_460
timestamp 1586364061
transform 1 0 43424 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43976 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43608 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43148 0 1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44160 0 1 35360
box -38 -48 866 592
use scs8hd_fill_2  FILLER_61_481
timestamp 1586364061
transform 1 0 45356 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_477
timestamp 1586364061
transform 1 0 44988 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45540 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45172 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46368 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_485
timestamp 1586364061
transform 1 0 45724 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_489
timestamp 1586364061
transform 1 0 46092 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_494
timestamp 1586364061
transform 1 0 46552 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_506
timestamp 1586364061
transform 1 0 47656 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 48852 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_514
timestamp 1586364061
transform 1 0 48392 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_62_135
timestamp 1586364061
transform 1 0 13524 0 -1 36448
box -38 -48 130 592
use scs8hd_nor2_4  _420_
timestamp 1586364061
transform 1 0 13616 0 -1 36448
box -38 -48 866 592
use scs8hd_fill_2  FILLER_62_149
timestamp 1586364061
transform 1 0 14812 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_157
timestamp 1586364061
transform 1 0 15548 0 -1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 -1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 36448
box -38 -48 314 592
use scs8hd_nor2_4  _422_
timestamp 1586364061
transform 1 0 17848 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_163
timestamp 1586364061
transform 1 0 16100 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_62_174
timestamp 1586364061
transform 1 0 17112 0 -1 36448
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_191
timestamp 1586364061
transform 1 0 18676 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_195
timestamp 1586364061
transform 1 0 19044 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_62_198
timestamp 1586364061
transform 1 0 19320 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_202
timestamp 1586364061
transform 1 0 19688 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_62_210
timestamp 1586364061
transform 1 0 20424 0 -1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _412_
timestamp 1586364061
transform 1 0 21436 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_62_215
timestamp 1586364061
transform 1 0 20884 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_220
timestamp 1586364061
transform 1 0 21344 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_230
timestamp 1586364061
transform 1 0 22264 0 -1 36448
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25760 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_247
timestamp 1586364061
transform 1 0 23828 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_251
timestamp 1586364061
transform 1 0 24196 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_8  FILLER_62_258
timestamp 1586364061
transform 1 0 24840 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_62_266
timestamp 1586364061
transform 1 0 25576 0 -1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_270
timestamp 1586364061
transform 1 0 25944 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_274
timestamp 1586364061
transform 1 0 26312 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  FILLER_62_285
timestamp 1586364061
transform 1 0 27324 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_62_290
timestamp 1586364061
transform 1 0 27784 0 -1 36448
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28336 0 -1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30176 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29624 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_305
timestamp 1586364061
transform 1 0 29164 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_309
timestamp 1586364061
transform 1 0 29532 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_312
timestamp 1586364061
transform 1 0 29808 0 -1 36448
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33028 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_325
timestamp 1586364061
transform 1 0 31004 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_62_333
timestamp 1586364061
transform 1 0 31740 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_337
timestamp 1586364061
transform 1 0 32108 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_341
timestamp 1586364061
transform 1 0 32476 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_345
timestamp 1586364061
transform 1 0 32844 0 -1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33580 0 -1 36448
box -38 -48 866 592
use scs8hd_decap_4  FILLER_62_349
timestamp 1586364061
transform 1 0 33212 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_362
timestamp 1586364061
transform 1 0 34408 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_62_374
timestamp 1586364061
transform 1 0 35512 0 -1 36448
box -38 -48 314 592
use scs8hd_nor2_4  _355_
timestamp 1586364061
transform 1 0 36064 0 -1 36448
box -38 -48 866 592
use scs8hd_buf_1  _386_
timestamp 1586364061
transform 1 0 37720 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__348__A
timestamp 1586364061
transform 1 0 35788 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37076 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_379
timestamp 1586364061
transform 1 0 35972 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_389
timestamp 1586364061
transform 1 0 36892 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_393
timestamp 1586364061
transform 1 0 37260 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_62_401
timestamp 1586364061
transform 1 0 37996 0 -1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _352_
timestamp 1586364061
transform 1 0 39100 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__354__B
timestamp 1586364061
transform 1 0 38548 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__386__A
timestamp 1586364061
transform 1 0 38180 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40572 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38916 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_405
timestamp 1586364061
transform 1 0 38364 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_409
timestamp 1586364061
transform 1 0 38732 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_62_422
timestamp 1586364061
transform 1 0 39928 0 -1 36448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_62_428
timestamp 1586364061
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41952 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_431
timestamp 1586364061
transform 1 0 40756 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_442
timestamp 1586364061
transform 1 0 41768 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_446
timestamp 1586364061
transform 1 0 42136 0 -1 36448
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43608 0 -1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44804 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44160 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44528 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_62_459
timestamp 1586364061
transform 1 0 43332 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_62_465
timestamp 1586364061
transform 1 0 43884 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_470
timestamp 1586364061
transform 1 0 44344 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_474
timestamp 1586364061
transform 1 0 44712 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46368 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_8  FILLER_62_484
timestamp 1586364061
transform 1 0 45632 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_12  FILLER_62_495
timestamp 1586364061
transform 1 0 46644 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_507
timestamp 1586364061
transform 1 0 47748 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 48852 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_515
timestamp 1586364061
transform 1 0 48484 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14536 0 1 36448
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_139
timestamp 1586364061
transform 1 0 13892 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_142
timestamp 1586364061
transform 1 0 14168 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_157
timestamp 1586364061
transform 1 0 15548 0 1 36448
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_163
timestamp 1586364061
transform 1 0 16100 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_174
timestamp 1586364061
transform 1 0 17112 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_179
timestamp 1586364061
transform 1 0 17572 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_184
timestamp 1586364061
transform 1 0 18032 0 1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_196
timestamp 1586364061
transform 1 0 19136 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_200
timestamp 1586364061
transform 1 0 19504 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_204
timestamp 1586364061
transform 1 0 19872 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_208
timestamp 1586364061
transform 1 0 20240 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__426__B
timestamp 1586364061
transform 1 0 23000 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_221
timestamp 1586364061
transform 1 0 21436 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_225
timestamp 1586364061
transform 1 0 21804 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_232
timestamp 1586364061
transform 1 0 22448 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_236
timestamp 1586364061
transform 1 0 22816 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_240
timestamp 1586364061
transform 1 0 23184 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__426__A
timestamp 1586364061
transform 1 0 23368 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 36448
box -38 -48 866 592
use scs8hd_decap_4  FILLER_63_258
timestamp 1586364061
transform 1 0 24840 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_254
timestamp 1586364061
transform 1 0 24472 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_265
timestamp 1586364061
transform 1 0 25484 0 1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_63_262
timestamp 1586364061
transform 1 0 25208 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25300 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25760 0 1 36448
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_277
timestamp 1586364061
transform 1 0 26588 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_281
timestamp 1586364061
transform 1 0 26956 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_294
timestamp 1586364061
transform 1 0 28152 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_302
timestamp 1586364061
transform 1 0 28888 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_298
timestamp 1586364061
transform 1 0 28520 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28704 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_306
timestamp 1586364061
transform 1 0 29256 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29624 0 1 36448
box -38 -48 866 592
use scs8hd_fill_2  FILLER_63_319
timestamp 1586364061
transform 1 0 30452 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30636 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_331
timestamp 1586364061
transform 1 0 31556 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_327
timestamp 1586364061
transform 1 0 31188 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_323
timestamp 1586364061
transform 1 0 30820 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__A
timestamp 1586364061
transform 1 0 31004 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_335
timestamp 1586364061
transform 1 0 31924 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32108 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32292 0 1 36448
box -38 -48 866 592
use scs8hd_decap_4  FILLER_63_348
timestamp 1586364061
transform 1 0 33120 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_354
timestamp 1586364061
transform 1 0 33672 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_358
timestamp 1586364061
transform 1 0 34040 0 1 36448
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_367
timestamp 1586364061
transform 1 0 34868 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__344__A
timestamp 1586364061
transform 1 0 34592 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use scs8hd_buf_1  _321_
timestamp 1586364061
transform 1 0 34960 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_375
timestamp 1586364061
transform 1 0 35604 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_371
timestamp 1586364061
transform 1 0 35236 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__321__A
timestamp 1586364061
transform 1 0 35420 0 1 36448
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 36800 0 1 36448
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 36616 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__344__B
timestamp 1586364061
transform 1 0 35788 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__397__A
timestamp 1586364061
transform 1 0 36248 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_379
timestamp 1586364061
transform 1 0 35972 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_384
timestamp 1586364061
transform 1 0 36432 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_399
timestamp 1586364061
transform 1 0 37812 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_403
timestamp 1586364061
transform 1 0 38180 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__354__A
timestamp 1586364061
transform 1 0 38364 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _354_
timestamp 1586364061
transform 1 0 38548 0 1 36448
box -38 -48 866 592
use scs8hd_decap_4  FILLER_63_420
timestamp 1586364061
transform 1 0 39744 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_416
timestamp 1586364061
transform 1 0 39376 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 39560 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_428
timestamp 1586364061
transform 1 0 40480 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_424
timestamp 1586364061
transform 1 0 40112 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42412 0 1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40848 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 40664 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42872 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41860 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_441
timestamp 1586364061
transform 1 0 41676 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_445
timestamp 1586364061
transform 1 0 42044 0 1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_63_452
timestamp 1586364061
transform 1 0 42688 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_456
timestamp 1586364061
transform 1 0 43056 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43424 0 1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44436 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43884 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44252 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45448 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43240 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_463
timestamp 1586364061
transform 1 0 43700 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_467
timestamp 1586364061
transform 1 0 44068 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_480
timestamp 1586364061
transform 1 0 45264 0 1 36448
box -38 -48 222 592
use scs8hd_conb_1  _654_
timestamp 1586364061
transform 1 0 46092 0 1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45816 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 46552 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_484
timestamp 1586364061
transform 1 0 45632 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_492
timestamp 1586364061
transform 1 0 46368 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_496
timestamp 1586364061
transform 1 0 46736 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_508
timestamp 1586364061
transform 1 0 47840 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 48852 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_68
timestamp 1586364061
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_80
timestamp 1586364061
transform 1 0 8464 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_93
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_105
timestamp 1586364061
transform 1 0 10764 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_117
timestamp 1586364061
transform 1 0 11868 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_129
timestamp 1586364061
transform 1 0 12972 0 -1 37536
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__432__B
timestamp 1586364061
transform 1 0 15456 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_141
timestamp 1586364061
transform 1 0 14076 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_64_154
timestamp 1586364061
transform 1 0 15272 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_158
timestamp 1586364061
transform 1 0 15640 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_170
timestamp 1586364061
transform 1 0 16744 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_174
timestamp 1586364061
transform 1 0 17112 0 -1 37536
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_189
timestamp 1586364061
transform 1 0 18492 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_193
timestamp 1586364061
transform 1 0 18860 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_8  FILLER_64_206
timestamp 1586364061
transform 1 0 20056 0 -1 37536
box -38 -48 774 592
use scs8hd_nor2_4  _426_
timestamp 1586364061
transform 1 0 22724 0 -1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__424__A
timestamp 1586364061
transform 1 0 21988 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_224
timestamp 1586364061
transform 1 0 21712 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_64_229
timestamp 1586364061
transform 1 0 22172 0 -1 37536
box -38 -48 590 592
use scs8hd_fill_2  FILLER_64_244
timestamp 1586364061
transform 1 0 23552 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_248
timestamp 1586364061
transform 1 0 23920 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23736 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_64_255
timestamp 1586364061
transform 1 0 24564 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_64_260
timestamp 1586364061
transform 1 0 25024 0 -1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_266
timestamp 1586364061
transform 1 0 25576 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25760 0 -1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28152 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__402__B
timestamp 1586364061
transform 1 0 27600 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_270
timestamp 1586364061
transform 1 0 25944 0 -1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_64_274
timestamp 1586364061
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_279
timestamp 1586364061
transform 1 0 26772 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_1  FILLER_64_287
timestamp 1586364061
transform 1 0 27508 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_290
timestamp 1586364061
transform 1 0 27784 0 -1 37536
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29900 0 -1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29164 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29532 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30452 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_303
timestamp 1586364061
transform 1 0 28980 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_307
timestamp 1586364061
transform 1 0 29348 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_311
timestamp 1586364061
transform 1 0 29716 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_316
timestamp 1586364061
transform 1 0 30176 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_321
timestamp 1586364061
transform 1 0 30636 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_328
timestamp 1586364061
transform 1 0 31280 0 -1 37536
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__400__B
timestamp 1586364061
transform 1 0 30820 0 -1 37536
box -38 -48 222 592
use scs8hd_buf_1  _384_
timestamp 1586364061
transform 1 0 31004 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_337
timestamp 1586364061
transform 1 0 32108 0 -1 37536
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use scs8hd_conb_1  _650_
timestamp 1586364061
transform 1 0 32200 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_345
timestamp 1586364061
transform 1 0 32844 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_341
timestamp 1586364061
transform 1 0 32476 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33028 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 -1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _344_
timestamp 1586364061
transform 1 0 35052 0 -1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33488 0 -1 37536
box -38 -48 866 592
use scs8hd_decap_3  FILLER_64_349
timestamp 1586364061
transform 1 0 33212 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_8  FILLER_64_361
timestamp 1586364061
transform 1 0 34316 0 -1 37536
box -38 -48 774 592
use scs8hd_buf_1  _397_
timestamp 1586364061
transform 1 0 36616 0 -1 37536
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37812 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37076 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_378
timestamp 1586364061
transform 1 0 35880 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_64_389
timestamp 1586364061
transform 1 0 36892 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_393
timestamp 1586364061
transform 1 0 37260 0 -1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_64_398
timestamp 1586364061
transform 1 0 37720 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_402
timestamp 1586364061
transform 1 0 38088 0 -1 37536
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 40572 0 -1 37536
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 38824 0 -1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__353__B
timestamp 1586364061
transform 1 0 38272 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_406
timestamp 1586364061
transform 1 0 38456 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_8  FILLER_64_421
timestamp 1586364061
transform 1 0 39836 0 -1 37536
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41768 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42320 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_440
timestamp 1586364061
transform 1 0 41584 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_444
timestamp 1586364061
transform 1 0 41952 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_8  FILLER_64_450
timestamp 1586364061
transform 1 0 42504 0 -1 37536
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44252 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43884 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_459
timestamp 1586364061
transform 1 0 43332 0 -1 37536
box -38 -48 590 592
use scs8hd_fill_2  FILLER_64_467
timestamp 1586364061
transform 1 0 44068 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_478
timestamp 1586364061
transform 1 0 45080 0 -1 37536
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45816 0 -1 37536
box -38 -48 866 592
use scs8hd_decap_12  FILLER_64_495
timestamp 1586364061
transform 1 0 46644 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_507
timestamp 1586364061
transform 1 0 47748 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 48852 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_515
timestamp 1586364061
transform 1 0 48484 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_74
timestamp 1586364061
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_86
timestamp 1586364061
transform 1 0 9016 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_98
timestamp 1586364061
transform 1 0 10120 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_110
timestamp 1586364061
transform 1 0 11224 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_123
timestamp 1586364061
transform 1 0 12420 0 1 37536
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__A
timestamp 1586364061
transform 1 0 15732 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_135
timestamp 1586364061
transform 1 0 13524 0 1 37536
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_65_147
timestamp 1586364061
transform 1 0 14628 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_153
timestamp 1586364061
transform 1 0 15180 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_157
timestamp 1586364061
transform 1 0 15548 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__435__B
timestamp 1586364061
transform 1 0 17756 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_170
timestamp 1586364061
transform 1 0 16744 0 1 37536
box -38 -48 406 592
use scs8hd_decap_4  FILLER_65_176
timestamp 1586364061
transform 1 0 17296 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_180
timestamp 1586364061
transform 1 0 17664 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_187
timestamp 1586364061
transform 1 0 18308 0 1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__435__A
timestamp 1586364061
transform 1 0 18860 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_191
timestamp 1586364061
transform 1 0 18676 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_195
timestamp 1586364061
transform 1 0 19044 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_209
timestamp 1586364061
transform 1 0 20332 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_213
timestamp 1586364061
transform 1 0 20700 0 1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _424_
timestamp 1586364061
transform 1 0 21988 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__424__B
timestamp 1586364061
transform 1 0 21804 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__437__A
timestamp 1586364061
transform 1 0 20884 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__437__B
timestamp 1586364061
transform 1 0 21252 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_217
timestamp 1586364061
transform 1 0 21068 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_221
timestamp 1586364061
transform 1 0 21436 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_236
timestamp 1586364061
transform 1 0 22816 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_240
timestamp 1586364061
transform 1 0 23184 0 1 37536
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 37536
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25576 0 1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_256
timestamp 1586364061
transform 1 0 24656 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_260
timestamp 1586364061
transform 1 0 25024 0 1 37536
box -38 -48 406 592
use scs8hd_nor2_4  _402_
timestamp 1586364061
transform 1 0 27600 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__402__A
timestamp 1586364061
transform 1 0 27416 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_275
timestamp 1586364061
transform 1 0 26404 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_279
timestamp 1586364061
transform 1 0 26772 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_283
timestamp 1586364061
transform 1 0 27140 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_301
timestamp 1586364061
transform 1 0 28796 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_297
timestamp 1586364061
transform 1 0 28428 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 37536
box -38 -48 866 592
use scs8hd_fill_2  FILLER_65_319
timestamp 1586364061
transform 1 0 30452 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_315
timestamp 1586364061
transform 1 0 30084 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__A
timestamp 1586364061
transform 1 0 30636 0 1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _400_
timestamp 1586364061
transform 1 0 30820 0 1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32568 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_332
timestamp 1586364061
transform 1 0 31648 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_336
timestamp 1586364061
transform 1 0 32016 0 1 37536
box -38 -48 130 592
use scs8hd_decap_3  FILLER_65_339
timestamp 1586364061
transform 1 0 32292 0 1 37536
box -38 -48 314 592
use scs8hd_decap_4  FILLER_65_359
timestamp 1586364061
transform 1 0 34132 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_355
timestamp 1586364061
transform 1 0 33764 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_351
timestamp 1586364061
transform 1 0 33396 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33580 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__322__A
timestamp 1586364061
transform 1 0 33948 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_371
timestamp 1586364061
transform 1 0 35236 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_367
timestamp 1586364061
transform 1 0 34868 0 1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_65_363
timestamp 1586364061
transform 1 0 34500 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__341__A
timestamp 1586364061
transform 1 0 34592 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__341__B
timestamp 1586364061
transform 1 0 35052 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35420 0 1 37536
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35604 0 1 37536
box -38 -48 1050 592
use scs8hd_nor2_4  _353_
timestamp 1586364061
transform 1 0 37996 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__353__A
timestamp 1586364061
transform 1 0 37812 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__A
timestamp 1586364061
transform 1 0 37444 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__370__A
timestamp 1586364061
transform 1 0 36800 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_386
timestamp 1586364061
transform 1 0 36616 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_390
timestamp 1586364061
transform 1 0 36984 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_394
timestamp 1586364061
transform 1 0 37352 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_397
timestamp 1586364061
transform 1 0 37628 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39560 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__B
timestamp 1586364061
transform 1 0 39008 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_410
timestamp 1586364061
transform 1 0 38824 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_414
timestamp 1586364061
transform 1 0 39192 0 1 37536
box -38 -48 406 592
use scs8hd_decap_4  FILLER_65_420
timestamp 1586364061
transform 1 0 39744 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_424
timestamp 1586364061
transform 1 0 40112 0 1 37536
box -38 -48 130 592
use scs8hd_decap_3  FILLER_65_428
timestamp 1586364061
transform 1 0 40480 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42320 0 1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40756 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42136 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_440
timestamp 1586364061
transform 1 0 41584 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_444
timestamp 1586364061
transform 1 0 41952 0 1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44068 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43884 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45080 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_457
timestamp 1586364061
transform 1 0 43148 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_463
timestamp 1586364061
transform 1 0 43700 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_476
timestamp 1586364061
transform 1 0 44896 0 1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_65_480
timestamp 1586364061
transform 1 0 45264 0 1 37536
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_492
timestamp 1586364061
transform 1 0 46368 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_496
timestamp 1586364061
transform 1 0 46736 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_508
timestamp 1586364061
transform 1 0 47840 0 1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 48852 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_80
timestamp 1586364061
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_93
timestamp 1586364061
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_105
timestamp 1586364061
transform 1 0 10764 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_86
timestamp 1586364061
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_98
timestamp 1586364061
transform 1 0 10120 0 1 38624
box -38 -48 1142 592
use scs8hd_nor2_4  _434_
timestamp 1586364061
transform 1 0 13156 0 1 38624
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__434__A
timestamp 1586364061
transform 1 0 12972 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__434__B
timestamp 1586364061
transform 1 0 13156 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_117
timestamp 1586364061
transform 1 0 11868 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_66_129
timestamp 1586364061
transform 1 0 12972 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_133
timestamp 1586364061
transform 1 0 13340 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_110
timestamp 1586364061
transform 1 0 11224 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_67_123
timestamp 1586364061
transform 1 0 12420 0 1 38624
box -38 -48 590 592
use scs8hd_decap_6  FILLER_67_140
timestamp 1586364061
transform 1 0 13984 0 1 38624
box -38 -48 590 592
use scs8hd_decap_3  FILLER_66_150
timestamp 1586364061
transform 1 0 14904 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  FILLER_66_145
timestamp 1586364061
transform 1 0 14444 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__431__B
timestamp 1586364061
transform 1 0 14720 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__431__A
timestamp 1586364061
transform 1 0 14536 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use scs8hd_nor2_4  _431_
timestamp 1586364061
transform 1 0 14720 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_161
timestamp 1586364061
transform 1 0 15916 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_157
timestamp 1586364061
transform 1 0 15548 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_154
timestamp 1586364061
transform 1 0 15272 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__433__A
timestamp 1586364061
transform 1 0 15732 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _432_
timestamp 1586364061
transform 1 0 15364 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_66_168
timestamp 1586364061
transform 1 0 16560 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_164
timestamp 1586364061
transform 1 0 16192 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__433__B
timestamp 1586364061
transform 1 0 16376 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _433_
timestamp 1586364061
transform 1 0 16284 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_179
timestamp 1586364061
transform 1 0 17572 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_174
timestamp 1586364061
transform 1 0 17112 0 1 38624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_66_177
timestamp 1586364061
transform 1 0 17388 0 -1 38624
box -38 -48 590 592
use scs8hd_fill_2  FILLER_66_172
timestamp 1586364061
transform 1 0 16928 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17112 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_184
timestamp 1586364061
transform 1 0 18032 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17940 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__430__B
timestamp 1586364061
transform 1 0 17756 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__430__A
timestamp 1586364061
transform 1 0 18216 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use scs8hd_nor2_4  _435_
timestamp 1586364061
transform 1 0 18124 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_197
timestamp 1586364061
transform 1 0 19228 0 1 38624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_66_194
timestamp 1586364061
transform 1 0 18952 0 -1 38624
box -38 -48 590 592
use scs8hd_nor2_4  _430_
timestamp 1586364061
transform 1 0 18400 0 1 38624
box -38 -48 866 592
use scs8hd_decap_6  FILLER_67_202
timestamp 1586364061
transform 1 0 19688 0 1 38624
box -38 -48 590 592
use scs8hd_decap_8  FILLER_66_206
timestamp 1586364061
transform 1 0 20056 0 -1 38624
box -38 -48 774 592
use scs8hd_fill_1  FILLER_66_202
timestamp 1586364061
transform 1 0 19688 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_211
timestamp 1586364061
transform 1 0 20516 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_67_208
timestamp 1586364061
transform 1 0 20240 0 1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__436__B
timestamp 1586364061
transform 1 0 20332 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__436__A
timestamp 1586364061
transform 1 0 20700 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_224
timestamp 1586364061
transform 1 0 21712 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_224
timestamp 1586364061
transform 1 0 21712 0 -1 38624
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21896 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _437_
timestamp 1586364061
transform 1 0 20884 0 -1 38624
box -38 -48 866 592
use scs8hd_nor2_4  _436_
timestamp 1586364061
transform 1 0 20884 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_239
timestamp 1586364061
transform 1 0 23092 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_235
timestamp 1586364061
transform 1 0 22724 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_228
timestamp 1586364061
transform 1 0 22080 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22816 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 38624
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23000 0 -1 38624
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23276 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_67_245
timestamp 1586364061
transform 1 0 23644 0 1 38624
box -38 -48 406 592
use scs8hd_fill_1  FILLER_67_243
timestamp 1586364061
transform 1 0 23460 0 1 38624
box -38 -48 130 592
use scs8hd_decap_8  FILLER_66_249
timestamp 1586364061
transform 1 0 24012 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__428__A
timestamp 1586364061
transform 1 0 24012 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_258
timestamp 1586364061
transform 1 0 24840 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_254
timestamp 1586364061
transform 1 0 24472 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_257
timestamp 1586364061
transform 1 0 24748 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 38624
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 25208 0 1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_66_267
timestamp 1586364061
transform 1 0 25668 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_67_273
timestamp 1586364061
transform 1 0 26220 0 1 38624
box -38 -48 406 592
use scs8hd_decap_4  FILLER_66_271
timestamp 1586364061
transform 1 0 26036 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__403__A
timestamp 1586364061
transform 1 0 26588 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_283
timestamp 1586364061
transform 1 0 27140 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_279
timestamp 1586364061
transform 1 0 26772 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_66_285
timestamp 1586364061
transform 1 0 27324 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__401__B
timestamp 1586364061
transform 1 0 27600 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__403__B
timestamp 1586364061
transform 1 0 26956 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__A
timestamp 1586364061
transform 1 0 27416 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _401_
timestamp 1586364061
transform 1 0 27600 0 1 38624
box -38 -48 866 592
use scs8hd_fill_1  FILLER_66_294
timestamp 1586364061
transform 1 0 28152 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_290
timestamp 1586364061
transform 1 0 27784 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28244 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_301
timestamp 1586364061
transform 1 0 28796 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_297
timestamp 1586364061
transform 1 0 28428 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_297
timestamp 1586364061
transform 1 0 28428 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 38624
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28520 0 -1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_67_315
timestamp 1586364061
transform 1 0 30084 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_317
timestamp 1586364061
transform 1 0 30268 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_309
timestamp 1586364061
transform 1 0 29532 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__398__A
timestamp 1586364061
transform 1 0 30268 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_319
timestamp 1586364061
transform 1 0 30452 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 30636 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_66_332
timestamp 1586364061
transform 1 0 31648 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_328
timestamp 1586364061
transform 1 0 31280 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31464 0 -1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 30820 0 1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_67_343
timestamp 1586364061
transform 1 0 32660 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_339
timestamp 1586364061
transform 1 0 32292 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_334
timestamp 1586364061
transform 1 0 31832 0 1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__399__B
timestamp 1586364061
transform 1 0 31832 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__332__A
timestamp 1586364061
transform 1 0 32476 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__332__B
timestamp 1586364061
transform 1 0 32844 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__399__A
timestamp 1586364061
transform 1 0 32108 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 38624
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_66_348
timestamp 1586364061
transform 1 0 33120 0 -1 38624
box -38 -48 590 592
use scs8hd_nor2_4  _332_
timestamp 1586364061
transform 1 0 33028 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_356
timestamp 1586364061
transform 1 0 33856 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_356
timestamp 1586364061
transform 1 0 33856 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 34040 0 1 38624
box -38 -48 222 592
use scs8hd_buf_1  _322_
timestamp 1586364061
transform 1 0 33948 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  FILLER_67_367
timestamp 1586364061
transform 1 0 34868 0 1 38624
box -38 -48 314 592
use scs8hd_decap_4  FILLER_67_360
timestamp 1586364061
transform 1 0 34224 0 1 38624
box -38 -48 406 592
use scs8hd_decap_8  FILLER_66_360
timestamp 1586364061
transform 1 0 34224 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use scs8hd_nor2_4  _341_
timestamp 1586364061
transform 1 0 34960 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_372
timestamp 1586364061
transform 1 0 35328 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35144 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 35512 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_387
timestamp 1586364061
transform 1 0 36708 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_385
timestamp 1586364061
transform 1 0 36524 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_381
timestamp 1586364061
transform 1 0 36156 0 -1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_66_377
timestamp 1586364061
transform 1 0 35788 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35972 0 -1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 35696 0 1 38624
box -38 -48 1050 592
use scs8hd_buf_1  _370_
timestamp 1586364061
transform 1 0 36616 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_398
timestamp 1586364061
transform 1 0 37720 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_391
timestamp 1586364061
transform 1 0 37076 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_389
timestamp 1586364061
transform 1 0 36892 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37260 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 38624
box -38 -48 314 592
use scs8hd_nor2_4  _378_
timestamp 1586364061
transform 1 0 37720 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_402
timestamp 1586364061
transform 1 0 38088 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__371__A
timestamp 1586364061
transform 1 0 37904 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_406
timestamp 1586364061
transform 1 0 38456 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_412
timestamp 1586364061
transform 1 0 39008 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_66_407
timestamp 1586364061
transform 1 0 38548 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__375__B
timestamp 1586364061
transform 1 0 38272 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__375__A
timestamp 1586364061
transform 1 0 38824 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 38640 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _375_
timestamp 1586364061
transform 1 0 38824 0 1 38624
box -38 -48 866 592
use scs8hd_decap_6  FILLER_67_419
timestamp 1586364061
transform 1 0 39652 0 1 38624
box -38 -48 590 592
use scs8hd_decap_8  FILLER_66_421
timestamp 1586364061
transform 1 0 39836 0 -1 38624
box -38 -48 774 592
use scs8hd_fill_2  FILLER_66_416
timestamp 1586364061
transform 1 0 39376 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39192 0 -1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39560 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_67_428
timestamp 1586364061
transform 1 0 40480 0 1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 -1 38624
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_436
timestamp 1586364061
transform 1 0 41216 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_432
timestamp 1586364061
transform 1 0 40848 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_436
timestamp 1586364061
transform 1 0 41216 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_432
timestamp 1586364061
transform 1 0 40848 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41400 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41400 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 41032 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_67_449
timestamp 1586364061
transform 1 0 42412 0 1 38624
box -38 -48 590 592
use scs8hd_decap_4  FILLER_67_443
timestamp 1586364061
transform 1 0 41860 0 1 38624
box -38 -48 406 592
use scs8hd_fill_1  FILLER_66_440
timestamp 1586364061
transform 1 0 41584 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41584 0 1 38624
box -38 -48 314 592
use scs8hd_decap_8  FILLER_66_450
timestamp 1586364061
transform 1 0 42504 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_467
timestamp 1586364061
transform 1 0 44068 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_461
timestamp 1586364061
transform 1 0 43516 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_457
timestamp 1586364061
transform 1 0 43148 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_66_459
timestamp 1586364061
transform 1 0 43332 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44252 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43884 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43792 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_67_471
timestamp 1586364061
transform 1 0 44436 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_474
timestamp 1586364061
transform 1 0 44712 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_67_483
timestamp 1586364061
transform 1 0 45540 0 1 38624
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_486
timestamp 1586364061
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_498
timestamp 1586364061
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_67_487
timestamp 1586364061
transform 1 0 45908 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_67_489
timestamp 1586364061
transform 1 0 46092 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_501
timestamp 1586364061
transform 1 0 47196 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 48852 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 48852 0 1 38624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_66_510
timestamp 1586364061
transform 1 0 48024 0 -1 38624
box -38 -48 590 592
use scs8hd_decap_3  FILLER_67_513
timestamp 1586364061
transform 1 0 48300 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_93
timestamp 1586364061
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_105
timestamp 1586364061
transform 1 0 10764 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_117
timestamp 1586364061
transform 1 0 11868 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_129
timestamp 1586364061
transform 1 0 12972 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_141
timestamp 1586364061
transform 1 0 14076 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_68_154
timestamp 1586364061
transform 1 0 15272 0 -1 39712
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 39712
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_68_162
timestamp 1586364061
transform 1 0 16008 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_175
timestamp 1586364061
transform 1 0 17204 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_68_192
timestamp 1586364061
transform 1 0 18768 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_68_197
timestamp 1586364061
transform 1 0 19228 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_8  FILLER_68_203
timestamp 1586364061
transform 1 0 19780 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_3  FILLER_68_211
timestamp 1586364061
transform 1 0 20516 0 -1 39712
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 39712
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23184 0 -1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_215
timestamp 1586364061
transform 1 0 20884 0 -1 39712
box -38 -48 590 592
use scs8hd_fill_2  FILLER_68_232
timestamp 1586364061
transform 1 0 22448 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_236
timestamp 1586364061
transform 1 0 22816 0 -1 39712
box -38 -48 406 592
use scs8hd_buf_1  _428_
timestamp 1586364061
transform 1 0 24196 0 -1 39712
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_243
timestamp 1586364061
transform 1 0 23460 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_4  FILLER_68_254
timestamp 1586364061
transform 1 0 24472 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_68_260
timestamp 1586364061
transform 1 0 25024 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_265
timestamp 1586364061
transform 1 0 25484 0 -1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _403_
timestamp 1586364061
transform 1 0 26588 0 -1 39712
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28244 0 -1 39712
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__390__B
timestamp 1586364061
transform 1 0 27600 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_269
timestamp 1586364061
transform 1 0 25852 0 -1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_68_276
timestamp 1586364061
transform 1 0 26496 0 -1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_68_286
timestamp 1586364061
transform 1 0 27416 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_290
timestamp 1586364061
transform 1 0 27784 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_68_294
timestamp 1586364061
transform 1 0 28152 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__394__B
timestamp 1586364061
transform 1 0 30452 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_306
timestamp 1586364061
transform 1 0 29256 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_310
timestamp 1586364061
transform 1 0 29624 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_1  FILLER_68_318
timestamp 1586364061
transform 1 0 30360 0 -1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_68_321
timestamp 1586364061
transform 1 0 30636 0 -1 39712
box -38 -48 222 592
use scs8hd_buf_1  _398_
timestamp 1586364061
transform 1 0 31004 0 -1 39712
box -38 -48 314 592
use scs8hd_nor2_4  _399_
timestamp 1586364061
transform 1 0 32108 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__395__A
timestamp 1586364061
transform 1 0 30820 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_328
timestamp 1586364061
transform 1 0 31280 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_3  FILLER_68_346
timestamp 1586364061
transform 1 0 32936 0 -1 39712
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 39712
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__329__A
timestamp 1586364061
transform 1 0 33212 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_68_351
timestamp 1586364061
transform 1 0 33396 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_8  FILLER_68_365
timestamp 1586364061
transform 1 0 34684 0 -1 39712
box -38 -48 774 592
use scs8hd_buf_1  _371_
timestamp 1586364061
transform 1 0 37720 0 -1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36800 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_382
timestamp 1586364061
transform 1 0 36248 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_386
timestamp 1586364061
transform 1 0 36616 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_390
timestamp 1586364061
transform 1 0 36984 0 -1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_68_396
timestamp 1586364061
transform 1 0 37536 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_8  FILLER_68_401
timestamp 1586364061
transform 1 0 37996 0 -1 39712
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 38732 0 -1 39712
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 40480 0 -1 39712
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_68_420
timestamp 1586364061
transform 1 0 39744 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41676 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_439
timestamp 1586364061
transform 1 0 41492 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_443
timestamp 1586364061
transform 1 0 41860 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_68_450
timestamp 1586364061
transform 1 0 42504 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_454
timestamp 1586364061
transform 1 0 42872 0 -1 39712
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_468
timestamp 1586364061
transform 1 0 44160 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_480
timestamp 1586364061
transform 1 0 45264 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_492
timestamp 1586364061
transform 1 0 46368 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_504
timestamp 1586364061
transform 1 0 47472 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 48852 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_86
timestamp 1586364061
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_98
timestamp 1586364061
transform 1 0 10120 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_110
timestamp 1586364061
transform 1 0 11224 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_123
timestamp 1586364061
transform 1 0 12420 0 1 39712
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_135
timestamp 1586364061
transform 1 0 13524 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_69_147
timestamp 1586364061
transform 1 0 14628 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_151
timestamp 1586364061
transform 1 0 14996 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_154
timestamp 1586364061
transform 1 0 15272 0 1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_69_158
timestamp 1586364061
transform 1 0 15640 0 1 39712
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16100 0 1 39712
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_174
timestamp 1586364061
transform 1 0 17112 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_178
timestamp 1586364061
transform 1 0 17480 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_182
timestamp 1586364061
transform 1 0 17848 0 1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_69_184
timestamp 1586364061
transform 1 0 18032 0 1 39712
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 19044 0 1 39712
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__429__A
timestamp 1586364061
transform 1 0 18492 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_188
timestamp 1586364061
transform 1 0 18400 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_191
timestamp 1586364061
transform 1 0 18676 0 1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_69_206
timestamp 1586364061
transform 1 0 20056 0 1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_69_214
timestamp 1586364061
transform 1 0 20792 0 1 39712
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20976 0 1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_219
timestamp 1586364061
transform 1 0 21252 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_223
timestamp 1586364061
transform 1 0 21620 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_236
timestamp 1586364061
transform 1 0 22816 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_240
timestamp 1586364061
transform 1 0 23184 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use scs8hd_buf_1  _410_
timestamp 1586364061
transform 1 0 23644 0 1 39712
box -38 -48 314 592
use scs8hd_fill_2  FILLER_69_248
timestamp 1586364061
transform 1 0 23920 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_252
timestamp 1586364061
transform 1 0 24288 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_256
timestamp 1586364061
transform 1 0 24656 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__410__A
timestamp 1586364061
transform 1 0 24472 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_260
timestamp 1586364061
transform 1 0 25024 0 1 39712
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 39712
box -38 -48 314 592
use scs8hd_fill_2  FILLER_69_264
timestamp 1586364061
transform 1 0 25392 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_268
timestamp 1586364061
transform 1 0 25760 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25576 0 1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _390_
timestamp 1586364061
transform 1 0 27508 0 1 39712
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__390__A
timestamp 1586364061
transform 1 0 27324 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__A
timestamp 1586364061
transform 1 0 26956 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__B
timestamp 1586364061
transform 1 0 26312 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25944 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_272
timestamp 1586364061
transform 1 0 26128 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_279
timestamp 1586364061
transform 1 0 26772 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_283
timestamp 1586364061
transform 1 0 27140 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_304
timestamp 1586364061
transform 1 0 29072 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_300
timestamp 1586364061
transform 1 0 28704 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_296
timestamp 1586364061
transform 1 0 28336 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28888 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28520 0 1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_69_306
timestamp 1586364061
transform 1 0 29256 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_321
timestamp 1586364061
transform 1 0 30636 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_317
timestamp 1586364061
transform 1 0 30268 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_314
timestamp 1586364061
transform 1 0 29992 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__395__B
timestamp 1586364061
transform 1 0 30084 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__A
timestamp 1586364061
transform 1 0 30452 0 1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _395_
timestamp 1586364061
transform 1 0 30820 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__335__B
timestamp 1586364061
transform 1 0 32108 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__329__B
timestamp 1586364061
transform 1 0 33028 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__A
timestamp 1586364061
transform 1 0 32476 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_332
timestamp 1586364061
transform 1 0 31648 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_336
timestamp 1586364061
transform 1 0 32016 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_339
timestamp 1586364061
transform 1 0 32292 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_343
timestamp 1586364061
transform 1 0 32660 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_358
timestamp 1586364061
transform 1 0 34040 0 1 39712
box -38 -48 222 592
use scs8hd_nor2_4  _329_
timestamp 1586364061
transform 1 0 33212 0 1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_69_367
timestamp 1586364061
transform 1 0 34868 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_362
timestamp 1586364061
transform 1 0 34408 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34592 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_375
timestamp 1586364061
transform 1 0 35604 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_371
timestamp 1586364061
transform 1 0 35236 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 35052 0 1 39712
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35328 0 1 39712
box -38 -48 314 592
use scs8hd_nor2_4  _379_
timestamp 1586364061
transform 1 0 37904 0 1 39712
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36340 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35788 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36156 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__A
timestamp 1586364061
transform 1 0 37720 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_379
timestamp 1586364061
transform 1 0 35972 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_392
timestamp 1586364061
transform 1 0 37168 0 1 39712
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 40480 0 1 39712
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__A
timestamp 1586364061
transform 1 0 39100 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__B
timestamp 1586364061
transform 1 0 39468 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_409
timestamp 1586364061
transform 1 0 38732 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_415
timestamp 1586364061
transform 1 0 39284 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_419
timestamp 1586364061
transform 1 0 39652 0 1 39712
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42688 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42504 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_439
timestamp 1586364061
transform 1 0 41492 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_443
timestamp 1586364061
transform 1 0 41860 0 1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_69_447
timestamp 1586364061
transform 1 0 42228 0 1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_461
timestamp 1586364061
transform 1 0 43516 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_465
timestamp 1586364061
transform 1 0 43884 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_477
timestamp 1586364061
transform 1 0 44988 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_69_485
timestamp 1586364061
transform 1 0 45724 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_489
timestamp 1586364061
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_501
timestamp 1586364061
transform 1 0 47196 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 48852 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_69_513
timestamp 1586364061
transform 1 0 48300 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_93
timestamp 1586364061
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_105
timestamp 1586364061
transform 1 0 10764 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_117
timestamp 1586364061
transform 1 0 11868 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_129
timestamp 1586364061
transform 1 0 12972 0 -1 40800
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 40800
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_141
timestamp 1586364061
transform 1 0 14076 0 -1 40800
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_70_154
timestamp 1586364061
transform 1 0 15272 0 -1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_167
timestamp 1586364061
transform 1 0 16468 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_171
timestamp 1586364061
transform 1 0 16836 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_184
timestamp 1586364061
transform 1 0 18032 0 -1 40800
box -38 -48 774 592
use scs8hd_buf_1  _429_
timestamp 1586364061
transform 1 0 18952 0 -1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_192
timestamp 1586364061
transform 1 0 18768 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_70_197
timestamp 1586364061
transform 1 0 19228 0 -1 40800
box -38 -48 590 592
use scs8hd_decap_8  FILLER_70_205
timestamp 1586364061
transform 1 0 19964 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_1  FILLER_70_213
timestamp 1586364061
transform 1 0 20700 0 -1 40800
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22172 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_70_215
timestamp 1586364061
transform 1 0 20884 0 -1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_70_221
timestamp 1586364061
transform 1 0 21436 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_225
timestamp 1586364061
transform 1 0 21804 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_238
timestamp 1586364061
transform 1 0 23000 0 -1 40800
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24656 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_70_249
timestamp 1586364061
transform 1 0 24012 0 -1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_70_254
timestamp 1586364061
transform 1 0 24472 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_267
timestamp 1586364061
transform 1 0 25668 0 -1 40800
box -38 -48 774 592
use scs8hd_nor2_4  _391_
timestamp 1586364061
transform 1 0 26680 0 -1 40800
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28244 0 -1 40800
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27784 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_276
timestamp 1586364061
transform 1 0 26496 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_70_287
timestamp 1586364061
transform 1 0 27508 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_3  FILLER_70_292
timestamp 1586364061
transform 1 0 27968 0 -1 40800
box -38 -48 314 592
use scs8hd_nor2_4  _394_
timestamp 1586364061
transform 1 0 30452 0 -1 40800
box -38 -48 866 592
use scs8hd_decap_12  FILLER_70_306
timestamp 1586364061
transform 1 0 29256 0 -1 40800
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_70_318
timestamp 1586364061
transform 1 0 30360 0 -1 40800
box -38 -48 130 592
use scs8hd_nor2_4  _335_
timestamp 1586364061
transform 1 0 32108 0 -1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_328
timestamp 1586364061
transform 1 0 31280 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_8  FILLER_70_346
timestamp 1586364061
transform 1 0 32936 0 -1 40800
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 34684 0 -1 40800
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_8  FILLER_70_357
timestamp 1586364061
transform 1 0 33948 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_4  FILLER_70_380
timestamp 1586364061
transform 1 0 36064 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_70_376
timestamp 1586364061
transform 1 0 35696 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_70_387
timestamp 1586364061
transform 1 0 36708 0 -1 40800
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37260 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_402
timestamp 1586364061
transform 1 0 38088 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_70_398
timestamp 1586364061
transform 1 0 37720 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_395
timestamp 1586364061
transform 1 0 37444 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__B
timestamp 1586364061
transform 1 0 37904 0 -1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use scs8hd_nor2_4  _374_
timestamp 1586364061
transform 1 0 39100 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__376__B
timestamp 1586364061
transform 1 0 38824 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_70_412
timestamp 1586364061
transform 1 0 39008 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_6  FILLER_70_422
timestamp 1586364061
transform 1 0 39928 0 -1 40800
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41492 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_430
timestamp 1586364061
transform 1 0 40664 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_1  FILLER_70_438
timestamp 1586364061
transform 1 0 41400 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_450
timestamp 1586364061
transform 1 0 42504 0 -1 40800
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_462
timestamp 1586364061
transform 1 0 43608 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_474
timestamp 1586364061
transform 1 0 44712 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_486
timestamp 1586364061
transform 1 0 45816 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_498
timestamp 1586364061
transform 1 0 46920 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 48852 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_70_510
timestamp 1586364061
transform 1 0 48024 0 -1 40800
box -38 -48 590 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_86
timestamp 1586364061
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_98
timestamp 1586364061
transform 1 0 10120 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_110
timestamp 1586364061
transform 1 0 11224 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_123
timestamp 1586364061
transform 1 0 12420 0 1 40800
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_135
timestamp 1586364061
transform 1 0 13524 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_147
timestamp 1586364061
transform 1 0 14628 0 1 40800
box -38 -48 774 592
use scs8hd_fill_1  FILLER_71_155
timestamp 1586364061
transform 1 0 15364 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_158
timestamp 1586364061
transform 1 0 15640 0 1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_162
timestamp 1586364061
transform 1 0 16008 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_175
timestamp 1586364061
transform 1 0 17204 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_179
timestamp 1586364061
transform 1 0 17572 0 1 40800
box -38 -48 406 592
use scs8hd_decap_6  FILLER_71_184
timestamp 1586364061
transform 1 0 18032 0 1 40800
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_192
timestamp 1586364061
transform 1 0 18768 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_196
timestamp 1586364061
transform 1 0 19136 0 1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_71_200
timestamp 1586364061
transform 1 0 19504 0 1 40800
box -38 -48 130 592
use scs8hd_decap_3  FILLER_71_212
timestamp 1586364061
transform 1 0 20608 0 1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_217
timestamp 1586364061
transform 1 0 21068 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_221
timestamp 1586364061
transform 1 0 21436 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_236
timestamp 1586364061
transform 1 0 22816 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_240
timestamp 1586364061
transform 1 0 23184 0 1 40800
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 24840 0 1 40800
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_245
timestamp 1586364061
transform 1 0 23644 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_250
timestamp 1586364061
transform 1 0 24104 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_254
timestamp 1586364061
transform 1 0 24472 0 1 40800
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 27416 0 1 40800
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_269
timestamp 1586364061
transform 1 0 25852 0 1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_71_273
timestamp 1586364061
transform 1 0 26220 0 1 40800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_71_278
timestamp 1586364061
transform 1 0 26680 0 1 40800
box -38 -48 590 592
use scs8hd_fill_2  FILLER_71_306
timestamp 1586364061
transform 1 0 29256 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_301
timestamp 1586364061
transform 1 0 28796 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_297
timestamp 1586364061
transform 1 0 28428 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_314
timestamp 1586364061
transform 1 0 29992 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_310
timestamp 1586364061
transform 1 0 29624 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29808 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 30176 0 1 40800
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 30360 0 1 40800
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32660 0 1 40800
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32476 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__387__A
timestamp 1586364061
transform 1 0 31556 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_329
timestamp 1586364061
transform 1 0 31372 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_333
timestamp 1586364061
transform 1 0 31740 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_339
timestamp 1586364061
transform 1 0 32292 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_354
timestamp 1586364061
transform 1 0 33672 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33856 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_358
timestamp 1586364061
transform 1 0 34040 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_362
timestamp 1586364061
transform 1 0 34408 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_367
timestamp 1586364061
transform 1 0 34868 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_371
timestamp 1586364061
transform 1 0 35236 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35052 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35420 0 1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_71_375
timestamp 1586364061
transform 1 0 35604 0 1 40800
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37260 0 1 40800
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35696 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__373__B
timestamp 1586364061
transform 1 0 37076 0 1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_71_385
timestamp 1586364061
transform 1 0 36524 0 1 40800
box -38 -48 590 592
use scs8hd_fill_2  FILLER_71_402
timestamp 1586364061
transform 1 0 38088 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_406
timestamp 1586364061
transform 1 0 38456 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__376__A
timestamp 1586364061
transform 1 0 38640 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__373__A
timestamp 1586364061
transform 1 0 38272 0 1 40800
box -38 -48 222 592
use scs8hd_nor2_4  _376_
timestamp 1586364061
transform 1 0 38824 0 1 40800
box -38 -48 866 592
use scs8hd_fill_2  FILLER_71_419
timestamp 1586364061
transform 1 0 39652 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_71_428
timestamp 1586364061
transform 1 0 40480 0 1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_71_423
timestamp 1586364061
transform 1 0 40020 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 40800
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40940 0 1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41952 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41400 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_436
timestamp 1586364061
transform 1 0 41216 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_440
timestamp 1586364061
transform 1 0 41584 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_453
timestamp 1586364061
transform 1 0 42780 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_457
timestamp 1586364061
transform 1 0 43148 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_461
timestamp 1586364061
transform 1 0 43516 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_473
timestamp 1586364061
transform 1 0 44620 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use scs8hd_decap_3  FILLER_71_485
timestamp 1586364061
transform 1 0 45724 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_489
timestamp 1586364061
transform 1 0 46092 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_501
timestamp 1586364061
transform 1 0 47196 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 48852 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  FILLER_71_513
timestamp 1586364061
transform 1 0 48300 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_93
timestamp 1586364061
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_105
timestamp 1586364061
transform 1 0 10764 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_86
timestamp 1586364061
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_98
timestamp 1586364061
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_117
timestamp 1586364061
transform 1 0 11868 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_129
timestamp 1586364061
transform 1 0 12972 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_110
timestamp 1586364061
transform 1 0 11224 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_123
timestamp 1586364061
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_73_143
timestamp 1586364061
transform 1 0 14260 0 1 41888
box -38 -48 314 592
use scs8hd_decap_8  FILLER_73_135
timestamp 1586364061
transform 1 0 13524 0 1 41888
box -38 -48 774 592
use scs8hd_decap_12  FILLER_72_141
timestamp 1586364061
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_153
timestamp 1586364061
transform 1 0 15180 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_149
timestamp 1586364061
transform 1 0 14812 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_159
timestamp 1586364061
transform 1 0 15732 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_154
timestamp 1586364061
transform 1 0 15272 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 41888
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15548 0 1 41888
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_172
timestamp 1586364061
transform 1 0 16928 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_168
timestamp 1586364061
transform 1 0 16560 0 1 41888
box -38 -48 222 592
use scs8hd_decap_4  FILLER_72_163
timestamp 1586364061
transform 1 0 16100 0 -1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 41888
box -38 -48 866 592
use scs8hd_decap_3  FILLER_73_184
timestamp 1586364061
transform 1 0 18032 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_73_182
timestamp 1586364061
transform 1 0 17848 0 1 41888
box -38 -48 130 592
use scs8hd_decap_6  FILLER_73_176
timestamp 1586364061
transform 1 0 17296 0 1 41888
box -38 -48 590 592
use scs8hd_decap_12  FILLER_72_176
timestamp 1586364061
transform 1 0 17296 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use scs8hd_conb_1  _648_
timestamp 1586364061
transform 1 0 18308 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_194
timestamp 1586364061
transform 1 0 18952 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_190
timestamp 1586364061
transform 1 0 18584 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_188
timestamp 1586364061
transform 1 0 18400 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 41888
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 41888
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_73_211
timestamp 1586364061
transform 1 0 20516 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_207
timestamp 1586364061
transform 1 0 20148 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_205
timestamp 1586364061
transform 1 0 19964 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_72_201
timestamp 1586364061
transform 1 0 19596 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_213
timestamp 1586364061
transform 1 0 20700 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_73_222
timestamp 1586364061
transform 1 0 21528 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_218
timestamp 1586364061
transform 1 0 21160 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_226
timestamp 1586364061
transform 1 0 21896 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 41888
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 41888
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_73_235
timestamp 1586364061
transform 1 0 22724 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_230
timestamp 1586364061
transform 1 0 22264 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_239
timestamp 1586364061
transform 1 0 23092 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_252
timestamp 1586364061
transform 1 0 24288 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_245
timestamp 1586364061
transform 1 0 23644 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_73_243
timestamp 1586364061
transform 1 0 23460 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_243
timestamp 1586364061
transform 1 0 23460 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_256
timestamp 1586364061
transform 1 0 24656 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_267
timestamp 1586364061
transform 1 0 25668 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_255
timestamp 1586364061
transform 1 0 24564 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 41888
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_273
timestamp 1586364061
transform 1 0 26220 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_269
timestamp 1586364061
transform 1 0 25852 0 1 41888
box -38 -48 222 592
use scs8hd_decap_4  FILLER_72_271
timestamp 1586364061
transform 1 0 26036 0 -1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__B
timestamp 1586364061
transform 1 0 26404 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_286
timestamp 1586364061
transform 1 0 27416 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_288
timestamp 1586364061
transform 1 0 27600 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_3  FILLER_72_283
timestamp 1586364061
transform 1 0 27140 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_72_279
timestamp 1586364061
transform 1 0 26772 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27416 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26956 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__A
timestamp 1586364061
transform 1 0 27600 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_290
timestamp 1586364061
transform 1 0 27784 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27784 0 -1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_301
timestamp 1586364061
transform 1 0 28796 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_297
timestamp 1586364061
transform 1 0 28428 0 1 41888
box -38 -48 222 592
use scs8hd_decap_4  FILLER_72_303
timestamp 1586364061
transform 1 0 28980 0 -1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_299
timestamp 1586364061
transform 1 0 28612 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28796 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_73_313
timestamp 1586364061
transform 1 0 29900 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_73_310
timestamp 1586364061
transform 1 0 29624 0 1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_73_306
timestamp 1586364061
transform 1 0 29256 0 1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__389__A
timestamp 1586364061
transform 1 0 29716 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29348 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_72_320
timestamp 1586364061
transform 1 0 30544 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_316
timestamp 1586364061
transform 1 0 30176 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30728 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__389__B
timestamp 1586364061
transform 1 0 30360 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 30084 0 1 41888
box -38 -48 222 592
use scs8hd_nor2_4  _389_
timestamp 1586364061
transform 1 0 30268 0 1 41888
box -38 -48 866 592
use scs8hd_decap_4  FILLER_73_326
timestamp 1586364061
transform 1 0 31096 0 1 41888
box -38 -48 406 592
use scs8hd_decap_8  FILLER_72_327
timestamp 1586364061
transform 1 0 31188 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__326__A
timestamp 1586364061
transform 1 0 31464 0 1 41888
box -38 -48 222 592
use scs8hd_buf_1  _387_
timestamp 1586364061
transform 1 0 30912 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_332
timestamp 1586364061
transform 1 0 31648 0 1 41888
box -38 -48 222 592
use scs8hd_decap_6  FILLER_72_337
timestamp 1586364061
transform 1 0 32108 0 -1 41888
box -38 -48 590 592
use scs8hd_fill_1  FILLER_72_335
timestamp 1586364061
transform 1 0 31924 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__326__B
timestamp 1586364061
transform 1 0 31832 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use scs8hd_nor2_4  _326_
timestamp 1586364061
transform 1 0 32016 0 1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_345
timestamp 1586364061
transform 1 0 32844 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_348
timestamp 1586364061
transform 1 0 33120 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 33028 0 1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32844 0 -1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_73_356
timestamp 1586364061
transform 1 0 33856 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_349
timestamp 1586364061
transform 1 0 33212 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33396 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34040 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 1 41888
box -38 -48 314 592
use scs8hd_decap_4  FILLER_73_360
timestamp 1586364061
transform 1 0 34224 0 1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_365
timestamp 1586364061
transform 1 0 34684 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_72_369
timestamp 1586364061
transform 1 0 35052 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_380
timestamp 1586364061
transform 1 0 36064 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_376
timestamp 1586364061
transform 1 0 35696 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_382
timestamp 1586364061
transform 1 0 36248 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 41888
box -38 -48 866 592
use scs8hd_decap_4  FILLER_73_393
timestamp 1586364061
transform 1 0 37260 0 1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_395
timestamp 1586364061
transform 1 0 37444 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_392
timestamp 1586364061
transform 1 0 37168 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_6  FILLER_72_386
timestamp 1586364061
transform 1 0 36616 0 -1 41888
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37260 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_400
timestamp 1586364061
transform 1 0 37904 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_73_397
timestamp 1586364061
transform 1 0 37628 0 1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_72_398
timestamp 1586364061
transform 1 0 37720 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use scs8hd_nor2_4  _373_
timestamp 1586364061
transform 1 0 37904 0 -1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_404
timestamp 1586364061
transform 1 0 38272 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_413
timestamp 1586364061
transform 1 0 39100 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_409
timestamp 1586364061
transform 1 0 38732 0 -1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39192 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 41888
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 38640 0 1 41888
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_73_423
timestamp 1586364061
transform 1 0 40020 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_419
timestamp 1586364061
transform 1 0 39652 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_420
timestamp 1586364061
transform 1 0 39744 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_416
timestamp 1586364061
transform 1 0 39376 0 -1 41888
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 41888
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 39836 0 -1 41888
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_73_428
timestamp 1586364061
transform 1 0 40480 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_73_439
timestamp 1586364061
transform 1 0 41492 0 1 41888
box -38 -48 222 592
use scs8hd_decap_4  FILLER_72_436
timestamp 1586364061
transform 1 0 41216 0 -1 41888
box -38 -48 406 592
use scs8hd_fill_2  FILLER_72_432
timestamp 1586364061
transform 1 0 40848 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41032 0 -1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 1 41888
box -38 -48 866 592
use scs8hd_fill_2  FILLER_73_443
timestamp 1586364061
transform 1 0 41860 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_440
timestamp 1586364061
transform 1 0 41584 0 -1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 41888
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 41888
box -38 -48 866 592
use scs8hd_decap_3  FILLER_73_456
timestamp 1586364061
transform 1 0 43056 0 1 41888
box -38 -48 314 592
use scs8hd_decap_8  FILLER_72_450
timestamp 1586364061
transform 1 0 42504 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_3  FILLER_73_461
timestamp 1586364061
transform 1 0 43516 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_72_466
timestamp 1586364061
transform 1 0 43976 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_462
timestamp 1586364061
transform 1 0 43608 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44160 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_8  FILLER_73_477
timestamp 1586364061
transform 1 0 44988 0 1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_73_473
timestamp 1586364061
transform 1 0 44620 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_72_470
timestamp 1586364061
transform 1 0 44344 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44804 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_72_482
timestamp 1586364061
transform 1 0 45448 0 -1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_494
timestamp 1586364061
transform 1 0 46552 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_72_506
timestamp 1586364061
transform 1 0 47656 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_3  FILLER_73_485
timestamp 1586364061
transform 1 0 45724 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_73_489
timestamp 1586364061
transform 1 0 46092 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_501
timestamp 1586364061
transform 1 0 47196 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 48852 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 48852 0 1 41888
box -38 -48 314 592
use scs8hd_fill_2  FILLER_72_514
timestamp 1586364061
transform 1 0 48392 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_3  FILLER_73_513
timestamp 1586364061
transform 1 0 48300 0 1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_93
timestamp 1586364061
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_105
timestamp 1586364061
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_117
timestamp 1586364061
transform 1 0 11868 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_129
timestamp 1586364061
transform 1 0 12972 0 -1 42976
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 42976
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_74_141
timestamp 1586364061
transform 1 0 14076 0 -1 42976
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_74_154
timestamp 1586364061
transform 1 0 15272 0 -1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_74_158
timestamp 1586364061
transform 1 0 15640 0 -1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 42976
box -38 -48 866 592
use scs8hd_decap_4  FILLER_74_162
timestamp 1586364061
transform 1 0 16008 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_8  FILLER_74_175
timestamp 1586364061
transform 1 0 17204 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_1  FILLER_74_183
timestamp 1586364061
transform 1 0 17940 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_6  FILLER_74_187
timestamp 1586364061
transform 1 0 18308 0 -1 42976
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_74_204
timestamp 1586364061
transform 1 0 19872 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_74_212
timestamp 1586364061
transform 1 0 20608 0 -1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 -1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_6  FILLER_74_218
timestamp 1586364061
transform 1 0 21160 0 -1 42976
box -38 -48 590 592
use scs8hd_decap_12  FILLER_74_235
timestamp 1586364061
transform 1 0 22724 0 -1 42976
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_6  FILLER_74_250
timestamp 1586364061
transform 1 0 24104 0 -1 42976
box -38 -48 590 592
use scs8hd_decap_8  FILLER_74_267
timestamp 1586364061
transform 1 0 25668 0 -1 42976
box -38 -48 774 592
use scs8hd_nor2_4  _392_
timestamp 1586364061
transform 1 0 26772 0 -1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_3  FILLER_74_276
timestamp 1586364061
transform 1 0 26496 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_8  FILLER_74_288
timestamp 1586364061
transform 1 0 27600 0 -1 42976
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 30176 0 -1 42976
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28612 0 -1 42976
box -38 -48 866 592
use scs8hd_decap_3  FILLER_74_296
timestamp 1586364061
transform 1 0 28336 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_8  FILLER_74_308
timestamp 1586364061
transform 1 0 29440 0 -1 42976
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 32660 0 -1 42976
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__323__B
timestamp 1586364061
transform 1 0 32292 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_74_327
timestamp 1586364061
transform 1 0 31188 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_1  FILLER_74_335
timestamp 1586364061
transform 1 0 31924 0 -1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_74_337
timestamp 1586364061
transform 1 0 32108 0 -1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_74_341
timestamp 1586364061
transform 1 0 32476 0 -1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34592 0 -1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35604 0 -1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34408 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_74_354
timestamp 1586364061
transform 1 0 33672 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_74_373
timestamp 1586364061
transform 1 0 35420 0 -1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 42976
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36248 0 -1 42976
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36708 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_4  FILLER_74_377
timestamp 1586364061
transform 1 0 35788 0 -1 42976
box -38 -48 406 592
use scs8hd_fill_1  FILLER_74_381
timestamp 1586364061
transform 1 0 36156 0 -1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_74_385
timestamp 1586364061
transform 1 0 36524 0 -1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_74_389
timestamp 1586364061
transform 1 0 36892 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_4  FILLER_74_401
timestamp 1586364061
transform 1 0 37996 0 -1 42976
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 39192 0 -1 42976
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__377__A
timestamp 1586364061
transform 1 0 38456 0 -1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_74_405
timestamp 1586364061
transform 1 0 38364 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_6  FILLER_74_408
timestamp 1586364061
transform 1 0 38640 0 -1 42976
box -38 -48 590 592
use scs8hd_decap_4  FILLER_74_425
timestamp 1586364061
transform 1 0 40204 0 -1 42976
box -38 -48 406 592
use scs8hd_fill_1  FILLER_74_429
timestamp 1586364061
transform 1 0 40572 0 -1 42976
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 -1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42228 0 -1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40664 0 -1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_74_432
timestamp 1586364061
transform 1 0 40848 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_442
timestamp 1586364061
transform 1 0 41768 0 -1 42976
box -38 -48 406 592
use scs8hd_fill_1  FILLER_74_446
timestamp 1586364061
transform 1 0 42136 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_74_449
timestamp 1586364061
transform 1 0 42412 0 -1 42976
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use scs8hd_fill_1  FILLER_74_457
timestamp 1586364061
transform 1 0 43148 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_468
timestamp 1586364061
transform 1 0 44160 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_480
timestamp 1586364061
transform 1 0 45264 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_492
timestamp 1586364061
transform 1 0 46368 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_504
timestamp 1586364061
transform 1 0 47472 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 48852 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_86
timestamp 1586364061
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_98
timestamp 1586364061
transform 1 0 10120 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_110
timestamp 1586364061
transform 1 0 11224 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_123
timestamp 1586364061
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_135
timestamp 1586364061
transform 1 0 13524 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_147
timestamp 1586364061
transform 1 0 14628 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_75_159
timestamp 1586364061
transform 1 0 15732 0 1 42976
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_75_163
timestamp 1586364061
transform 1 0 16100 0 1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_75_175
timestamp 1586364061
transform 1 0 17204 0 1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_75_187
timestamp 1586364061
transform 1 0 18308 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_191
timestamp 1586364061
transform 1 0 18676 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 42976
box -38 -48 866 592
use scs8hd_fill_2  FILLER_75_204
timestamp 1586364061
transform 1 0 19872 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_212
timestamp 1586364061
transform 1 0 20608 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_208
timestamp 1586364061
transform 1 0 20240 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22816 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_217
timestamp 1586364061
transform 1 0 21068 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_221
timestamp 1586364061
transform 1 0 21436 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_234
timestamp 1586364061
transform 1 0 22632 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_238
timestamp 1586364061
transform 1 0 23000 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_250
timestamp 1586364061
transform 1 0 24104 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_245
timestamp 1586364061
transform 1 0 23644 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_242
timestamp 1586364061
transform 1 0 23368 0 1 42976
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 1 42976
box -38 -48 314 592
use scs8hd_fill_2  FILLER_75_254
timestamp 1586364061
transform 1 0 24472 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 1 42976
box -38 -48 866 592
use scs8hd_fill_2  FILLER_75_267
timestamp 1586364061
transform 1 0 25668 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_278
timestamp 1586364061
transform 1 0 26680 0 1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_75_275
timestamp 1586364061
transform 1 0 26404 0 1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_75_271
timestamp 1586364061
transform 1 0 26036 0 1 42976
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26496 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25852 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_282
timestamp 1586364061
transform 1 0 27048 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26864 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 1 42976
box -38 -48 866 592
use scs8hd_fill_2  FILLER_75_293
timestamp 1586364061
transform 1 0 28060 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28244 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_301
timestamp 1586364061
transform 1 0 28796 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_297
timestamp 1586364061
transform 1 0 28428 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 42976
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 42976
box -38 -48 866 592
use scs8hd_fill_2  FILLER_75_319
timestamp 1586364061
transform 1 0 30452 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_315
timestamp 1586364061
transform 1 0 30084 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 42976
box -38 -48 222 592
use scs8hd_nor2_4  _323_
timestamp 1586364061
transform 1 0 32292 0 1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__323__A
timestamp 1586364061
transform 1 0 32108 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_323
timestamp 1586364061
transform 1 0 30820 0 1 42976
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_75_335
timestamp 1586364061
transform 1 0 31924 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_348
timestamp 1586364061
transform 1 0 33120 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 42976
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 33304 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_352
timestamp 1586364061
transform 1 0 33488 0 1 42976
box -38 -48 222 592
use scs8hd_decap_4  FILLER_75_356
timestamp 1586364061
transform 1 0 33856 0 1 42976
box -38 -48 406 592
use scs8hd_fill_2  FILLER_75_362
timestamp 1586364061
transform 1 0 34408 0 1 42976
box -38 -48 222 592
use scs8hd_fill_1  FILLER_75_383
timestamp 1586364061
transform 1 0 36340 0 1 42976
box -38 -48 130 592
use scs8hd_fill_1  FILLER_75_380
timestamp 1586364061
transform 1 0 36064 0 1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_75_376
timestamp 1586364061
transform 1 0 35696 0 1 42976
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36156 0 1 42976
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 42976
box -38 -48 866 592
use scs8hd_fill_2  FILLER_75_393
timestamp 1586364061
transform 1 0 37260 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__B
timestamp 1586364061
transform 1 0 37444 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_401
timestamp 1586364061
transform 1 0 37996 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_397
timestamp 1586364061
transform 1 0 37628 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__377__B
timestamp 1586364061
transform 1 0 37812 0 1 42976
box -38 -48 222 592
use scs8hd_nor2_4  _372_
timestamp 1586364061
transform 1 0 38364 0 1 42976
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 42976
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__A
timestamp 1586364061
transform 1 0 38180 0 1 42976
box -38 -48 222 592
use scs8hd_decap_8  FILLER_75_414
timestamp 1586364061
transform 1 0 39192 0 1 42976
box -38 -48 774 592
use scs8hd_decap_3  FILLER_75_422
timestamp 1586364061
transform 1 0 39928 0 1 42976
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 1 42976
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42688 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41032 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 1 42976
box -38 -48 222 592
use scs8hd_decap_3  FILLER_75_431
timestamp 1586364061
transform 1 0 40756 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_436
timestamp 1586364061
transform 1 0 41216 0 1 42976
box -38 -48 314 592
use scs8hd_fill_2  FILLER_75_450
timestamp 1586364061
transform 1 0 42504 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_454
timestamp 1586364061
transform 1 0 42872 0 1 42976
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43240 0 1 42976
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 42976
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44068 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_461
timestamp 1586364061
transform 1 0 43516 0 1 42976
box -38 -48 222 592
use scs8hd_fill_2  FILLER_75_465
timestamp 1586364061
transform 1 0 43884 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_469
timestamp 1586364061
transform 1 0 44252 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_75_481
timestamp 1586364061
transform 1 0 45356 0 1 42976
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use scs8hd_fill_1  FILLER_75_487
timestamp 1586364061
transform 1 0 45908 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_489
timestamp 1586364061
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_501
timestamp 1586364061
transform 1 0 47196 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 48852 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_513
timestamp 1586364061
transform 1 0 48300 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_93
timestamp 1586364061
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_105
timestamp 1586364061
transform 1 0 10764 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_117
timestamp 1586364061
transform 1 0 11868 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_129
timestamp 1586364061
transform 1 0 12972 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_141
timestamp 1586364061
transform 1 0 14076 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_154
timestamp 1586364061
transform 1 0 15272 0 -1 44064
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_76_168
timestamp 1586364061
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_180
timestamp 1586364061
transform 1 0 17664 0 -1 44064
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 44064
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_3  FILLER_76_192
timestamp 1586364061
transform 1 0 18768 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_8  FILLER_76_204
timestamp 1586364061
transform 1 0 19872 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_2  FILLER_76_212
timestamp 1586364061
transform 1 0 20608 0 -1 44064
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 -1 44064
box -38 -48 866 592
use scs8hd_decap_8  FILLER_76_215
timestamp 1586364061
transform 1 0 20884 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_2  FILLER_76_223
timestamp 1586364061
transform 1 0 21620 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_76_234
timestamp 1586364061
transform 1 0 22632 0 -1 44064
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24840 0 -1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_76_246
timestamp 1586364061
transform 1 0 23736 0 -1 44064
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_76_261
timestamp 1586364061
transform 1 0 25116 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_265
timestamp 1586364061
transform 1 0 25484 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_76_276
timestamp 1586364061
transform 1 0 26496 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_6  FILLER_76_269
timestamp 1586364061
transform 1 0 25852 0 -1 44064
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_76_287
timestamp 1586364061
transform 1 0 27508 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_283
timestamp 1586364061
transform 1 0 27140 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27324 0 -1 44064
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_4  FILLER_76_291
timestamp 1586364061
transform 1 0 27876 0 -1 44064
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 -1 44064
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 44064
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 29992 0 -1 44064
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_304
timestamp 1586364061
transform 1 0 29072 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_6  FILLER_76_308
timestamp 1586364061
transform 1 0 29440 0 -1 44064
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 33028 0 -1 44064
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__338__A
timestamp 1586364061
transform 1 0 32292 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__388__B
timestamp 1586364061
transform 1 0 31188 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_325
timestamp 1586364061
transform 1 0 31004 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_6  FILLER_76_329
timestamp 1586364061
transform 1 0 31372 0 -1 44064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_76_335
timestamp 1586364061
transform 1 0 31924 0 -1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_76_337
timestamp 1586364061
transform 1 0 32108 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_6  FILLER_76_341
timestamp 1586364061
transform 1 0 32476 0 -1 44064
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34776 0 -1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35236 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_8  FILLER_76_358
timestamp 1586364061
transform 1 0 34040 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_2  FILLER_76_369
timestamp 1586364061
transform 1 0 35052 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_6  FILLER_76_373
timestamp 1586364061
transform 1 0 35420 0 -1 44064
box -38 -48 590 592
use scs8hd_fill_2  FILLER_76_384
timestamp 1586364061
transform 1 0 36432 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35972 0 -1 44064
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36156 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_4  FILLER_76_392
timestamp 1586364061
transform 1 0 37168 0 -1 44064
box -38 -48 406 592
use scs8hd_fill_2  FILLER_76_388
timestamp 1586364061
transform 1 0 36800 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36984 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_8  FILLER_76_398
timestamp 1586364061
transform 1 0 37720 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_1  FILLER_76_396
timestamp 1586364061
transform 1 0 37536 0 -1 44064
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use scs8hd_nor2_4  _377_
timestamp 1586364061
transform 1 0 38456 0 -1 44064
box -38 -48 866 592
use scs8hd_conb_1  _652_
timestamp 1586364061
transform 1 0 40020 0 -1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39468 0 -1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_76_415
timestamp 1586364061
transform 1 0 39284 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_76_419
timestamp 1586364061
transform 1 0 39652 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_8  FILLER_76_426
timestamp 1586364061
transform 1 0 40296 0 -1 44064
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41032 0 -1 44064
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42688 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_76_437
timestamp 1586364061
transform 1 0 41308 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_4  FILLER_76_443
timestamp 1586364061
transform 1 0 41860 0 -1 44064
box -38 -48 406 592
use scs8hd_fill_2  FILLER_76_450
timestamp 1586364061
transform 1 0 42504 0 -1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_76_454
timestamp 1586364061
transform 1 0 42872 0 -1 44064
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 44064
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 43240 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_468
timestamp 1586364061
transform 1 0 44160 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_480
timestamp 1586364061
transform 1 0 45264 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_492
timestamp 1586364061
transform 1 0 46368 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_504
timestamp 1586364061
transform 1 0 47472 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 48852 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_86
timestamp 1586364061
transform 1 0 9016 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_98
timestamp 1586364061
transform 1 0 10120 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_110
timestamp 1586364061
transform 1 0 11224 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_123
timestamp 1586364061
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_135
timestamp 1586364061
transform 1 0 13524 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_147
timestamp 1586364061
transform 1 0 14628 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_159
timestamp 1586364061
transform 1 0 15732 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_171
timestamp 1586364061
transform 1 0 16836 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_77_184
timestamp 1586364061
transform 1 0 18032 0 1 44064
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 44064
box -38 -48 222 592
use scs8hd_fill_1  FILLER_77_190
timestamp 1586364061
transform 1 0 18584 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_194
timestamp 1586364061
transform 1 0 18952 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_198
timestamp 1586364061
transform 1 0 19320 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_210
timestamp 1586364061
transform 1 0 20424 0 1 44064
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21712 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_222
timestamp 1586364061
transform 1 0 21528 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_227
timestamp 1586364061
transform 1 0 21988 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_231
timestamp 1586364061
transform 1 0 22356 0 1 44064
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_77_249
timestamp 1586364061
transform 1 0 24012 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_245
timestamp 1586364061
transform 1 0 23644 0 1 44064
box -38 -48 222 592
use scs8hd_fill_1  FILLER_77_243
timestamp 1586364061
transform 1 0 23460 0 1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 44064
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24104 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_257
timestamp 1586364061
transform 1 0 24748 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_253
timestamp 1586364061
transform 1 0 24380 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 44064
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25116 0 1 44064
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 44064
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26956 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_270
timestamp 1586364061
transform 1 0 25944 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_77_274
timestamp 1586364061
transform 1 0 26312 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_279
timestamp 1586364061
transform 1 0 26772 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_283
timestamp 1586364061
transform 1 0 27140 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_294
timestamp 1586364061
transform 1 0 28152 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_77_302
timestamp 1586364061
transform 1 0 28888 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_298
timestamp 1586364061
transform 1 0 28520 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28704 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28336 0 1 44064
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_318
timestamp 1586364061
transform 1 0 30360 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_77_313
timestamp 1586364061
transform 1 0 29900 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_309
timestamp 1586364061
transform 1 0 29532 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__388__A
timestamp 1586364061
transform 1 0 30176 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 30544 0 1 44064
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 30728 0 1 44064
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32476 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32936 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__338__B
timestamp 1586364061
transform 1 0 32108 0 1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_77_333
timestamp 1586364061
transform 1 0 31740 0 1 44064
box -38 -48 406 592
use scs8hd_fill_2  FILLER_77_339
timestamp 1586364061
transform 1 0 32292 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_344
timestamp 1586364061
transform 1 0 32752 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_348
timestamp 1586364061
transform 1 0 33120 0 1 44064
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33488 0 1 44064
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 44064
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34316 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_355
timestamp 1586364061
transform 1 0 33764 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_359
timestamp 1586364061
transform 1 0 34132 0 1 44064
box -38 -48 222 592
use scs8hd_decap_3  FILLER_77_363
timestamp 1586364061
transform 1 0 34500 0 1 44064
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 44064
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_376
timestamp 1586364061
transform 1 0 35696 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_380
timestamp 1586364061
transform 1 0 36064 0 1 44064
box -38 -48 222 592
use scs8hd_decap_4  FILLER_77_393
timestamp 1586364061
transform 1 0 37260 0 1 44064
box -38 -48 406 592
use scs8hd_fill_1  FILLER_77_397
timestamp 1586364061
transform 1 0 37628 0 1 44064
box -38 -48 130 592
use scs8hd_decap_6  FILLER_77_400
timestamp 1586364061
transform 1 0 37904 0 1 44064
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 38640 0 1 44064
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 44064
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 40388 0 1 44064
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 38456 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_419
timestamp 1586364061
transform 1 0 39652 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_423
timestamp 1586364061
transform 1 0 40020 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_435
timestamp 1586364061
transform 1 0 41124 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_431
timestamp 1586364061
transform 1 0 40756 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 44064
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41492 0 1 44064
box -38 -48 314 592
use scs8hd_fill_2  FILLER_77_446
timestamp 1586364061
transform 1 0 42136 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_442
timestamp 1586364061
transform 1 0 41768 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42320 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41952 0 1 44064
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42504 0 1 44064
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44068 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44528 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 44064
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43884 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_459
timestamp 1586364061
transform 1 0 43332 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_463
timestamp 1586364061
transform 1 0 43700 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_470
timestamp 1586364061
transform 1 0 44344 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_474
timestamp 1586364061
transform 1 0 44712 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 46000 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_486
timestamp 1586364061
transform 1 0 45816 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_489
timestamp 1586364061
transform 1 0 46092 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_501
timestamp 1586364061
transform 1 0 47196 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 48852 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  FILLER_77_513
timestamp 1586364061
transform 1 0 48300 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_93
timestamp 1586364061
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_105
timestamp 1586364061
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_117
timestamp 1586364061
transform 1 0 11868 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_129
timestamp 1586364061
transform 1 0 12972 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_141
timestamp 1586364061
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_154
timestamp 1586364061
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_166
timestamp 1586364061
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_178
timestamp 1586364061
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_190
timestamp 1586364061
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_202
timestamp 1586364061
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_215
timestamp 1586364061
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_227
timestamp 1586364061
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_78_239
timestamp 1586364061
transform 1 0 23092 0 -1 45152
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 45152
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 45152
box -38 -48 866 592
use scs8hd_decap_8  FILLER_78_250
timestamp 1586364061
transform 1 0 24104 0 -1 45152
box -38 -48 774 592
use scs8hd_decap_8  FILLER_78_267
timestamp 1586364061
transform 1 0 25668 0 -1 45152
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26956 0 -1 45152
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 45152
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27600 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_4  FILLER_78_276
timestamp 1586364061
transform 1 0 26496 0 -1 45152
box -38 -48 406 592
use scs8hd_fill_1  FILLER_78_280
timestamp 1586364061
transform 1 0 26864 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_284
timestamp 1586364061
transform 1 0 27232 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_4  FILLER_78_290
timestamp 1586364061
transform 1 0 27784 0 -1 45152
box -38 -48 406 592
use scs8hd_fill_1  FILLER_78_294
timestamp 1586364061
transform 1 0 28152 0 -1 45152
box -38 -48 130 592
use scs8hd_nor2_4  _388_
timestamp 1586364061
transform 1 0 30360 0 -1 45152
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29256 0 -1 45152
box -38 -48 222 592
use scs8hd_fill_2  FILLER_78_304
timestamp 1586364061
transform 1 0 29072 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_8  FILLER_78_308
timestamp 1586364061
transform 1 0 29440 0 -1 45152
box -38 -48 774 592
use scs8hd_fill_2  FILLER_78_316
timestamp 1586364061
transform 1 0 30176 0 -1 45152
box -38 -48 222 592
use scs8hd_nor2_4  _338_
timestamp 1586364061
transform 1 0 32108 0 -1 45152
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31372 0 -1 45152
box -38 -48 222 592
use scs8hd_fill_2  FILLER_78_327
timestamp 1586364061
transform 1 0 31188 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_4  FILLER_78_331
timestamp 1586364061
transform 1 0 31556 0 -1 45152
box -38 -48 406 592
use scs8hd_fill_1  FILLER_78_335
timestamp 1586364061
transform 1 0 31924 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_8  FILLER_78_346
timestamp 1586364061
transform 1 0 32936 0 -1 45152
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33948 0 -1 45152
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34960 0 -1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_3  FILLER_78_354
timestamp 1586364061
transform 1 0 33672 0 -1 45152
box -38 -48 314 592
use scs8hd_fill_2  FILLER_78_366
timestamp 1586364061
transform 1 0 34776 0 -1 45152
box -38 -48 222 592
use scs8hd_fill_2  FILLER_78_370
timestamp 1586364061
transform 1 0 35144 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_6  FILLER_78_374
timestamp 1586364061
transform 1 0 35512 0 -1 45152
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 45152
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 45152
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_8  FILLER_78_389
timestamp 1586364061
transform 1 0 36892 0 -1 45152
box -38 -48 774 592
use scs8hd_decap_6  FILLER_78_401
timestamp 1586364061
transform 1 0 37996 0 -1 45152
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 39284 0 -1 45152
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38640 0 -1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40480 0 -1 45152
box -38 -48 222 592
use scs8hd_fill_1  FILLER_78_407
timestamp 1586364061
transform 1 0 38548 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_410
timestamp 1586364061
transform 1 0 38824 0 -1 45152
box -38 -48 406 592
use scs8hd_fill_1  FILLER_78_414
timestamp 1586364061
transform 1 0 39192 0 -1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_78_426
timestamp 1586364061
transform 1 0 40296 0 -1 45152
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41032 0 -1 45152
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42320 0 -1 45152
box -38 -48 222 592
use scs8hd_decap_4  FILLER_78_430
timestamp 1586364061
transform 1 0 40664 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_4  FILLER_78_443
timestamp 1586364061
transform 1 0 41860 0 -1 45152
box -38 -48 406 592
use scs8hd_fill_1  FILLER_78_447
timestamp 1586364061
transform 1 0 42228 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_8  FILLER_78_450
timestamp 1586364061
transform 1 0 42504 0 -1 45152
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 45152
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 43240 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_468
timestamp 1586364061
transform 1 0 44160 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_480
timestamp 1586364061
transform 1 0 45264 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_492
timestamp 1586364061
transform 1 0 46368 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_504
timestamp 1586364061
transform 1 0 47472 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 48852 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_86
timestamp 1586364061
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_98
timestamp 1586364061
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_93
timestamp 1586364061
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_105
timestamp 1586364061
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_110
timestamp 1586364061
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_123
timestamp 1586364061
transform 1 0 12420 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_117
timestamp 1586364061
transform 1 0 11868 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_129
timestamp 1586364061
transform 1 0 12972 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_135
timestamp 1586364061
transform 1 0 13524 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_147
timestamp 1586364061
transform 1 0 14628 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_159
timestamp 1586364061
transform 1 0 15732 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_141
timestamp 1586364061
transform 1 0 14076 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_154
timestamp 1586364061
transform 1 0 15272 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_171
timestamp 1586364061
transform 1 0 16836 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_184
timestamp 1586364061
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_166
timestamp 1586364061
transform 1 0 16376 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_178
timestamp 1586364061
transform 1 0 17480 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_196
timestamp 1586364061
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_208
timestamp 1586364061
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_190
timestamp 1586364061
transform 1 0 18584 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_202
timestamp 1586364061
transform 1 0 19688 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_220
timestamp 1586364061
transform 1 0 21344 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_232
timestamp 1586364061
transform 1 0 22448 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_215
timestamp 1586364061
transform 1 0 20884 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_227
timestamp 1586364061
transform 1 0 21988 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_239
timestamp 1586364061
transform 1 0 23092 0 -1 46240
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 45152
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 -1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_245
timestamp 1586364061
transform 1 0 23644 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_79_257
timestamp 1586364061
transform 1 0 24748 0 1 45152
box -38 -48 314 592
use scs8hd_decap_8  FILLER_80_251
timestamp 1586364061
transform 1 0 24196 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  FILLER_80_259
timestamp 1586364061
transform 1 0 24932 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_8  FILLER_80_264
timestamp 1586364061
transform 1 0 25392 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_8  FILLER_80_276
timestamp 1586364061
transform 1 0 26496 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  FILLER_80_272
timestamp 1586364061
transform 1 0 26128 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_8  FILLER_79_271
timestamp 1586364061
transform 1 0 26036 0 1 45152
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_8  FILLER_80_287
timestamp 1586364061
transform 1 0 27508 0 -1 46240
box -38 -48 774 592
use scs8hd_fill_2  FILLER_79_284
timestamp 1586364061
transform 1 0 27232 0 1 45152
box -38 -48 222 592
use scs8hd_decap_3  FILLER_79_279
timestamp 1586364061
transform 1 0 26772 0 1 45152
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 45152
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 45152
box -38 -48 866 592
use scs8hd_conb_1  _651_
timestamp 1586364061
transform 1 0 27232 0 -1 46240
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 46240
box -38 -48 866 592
use scs8hd_decap_8  FILLER_80_304
timestamp 1586364061
transform 1 0 29072 0 -1 46240
box -38 -48 774 592
use scs8hd_fill_2  FILLER_79_301
timestamp 1586364061
transform 1 0 28796 0 1 45152
box -38 -48 222 592
use scs8hd_fill_2  FILLER_79_297
timestamp 1586364061
transform 1 0 28428 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29256 0 1 45152
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_80_312
timestamp 1586364061
transform 1 0 29808 0 -1 46240
box -38 -48 314 592
use scs8hd_fill_2  FILLER_79_317
timestamp 1586364061
transform 1 0 30268 0 1 45152
box -38 -48 222 592
use scs8hd_nor2_4  _393_
timestamp 1586364061
transform 1 0 30084 0 -1 46240
box -38 -48 866 592
use scs8hd_fill_2  FILLER_79_321
timestamp 1586364061
transform 1 0 30636 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__393__A
timestamp 1586364061
transform 1 0 30452 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_80_324
timestamp 1586364061
transform 1 0 30912 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_325
timestamp 1586364061
transform 1 0 31004 0 1 45152
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__393__B
timestamp 1586364061
transform 1 0 30820 0 1 45152
box -38 -48 222 592
use scs8hd_decap_8  FILLER_80_346
timestamp 1586364061
transform 1 0 32936 0 -1 46240
box -38 -48 774 592
use scs8hd_fill_1  FILLER_80_343
timestamp 1586364061
transform 1 0 32660 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_6  FILLER_80_337
timestamp 1586364061
transform 1 0 32108 0 -1 46240
box -38 -48 590 592
use scs8hd_fill_1  FILLER_79_341
timestamp 1586364061
transform 1 0 32476 0 1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_79_337
timestamp 1586364061
transform 1 0 32108 0 1 45152
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32752 0 -1 46240
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32752 0 1 45152
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_80_354
timestamp 1586364061
transform 1 0 33672 0 -1 46240
box -38 -48 222 592
use scs8hd_decap_4  FILLER_79_360
timestamp 1586364061
transform 1 0 34224 0 1 45152
box -38 -48 406 592
use scs8hd_decap_3  FILLER_79_355
timestamp 1586364061
transform 1 0 33764 0 1 45152
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 -1 46240
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34040 0 1 45152
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34040 0 -1 46240
box -38 -48 866 592
use scs8hd_decap_12  FILLER_80_367
timestamp 1586364061
transform 1 0 34868 0 -1 46240
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 45152
box -38 -48 866 592
use scs8hd_fill_2  FILLER_80_383
timestamp 1586364061
transform 1 0 36340 0 -1 46240
box -38 -48 222 592
use scs8hd_fill_1  FILLER_80_379
timestamp 1586364061
transform 1 0 35972 0 -1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_382
timestamp 1586364061
transform 1 0 36248 0 1 45152
box -38 -48 222 592
use scs8hd_decap_4  FILLER_79_376
timestamp 1586364061
transform 1 0 35696 0 1 45152
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36524 0 -1 46240
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36064 0 1 45152
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 45152
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36064 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_6  FILLER_80_391
timestamp 1586364061
transform 1 0 37076 0 -1 46240
box -38 -48 590 592
use scs8hd_fill_2  FILLER_80_387
timestamp 1586364061
transform 1 0 36708 0 -1 46240
box -38 -48 222 592
use scs8hd_decap_6  FILLER_79_393
timestamp 1586364061
transform 1 0 37260 0 1 45152
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 -1 46240
box -38 -48 222 592
use scs8hd_decap_3  FILLER_80_398
timestamp 1586364061
transform 1 0 37720 0 -1 46240
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37996 0 -1 46240
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37812 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37996 0 1 45152
box -38 -48 866 592
use scs8hd_decap_6  FILLER_80_415
timestamp 1586364061
transform 1 0 39284 0 -1 46240
box -38 -48 590 592
use scs8hd_decap_12  FILLER_80_403
timestamp 1586364061
transform 1 0 38180 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_410
timestamp 1586364061
transform 1 0 38824 0 1 45152
box -38 -48 774 592
use scs8hd_decap_12  FILLER_80_424
timestamp 1586364061
transform 1 0 40112 0 -1 46240
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_79_423
timestamp 1586364061
transform 1 0 40020 0 1 45152
box -38 -48 222 592
use scs8hd_decap_3  FILLER_79_418
timestamp 1586364061
transform 1 0 39560 0 1 45152
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 40388 0 1 45152
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 45152
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39836 0 -1 46240
box -38 -48 314 592
use scs8hd_fill_2  FILLER_80_436
timestamp 1586364061
transform 1 0 41216 0 -1 46240
box -38 -48 222 592
use scs8hd_decap_4  FILLER_79_437
timestamp 1586364061
transform 1 0 41308 0 1 45152
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41400 0 -1 46240
box -38 -48 222 592
use scs8hd_fill_1  FILLER_80_440
timestamp 1586364061
transform 1 0 41584 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  FILLER_79_443
timestamp 1586364061
transform 1 0 41860 0 1 45152
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42136 0 1 45152
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 46240
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42320 0 1 45152
box -38 -48 866 592
use scs8hd_decap_8  FILLER_80_450
timestamp 1586364061
transform 1 0 42504 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_12  FILLER_80_459
timestamp 1586364061
transform 1 0 43332 0 -1 46240
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_79_468
timestamp 1586364061
transform 1 0 44160 0 1 45152
box -38 -48 222 592
use scs8hd_decap_4  FILLER_79_461
timestamp 1586364061
transform 1 0 43516 0 1 45152
box -38 -48 406 592
use scs8hd_fill_2  FILLER_79_457
timestamp 1586364061
transform 1 0 43148 0 1 45152
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43332 0 1 45152
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 43240 0 -1 46240
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43884 0 1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_80_471
timestamp 1586364061
transform 1 0 44436 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_472
timestamp 1586364061
transform 1 0 44528 0 1 45152
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44344 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_80_483
timestamp 1586364061
transform 1 0 45540 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 46000 0 1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_79_484
timestamp 1586364061
transform 1 0 45632 0 1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_79_489
timestamp 1586364061
transform 1 0 46092 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_501
timestamp 1586364061
transform 1 0 47196 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_495
timestamp 1586364061
transform 1 0 46644 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_80_507
timestamp 1586364061
transform 1 0 47748 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 48852 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 48852 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_79_513
timestamp 1586364061
transform 1 0 48300 0 1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_80_515
timestamp 1586364061
transform 1 0 48484 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_86
timestamp 1586364061
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_98
timestamp 1586364061
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_110
timestamp 1586364061
transform 1 0 11224 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_123
timestamp 1586364061
transform 1 0 12420 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_135
timestamp 1586364061
transform 1 0 13524 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_147
timestamp 1586364061
transform 1 0 14628 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_159
timestamp 1586364061
transform 1 0 15732 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_171
timestamp 1586364061
transform 1 0 16836 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_184
timestamp 1586364061
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_196
timestamp 1586364061
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_208
timestamp 1586364061
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_220
timestamp 1586364061
transform 1 0 21344 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_232
timestamp 1586364061
transform 1 0 22448 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_245
timestamp 1586364061
transform 1 0 23644 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_257
timestamp 1586364061
transform 1 0 24748 0 1 46240
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_269
timestamp 1586364061
transform 1 0 25852 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_281
timestamp 1586364061
transform 1 0 26956 0 1 46240
box -38 -48 774 592
use scs8hd_fill_2  FILLER_81_289
timestamp 1586364061
transform 1 0 27692 0 1 46240
box -38 -48 222 592
use scs8hd_fill_2  FILLER_81_294
timestamp 1586364061
transform 1 0 28152 0 1 46240
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 1 46240
box -38 -48 222 592
use scs8hd_decap_6  FILLER_81_298
timestamp 1586364061
transform 1 0 28520 0 1 46240
box -38 -48 590 592
use scs8hd_fill_1  FILLER_81_304
timestamp 1586364061
transform 1 0 29072 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_306
timestamp 1586364061
transform 1 0 29256 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_318
timestamp 1586364061
transform 1 0 30360 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_330
timestamp 1586364061
transform 1 0 31464 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_342
timestamp 1586364061
transform 1 0 32568 0 1 46240
box -38 -48 1142 592
use scs8hd_conb_1  _655_
timestamp 1586364061
transform 1 0 34868 0 1 46240
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_354
timestamp 1586364061
transform 1 0 33672 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_370
timestamp 1586364061
transform 1 0 35144 0 1 46240
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35972 0 1 46240
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36432 0 1 46240
box -38 -48 222 592
use scs8hd_fill_1  FILLER_81_378
timestamp 1586364061
transform 1 0 35880 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_382
timestamp 1586364061
transform 1 0 36248 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_386
timestamp 1586364061
transform 1 0 36616 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_398
timestamp 1586364061
transform 1 0 37720 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 40388 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_410
timestamp 1586364061
transform 1 0 38824 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_81_422
timestamp 1586364061
transform 1 0 39928 0 1 46240
box -38 -48 406 592
use scs8hd_fill_1  FILLER_81_426
timestamp 1586364061
transform 1 0 40296 0 1 46240
box -38 -48 130 592
use scs8hd_decap_3  FILLER_81_428
timestamp 1586364061
transform 1 0 40480 0 1 46240
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41400 0 1 46240
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 1 46240
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40756 0 1 46240
box -38 -48 222 592
use scs8hd_fill_2  FILLER_81_433
timestamp 1586364061
transform 1 0 40940 0 1 46240
box -38 -48 222 592
use scs8hd_fill_1  FILLER_81_437
timestamp 1586364061
transform 1 0 41308 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_447
timestamp 1586364061
transform 1 0 42228 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_459
timestamp 1586364061
transform 1 0 43332 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_471
timestamp 1586364061
transform 1 0 44436 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_81_483
timestamp 1586364061
transform 1 0 45540 0 1 46240
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 46000 0 1 46240
box -38 -48 130 592
use scs8hd_fill_1  FILLER_81_487
timestamp 1586364061
transform 1 0 45908 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_489
timestamp 1586364061
transform 1 0 46092 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_501
timestamp 1586364061
transform 1 0 47196 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 48852 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_81_513
timestamp 1586364061
transform 1 0 48300 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 6808 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_63
timestamp 1586364061
transform 1 0 6900 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_75
timestamp 1586364061
transform 1 0 8004 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 9660 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_87
timestamp 1586364061
transform 1 0 9108 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_94
timestamp 1586364061
transform 1 0 9752 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_106
timestamp 1586364061
transform 1 0 10856 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 12512 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_118
timestamp 1586364061
transform 1 0 11960 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_125
timestamp 1586364061
transform 1 0 12604 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 15364 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_137
timestamp 1586364061
transform 1 0 13708 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_149
timestamp 1586364061
transform 1 0 14812 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_156
timestamp 1586364061
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 18216 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_168
timestamp 1586364061
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_180
timestamp 1586364061
transform 1 0 17664 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_187
timestamp 1586364061
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_199
timestamp 1586364061
transform 1 0 19412 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_211
timestamp 1586364061
transform 1 0 20516 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 21068 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_218
timestamp 1586364061
transform 1 0 21160 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_230
timestamp 1586364061
transform 1 0 22264 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 23920 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_242
timestamp 1586364061
transform 1 0 23368 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_249
timestamp 1586364061
transform 1 0 24012 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_261
timestamp 1586364061
transform 1 0 25116 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 26772 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_273
timestamp 1586364061
transform 1 0 26220 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_280
timestamp 1586364061
transform 1 0 26864 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_292
timestamp 1586364061
transform 1 0 27968 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 29624 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_304
timestamp 1586364061
transform 1 0 29072 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_311
timestamp 1586364061
transform 1 0 29716 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 32476 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_323
timestamp 1586364061
transform 1 0 30820 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_335
timestamp 1586364061
transform 1 0 31924 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_342
timestamp 1586364061
transform 1 0 32568 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 35328 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_354
timestamp 1586364061
transform 1 0 33672 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_366
timestamp 1586364061
transform 1 0 34776 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_373
timestamp 1586364061
transform 1 0 35420 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_385
timestamp 1586364061
transform 1 0 36524 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_397
timestamp 1586364061
transform 1 0 37628 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 38180 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_404
timestamp 1586364061
transform 1 0 38272 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_416
timestamp 1586364061
transform 1 0 39376 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_428
timestamp 1586364061
transform 1 0 40480 0 -1 47328
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41124 0 -1 47328
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 41032 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_438
timestamp 1586364061
transform 1 0 41400 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_450
timestamp 1586364061
transform 1 0 42504 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 43884 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_3  FILLER_82_462
timestamp 1586364061
transform 1 0 43608 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_466
timestamp 1586364061
transform 1 0 43976 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_478
timestamp 1586364061
transform 1 0 45080 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 46736 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_490
timestamp 1586364061
transform 1 0 46184 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_497
timestamp 1586364061
transform 1 0 46828 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_509
timestamp 1586364061
transform 1 0 47932 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 48852 0 -1 47328
box -38 -48 314 592
use scs8hd_fill_1  FILLER_82_515
timestamp 1586364061
transform 1 0 48484 0 -1 47328
box -38 -48 130 592
<< labels >>
rlabel metal3 s 49520 17144 50000 17264 6 address[0]
port 0 nsew default input
rlabel metal3 s 49520 20272 50000 20392 6 address[1]
port 1 nsew default input
rlabel metal3 s 49520 23400 50000 23520 6 address[2]
port 2 nsew default input
rlabel metal3 s 49520 26528 50000 26648 6 address[3]
port 3 nsew default input
rlabel metal3 s 49520 29656 50000 29776 6 address[4]
port 4 nsew default input
rlabel metal3 s 49520 32784 50000 32904 6 address[5]
port 5 nsew default input
rlabel metal3 s 49520 35912 50000 36032 6 address[6]
port 6 nsew default input
rlabel metal3 s 49520 39040 50000 39160 6 address[7]
port 7 nsew default input
rlabel metal3 s 49520 42168 50000 42288 6 address[8]
port 8 nsew default input
rlabel metal3 s 49520 45296 50000 45416 6 address[9]
port 9 nsew default input
rlabel metal2 s 39118 0 39174 480 6 bottom_width_0_height_0__pin_10_
port 10 nsew default tristate
rlabel metal2 s 46294 0 46350 480 6 bottom_width_0_height_0__pin_14_
port 11 nsew default input
rlabel metal2 s 24858 0 24914 480 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal2 s 32034 0 32090 480 6 bottom_width_0_height_0__pin_6_
port 13 nsew default input
rlabel metal2 s 17774 0 17830 480 6 clk
port 14 nsew default input
rlabel metal3 s 49520 48424 50000 48544 6 data_in
port 15 nsew default input
rlabel metal3 s 49520 14016 50000 14136 6 enable
port 16 nsew default input
rlabel metal3 s 0 41624 480 41744 6 left_width_0_height_0__pin_11_
port 17 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 left_width_0_height_0__pin_3_
port 18 nsew default input
rlabel metal3 s 0 24896 480 25016 6 left_width_0_height_0__pin_7_
port 19 nsew default input
rlabel metal2 s 10598 0 10654 480 6 reset
port 20 nsew default input
rlabel metal3 s 49520 10888 50000 11008 6 right_width_0_height_0__pin_13_
port 21 nsew default tristate
rlabel metal3 s 49520 1504 50000 1624 6 right_width_0_height_0__pin_1_
port 22 nsew default input
rlabel metal3 s 49520 4632 50000 4752 6 right_width_0_height_0__pin_5_
port 23 nsew default input
rlabel metal3 s 49520 7760 50000 7880 6 right_width_0_height_0__pin_9_
port 24 nsew default input
rlabel metal2 s 3514 0 3570 480 6 set
port 25 nsew default input
rlabel metal2 s 6182 49520 6238 50000 6 top_width_0_height_0__pin_0_
port 26 nsew default input
rlabel metal2 s 43626 49520 43682 50000 6 top_width_0_height_0__pin_12_
port 27 nsew default tristate
rlabel metal2 s 18602 49520 18658 50000 6 top_width_0_height_0__pin_4_
port 28 nsew default input
rlabel metal2 s 31114 49520 31170 50000 6 top_width_0_height_0__pin_8_
port 29 nsew default input
rlabel metal4 s 4208 2128 4528 47376 6 vpwr
port 30 nsew default input
rlabel metal4 s 19568 2128 19888 47376 6 vgnd
port 31 nsew default input
<< end >>
