magic
tech sky130A
magscale 1 2
timestamp 1606475217
<< locali >>
rect 1961 14263 1995 14433
rect 4629 12767 4663 12869
rect 6653 12631 6687 12869
rect 13829 12631 13863 12937
rect 5917 11135 5951 11305
rect 7573 11135 7607 11305
rect 12265 10455 12299 10761
rect 18429 9911 18463 10149
rect 7757 8891 7791 9061
rect 16681 8279 16715 8381
rect 9505 7735 9539 7837
rect 13553 7803 13587 8041
rect 10057 7191 10091 7429
rect 13645 7191 13679 7293
rect 17509 6647 17543 6885
rect 17601 6647 17635 6749
rect 13921 6171 13955 6341
rect 17601 5763 17635 5865
rect 19257 5627 19291 5865
rect 6561 5083 6595 5253
rect 18245 4607 18279 4777
rect 5457 4063 5491 4233
rect 12357 3383 12391 3689
rect 6653 2907 6687 3145
rect 13001 2907 13035 3145
<< viali >>
rect 1961 19465 1995 19499
rect 5825 19465 5859 19499
rect 19165 19465 19199 19499
rect 20729 19465 20763 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 5641 19261 5675 19295
rect 18981 19261 19015 19295
rect 20545 19261 20579 19295
rect 2513 19125 2547 19159
rect 1961 18921 1995 18955
rect 6285 18853 6319 18887
rect 18429 18853 18463 18887
rect 1777 18785 1811 18819
rect 6009 18785 6043 18819
rect 18153 18785 18187 18819
rect 1961 18377 1995 18411
rect 20729 18377 20763 18411
rect 1777 18173 1811 18207
rect 20545 18173 20579 18207
rect 2421 17765 2455 17799
rect 19901 17765 19935 17799
rect 1593 17697 1627 17731
rect 2145 17697 2179 17731
rect 19625 17697 19659 17731
rect 1777 17561 1811 17595
rect 1961 17289 1995 17323
rect 20729 17289 20763 17323
rect 1777 17085 1811 17119
rect 20545 17085 20579 17119
rect 1961 16745 1995 16779
rect 20453 16745 20487 16779
rect 1777 16609 1811 16643
rect 20269 16609 20303 16643
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 3341 16201 3375 16235
rect 13553 16201 13587 16235
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 1777 15997 1811 16031
rect 2335 15997 2369 16031
rect 3157 15997 3191 16031
rect 13369 15997 13403 16031
rect 19993 15997 20027 16031
rect 20545 15997 20579 16031
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 20453 15657 20487 15691
rect 4353 15589 4387 15623
rect 12817 15589 12851 15623
rect 1777 15521 1811 15555
rect 2335 15521 2369 15555
rect 4077 15521 4111 15555
rect 12541 15521 12575 15555
rect 19717 15521 19751 15555
rect 20269 15521 20303 15555
rect 19901 15317 19935 15351
rect 2513 15113 2547 15147
rect 20177 15113 20211 15147
rect 20729 15113 20763 15147
rect 1961 15045 1995 15079
rect 19625 15045 19659 15079
rect 2973 14977 3007 15011
rect 16773 14977 16807 15011
rect 1777 14909 1811 14943
rect 2335 14909 2369 14943
rect 19441 14909 19475 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 3240 14841 3274 14875
rect 16681 14841 16715 14875
rect 4353 14773 4387 14807
rect 16221 14773 16255 14807
rect 16589 14773 16623 14807
rect 1685 14569 1719 14603
rect 4261 14569 4295 14603
rect 19349 14569 19383 14603
rect 2329 14501 2363 14535
rect 7573 14501 7607 14535
rect 19993 14501 20027 14535
rect 1501 14433 1535 14467
rect 1961 14433 1995 14467
rect 2053 14433 2087 14467
rect 3249 14433 3283 14467
rect 4077 14433 4111 14467
rect 10425 14433 10459 14467
rect 11805 14433 11839 14467
rect 12061 14433 12095 14467
rect 14289 14433 14323 14467
rect 14381 14433 14415 14467
rect 16028 14433 16062 14467
rect 18613 14433 18647 14467
rect 19165 14433 19199 14467
rect 19717 14433 19751 14467
rect 3341 14365 3375 14399
rect 3525 14365 3559 14399
rect 7665 14365 7699 14399
rect 7757 14365 7791 14399
rect 10517 14365 10551 14399
rect 10701 14365 10735 14399
rect 14565 14365 14599 14399
rect 15761 14365 15795 14399
rect 1961 14229 1995 14263
rect 2881 14229 2915 14263
rect 7205 14229 7239 14263
rect 10057 14229 10091 14263
rect 13185 14229 13219 14263
rect 13921 14229 13955 14263
rect 17141 14229 17175 14263
rect 18797 14229 18831 14263
rect 11437 14025 11471 14059
rect 14749 14025 14783 14059
rect 5457 13957 5491 13991
rect 9781 13957 9815 13991
rect 16681 13957 16715 13991
rect 2421 13889 2455 13923
rect 4077 13889 4111 13923
rect 7481 13889 7515 13923
rect 17233 13889 17267 13923
rect 20085 13889 20119 13923
rect 20821 13889 20855 13923
rect 1685 13821 1719 13855
rect 1961 13821 1995 13855
rect 4333 13821 4367 13855
rect 7297 13821 7331 13855
rect 8401 13821 8435 13855
rect 8668 13821 8702 13855
rect 10057 13821 10091 13855
rect 10313 13821 10347 13855
rect 13369 13821 13403 13855
rect 13636 13821 13670 13855
rect 15025 13821 15059 13855
rect 15281 13821 15315 13855
rect 17049 13821 17083 13855
rect 18061 13821 18095 13855
rect 18797 13821 18831 13855
rect 19901 13821 19935 13855
rect 20637 13821 20671 13855
rect 2688 13753 2722 13787
rect 7205 13753 7239 13787
rect 7849 13753 7883 13787
rect 17141 13753 17175 13787
rect 18337 13753 18371 13787
rect 19073 13753 19107 13787
rect 3801 13685 3835 13719
rect 6837 13685 6871 13719
rect 16405 13685 16439 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 2973 13481 3007 13515
rect 4261 13481 4295 13515
rect 5089 13481 5123 13515
rect 6285 13481 6319 13515
rect 6653 13481 6687 13515
rect 8677 13481 8711 13515
rect 14473 13481 14507 13515
rect 15301 13481 15335 13515
rect 16405 13481 16439 13515
rect 20453 13481 20487 13515
rect 6745 13413 6779 13447
rect 10425 13413 10459 13447
rect 11222 13413 11256 13447
rect 17202 13413 17236 13447
rect 1409 13345 1443 13379
rect 2329 13345 2363 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 7297 13345 7331 13379
rect 7564 13345 7598 13379
rect 10333 13345 10367 13379
rect 13093 13345 13127 13379
rect 13360 13345 13394 13379
rect 15669 13345 15703 13379
rect 16957 13345 16991 13379
rect 18880 13345 18914 13379
rect 20269 13345 20303 13379
rect 2421 13277 2455 13311
rect 2605 13277 2639 13311
rect 3433 13277 3467 13311
rect 3525 13277 3559 13311
rect 5181 13277 5215 13311
rect 5365 13277 5399 13311
rect 6929 13277 6963 13311
rect 9137 13277 9171 13311
rect 10609 13277 10643 13311
rect 10977 13277 11011 13311
rect 12633 13277 12667 13311
rect 14749 13277 14783 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 18613 13277 18647 13311
rect 18337 13209 18371 13243
rect 4721 13141 4755 13175
rect 9965 13141 9999 13175
rect 12357 13141 12391 13175
rect 19993 13141 20027 13175
rect 2513 12937 2547 12971
rect 3801 12937 3835 12971
rect 6837 12937 6871 12971
rect 9137 12937 9171 12971
rect 13829 12937 13863 12971
rect 13921 12937 13955 12971
rect 16865 12937 16899 12971
rect 18337 12937 18371 12971
rect 4629 12869 4663 12903
rect 6193 12869 6227 12903
rect 6653 12869 6687 12903
rect 7849 12869 7883 12903
rect 12449 12869 12483 12903
rect 2053 12801 2087 12835
rect 2973 12801 3007 12835
rect 3157 12801 3191 12835
rect 4445 12801 4479 12835
rect 1777 12733 1811 12767
rect 4629 12733 4663 12767
rect 4813 12733 4847 12767
rect 2881 12665 2915 12699
rect 4169 12665 4203 12699
rect 5080 12665 5114 12699
rect 7389 12801 7423 12835
rect 8309 12801 8343 12835
rect 8493 12801 8527 12835
rect 9597 12801 9631 12835
rect 9781 12801 9815 12835
rect 10701 12801 10735 12835
rect 11897 12801 11931 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 9505 12733 9539 12767
rect 7297 12665 7331 12699
rect 8217 12665 8251 12699
rect 10517 12665 10551 12699
rect 11713 12665 11747 12699
rect 12817 12665 12851 12699
rect 14473 12801 14507 12835
rect 16313 12801 16347 12835
rect 16497 12801 16531 12835
rect 17417 12801 17451 12835
rect 18981 12801 19015 12835
rect 19901 12801 19935 12835
rect 20913 12801 20947 12835
rect 14289 12733 14323 12767
rect 20821 12733 20855 12767
rect 14381 12665 14415 12699
rect 18705 12665 18739 12699
rect 19717 12665 19751 12699
rect 20729 12665 20763 12699
rect 4261 12597 4295 12631
rect 6653 12597 6687 12631
rect 7205 12597 7239 12631
rect 10149 12597 10183 12631
rect 10609 12597 10643 12631
rect 11345 12597 11379 12631
rect 11805 12597 11839 12631
rect 13829 12597 13863 12631
rect 15853 12597 15887 12631
rect 16221 12597 16255 12631
rect 17233 12597 17267 12631
rect 17325 12597 17359 12631
rect 18797 12597 18831 12631
rect 19349 12597 19383 12631
rect 19809 12597 19843 12631
rect 20361 12597 20395 12631
rect 2421 12393 2455 12427
rect 3617 12393 3651 12427
rect 5457 12393 5491 12427
rect 7481 12393 7515 12427
rect 8125 12393 8159 12427
rect 8585 12393 8619 12427
rect 9873 12393 9907 12427
rect 10333 12393 10367 12427
rect 13001 12393 13035 12427
rect 17601 12393 17635 12427
rect 19717 12393 19751 12427
rect 20913 12393 20947 12427
rect 1961 12325 1995 12359
rect 10241 12325 10275 12359
rect 18604 12325 18638 12359
rect 1685 12257 1719 12291
rect 2789 12257 2823 12291
rect 3433 12257 3467 12291
rect 4333 12257 4367 12291
rect 6368 12257 6402 12291
rect 8493 12257 8527 12291
rect 10885 12257 10919 12291
rect 11152 12257 11186 12291
rect 12909 12257 12943 12291
rect 13553 12257 13587 12291
rect 15844 12257 15878 12291
rect 18337 12257 18371 12291
rect 19993 12257 20027 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 4077 12189 4111 12223
rect 6101 12189 6135 12223
rect 8769 12189 8803 12223
rect 10425 12189 10459 12223
rect 13093 12189 13127 12223
rect 15577 12189 15611 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 20269 12189 20303 12223
rect 12265 12121 12299 12155
rect 16957 12121 16991 12155
rect 12541 12053 12575 12087
rect 17233 12053 17267 12087
rect 7481 11849 7515 11883
rect 11805 11849 11839 11883
rect 15669 11849 15703 11883
rect 18061 11849 18095 11883
rect 20913 11849 20947 11883
rect 4997 11781 5031 11815
rect 8493 11781 8527 11815
rect 12449 11781 12483 11815
rect 16037 11781 16071 11815
rect 2513 11713 2547 11747
rect 3433 11713 3467 11747
rect 4445 11713 4479 11747
rect 5549 11713 5583 11747
rect 8033 11713 8067 11747
rect 8769 11713 8803 11747
rect 13001 11713 13035 11747
rect 14289 11713 14323 11747
rect 16313 11713 16347 11747
rect 18613 11713 18647 11747
rect 5365 11645 5399 11679
rect 6193 11645 6227 11679
rect 8677 11645 8711 11679
rect 10425 11645 10459 11679
rect 12265 11645 12299 11679
rect 12817 11645 12851 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 16580 11645 16614 11679
rect 18429 11645 18463 11679
rect 19073 11645 19107 11679
rect 19340 11645 19374 11679
rect 20729 11645 20763 11679
rect 3249 11577 3283 11611
rect 4353 11577 4387 11611
rect 5457 11577 5491 11611
rect 7849 11577 7883 11611
rect 7941 11577 7975 11611
rect 9036 11577 9070 11611
rect 10670 11577 10704 11611
rect 13737 11577 13771 11611
rect 14556 11577 14590 11611
rect 1869 11509 1903 11543
rect 2237 11509 2271 11543
rect 2329 11509 2363 11543
rect 2881 11509 2915 11543
rect 3341 11509 3375 11543
rect 3893 11509 3927 11543
rect 4261 11509 4295 11543
rect 6009 11509 6043 11543
rect 10149 11509 10183 11543
rect 12081 11509 12115 11543
rect 12909 11509 12943 11543
rect 17693 11509 17727 11543
rect 18521 11509 18555 11543
rect 20453 11509 20487 11543
rect 3525 11305 3559 11339
rect 5917 11305 5951 11339
rect 7389 11305 7423 11339
rect 7573 11305 7607 11339
rect 8125 11305 8159 11339
rect 12909 11305 12943 11339
rect 15761 11305 15795 11339
rect 16313 11305 16347 11339
rect 17785 11305 17819 11339
rect 18429 11305 18463 11339
rect 18889 11305 18923 11339
rect 1869 11169 1903 11203
rect 2136 11169 2170 11203
rect 4353 11169 4387 11203
rect 4620 11169 4654 11203
rect 6265 11169 6299 11203
rect 11796 11237 11830 11271
rect 13614 11237 13648 11271
rect 15669 11237 15703 11271
rect 8033 11169 8067 11203
rect 10057 11169 10091 11203
rect 11529 11169 11563 11203
rect 13369 11169 13403 11203
rect 16681 11169 16715 11203
rect 17693 11169 17727 11203
rect 18797 11169 18831 11203
rect 20177 11169 20211 11203
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 7573 11101 7607 11135
rect 8217 11101 8251 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 15945 11101 15979 11135
rect 16773 11101 16807 11135
rect 16865 11101 16899 11135
rect 17877 11101 17911 11135
rect 18981 11101 19015 11135
rect 20269 11101 20303 11135
rect 20361 11101 20395 11135
rect 3249 11033 3283 11067
rect 5733 11033 5767 11067
rect 7665 11033 7699 11067
rect 14749 11033 14783 11067
rect 15301 11033 15335 11067
rect 17325 11033 17359 11067
rect 9689 10965 9723 10999
rect 19809 10965 19843 10999
rect 2053 10761 2087 10795
rect 3065 10761 3099 10795
rect 5457 10761 5491 10795
rect 9045 10761 9079 10795
rect 10057 10761 10091 10795
rect 12265 10761 12299 10795
rect 18705 10761 18739 10795
rect 11345 10693 11379 10727
rect 2697 10625 2731 10659
rect 3617 10625 3651 10659
rect 6193 10625 6227 10659
rect 6285 10625 6319 10659
rect 6837 10625 6871 10659
rect 9597 10625 9631 10659
rect 10609 10625 10643 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 2513 10557 2547 10591
rect 4077 10557 4111 10591
rect 9505 10557 9539 10591
rect 3433 10489 3467 10523
rect 4344 10489 4378 10523
rect 6101 10489 6135 10523
rect 7104 10489 7138 10523
rect 8585 10489 8619 10523
rect 9413 10489 9447 10523
rect 10425 10489 10459 10523
rect 15301 10693 15335 10727
rect 16405 10693 16439 10727
rect 14841 10625 14875 10659
rect 15945 10625 15979 10659
rect 16957 10625 16991 10659
rect 19165 10625 19199 10659
rect 19349 10625 19383 10659
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 15485 10557 15519 10591
rect 19073 10557 19107 10591
rect 19717 10557 19751 10591
rect 19984 10557 20018 10591
rect 14657 10489 14691 10523
rect 16773 10489 16807 10523
rect 2421 10421 2455 10455
rect 3525 10421 3559 10455
rect 5733 10421 5767 10455
rect 8217 10421 8251 10455
rect 10517 10421 10551 10455
rect 11713 10421 11747 10455
rect 12265 10421 12299 10455
rect 13829 10421 13863 10455
rect 14289 10421 14323 10455
rect 14749 10421 14783 10455
rect 16865 10421 16899 10455
rect 21097 10421 21131 10455
rect 3157 10217 3191 10251
rect 4261 10217 4295 10251
rect 4629 10217 4663 10251
rect 5273 10217 5307 10251
rect 7849 10217 7883 10251
rect 8125 10217 8159 10251
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 11989 10217 12023 10251
rect 12633 10217 12667 10251
rect 13645 10217 13679 10251
rect 14013 10217 14047 10251
rect 14473 10217 14507 10251
rect 15301 10217 15335 10251
rect 18337 10217 18371 10251
rect 20913 10217 20947 10251
rect 4721 10149 4755 10183
rect 18429 10149 18463 10183
rect 1777 10081 1811 10115
rect 2044 10081 2078 10115
rect 5641 10081 5675 10115
rect 6469 10081 6503 10115
rect 6736 10081 6770 10115
rect 8309 10081 8343 10115
rect 8861 10081 8895 10115
rect 9956 10081 9990 10115
rect 13001 10081 13035 10115
rect 13829 10081 13863 10115
rect 14381 10081 14415 10115
rect 15669 10081 15703 10115
rect 17224 10081 17258 10115
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 9137 10013 9171 10047
rect 9689 10013 9723 10047
rect 12081 10013 12115 10047
rect 12265 10013 12299 10047
rect 13093 10013 13127 10047
rect 13185 10013 13219 10047
rect 14565 10013 14599 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16957 10013 16991 10047
rect 18613 10081 18647 10115
rect 18880 10081 18914 10115
rect 20269 10081 20303 10115
rect 20453 9945 20487 9979
rect 18429 9877 18463 9911
rect 19993 9877 20027 9911
rect 1869 9673 1903 9707
rect 10241 9673 10275 9707
rect 10517 9673 10551 9707
rect 16957 9673 16991 9707
rect 18061 9673 18095 9707
rect 2881 9605 2915 9639
rect 4813 9605 4847 9639
rect 6837 9605 6871 9639
rect 14197 9605 14231 9639
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 3433 9537 3467 9571
rect 5273 9537 5307 9571
rect 5457 9537 5491 9571
rect 7481 9537 7515 9571
rect 8401 9537 8435 9571
rect 8861 9537 8895 9571
rect 11069 9537 11103 9571
rect 14749 9537 14783 9571
rect 15853 9537 15887 9571
rect 17509 9537 17543 9571
rect 18705 9537 18739 9571
rect 19717 9537 19751 9571
rect 2237 9469 2271 9503
rect 3249 9469 3283 9503
rect 8309 9469 8343 9503
rect 10977 9469 11011 9503
rect 12449 9469 12483 9503
rect 15669 9469 15703 9503
rect 19984 9469 20018 9503
rect 1409 9401 1443 9435
rect 9128 9401 9162 9435
rect 10885 9401 10919 9435
rect 12716 9401 12750 9435
rect 14565 9401 14599 9435
rect 15577 9401 15611 9435
rect 16221 9401 16255 9435
rect 17417 9401 17451 9435
rect 18521 9401 18555 9435
rect 3341 9333 3375 9367
rect 5181 9333 5215 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 7849 9333 7883 9367
rect 8217 9333 8251 9367
rect 13829 9333 13863 9367
rect 14657 9333 14691 9367
rect 15209 9333 15243 9367
rect 17325 9333 17359 9367
rect 18429 9333 18463 9367
rect 21097 9333 21131 9367
rect 2053 9129 2087 9163
rect 4537 9129 4571 9163
rect 7573 9129 7607 9163
rect 13921 9129 13955 9163
rect 14197 9129 14231 9163
rect 16681 9129 16715 9163
rect 16957 9129 16991 9163
rect 17417 9129 17451 9163
rect 19809 9129 19843 9163
rect 7757 9061 7791 9095
rect 10057 9061 10091 9095
rect 10149 9061 10183 9095
rect 12786 9061 12820 9095
rect 14565 9061 14599 9095
rect 2421 8993 2455 9027
rect 4905 8993 4939 9027
rect 5549 8993 5583 9027
rect 6193 8993 6227 9027
rect 6460 8993 6494 9027
rect 2513 8925 2547 8959
rect 2697 8925 2731 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 8217 8993 8251 9027
rect 8309 8993 8343 9027
rect 9137 8993 9171 9027
rect 10701 8993 10735 9027
rect 15557 8993 15591 9027
rect 17325 8993 17359 9027
rect 18696 8993 18730 9027
rect 20269 8993 20303 9027
rect 8493 8925 8527 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 10241 8925 10275 8959
rect 12548 8925 12582 8959
rect 14657 8925 14691 8959
rect 14749 8925 14783 8959
rect 15301 8925 15335 8959
rect 17509 8925 17543 8959
rect 18429 8925 18463 8959
rect 7757 8857 7791 8891
rect 7849 8857 7883 8891
rect 9689 8857 9723 8891
rect 20453 8857 20487 8891
rect 8769 8789 8803 8823
rect 11989 8789 12023 8823
rect 3249 8585 3283 8619
rect 4077 8585 4111 8619
rect 7941 8585 7975 8619
rect 9873 8585 9907 8619
rect 12081 8585 12115 8619
rect 12449 8585 12483 8619
rect 15853 8585 15887 8619
rect 16865 8585 16899 8619
rect 19441 8585 19475 8619
rect 19717 8585 19751 8619
rect 5089 8517 5123 8551
rect 6837 8517 6871 8551
rect 14841 8517 14875 8551
rect 4629 8449 4663 8483
rect 5641 8449 5675 8483
rect 7481 8449 7515 8483
rect 13001 8449 13035 8483
rect 13461 8449 13495 8483
rect 16405 8449 16439 8483
rect 17509 8449 17543 8483
rect 20269 8449 20303 8483
rect 1869 8381 1903 8415
rect 5457 8381 5491 8415
rect 5549 8381 5583 8415
rect 7297 8381 7331 8415
rect 8125 8381 8159 8415
rect 8493 8381 8527 8415
rect 10701 8381 10735 8415
rect 12817 8381 12851 8415
rect 16313 8381 16347 8415
rect 16681 8381 16715 8415
rect 18061 8381 18095 8415
rect 18317 8381 18351 8415
rect 20177 8381 20211 8415
rect 20729 8381 20763 8415
rect 2136 8313 2170 8347
rect 7205 8313 7239 8347
rect 8217 8313 8251 8347
rect 8760 8313 8794 8347
rect 10968 8313 11002 8347
rect 13728 8313 13762 8347
rect 20085 8313 20119 8347
rect 4445 8245 4479 8279
rect 4537 8245 4571 8279
rect 6285 8245 6319 8279
rect 12909 8245 12943 8279
rect 16221 8245 16255 8279
rect 16681 8245 16715 8279
rect 17233 8245 17267 8279
rect 17325 8245 17359 8279
rect 20913 8245 20947 8279
rect 1961 8041 1995 8075
rect 3341 8041 3375 8075
rect 4261 8041 4295 8075
rect 5273 8041 5307 8075
rect 6837 8041 6871 8075
rect 7941 8041 7975 8075
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 9873 8041 9907 8075
rect 10241 8041 10275 8075
rect 10333 8041 10367 8075
rect 11161 8041 11195 8075
rect 11529 8041 11563 8075
rect 12633 8041 12667 8075
rect 13093 8041 13127 8075
rect 13553 8041 13587 8075
rect 13645 8041 13679 8075
rect 14013 8041 14047 8075
rect 18705 8041 18739 8075
rect 3433 7973 3467 8007
rect 4629 7973 4663 8007
rect 11897 7973 11931 8007
rect 2329 7905 2363 7939
rect 5641 7905 5675 7939
rect 7849 7905 7883 7939
rect 11069 7905 11103 7939
rect 13001 7905 13035 7939
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 4721 7837 4755 7871
rect 4813 7837 4847 7871
rect 5733 7837 5767 7871
rect 5825 7837 5859 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 8033 7837 8067 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 10425 7837 10459 7871
rect 11253 7837 11287 7871
rect 11989 7837 12023 7871
rect 12173 7837 12207 7871
rect 13185 7837 13219 7871
rect 2973 7769 3007 7803
rect 6469 7769 6503 7803
rect 15936 7973 15970 8007
rect 17570 7973 17604 8007
rect 14841 7905 14875 7939
rect 15669 7905 15703 7939
rect 17325 7905 17359 7939
rect 20085 7905 20119 7939
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 19257 7837 19291 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 10701 7769 10735 7803
rect 13553 7769 13587 7803
rect 7481 7701 7515 7735
rect 9505 7701 9539 7735
rect 14657 7701 14691 7735
rect 17049 7701 17083 7735
rect 19717 7701 19751 7735
rect 2145 7497 2179 7531
rect 4905 7497 4939 7531
rect 9965 7497 9999 7531
rect 10241 7497 10275 7531
rect 15117 7497 15151 7531
rect 16221 7497 16255 7531
rect 10057 7429 10091 7463
rect 2789 7361 2823 7395
rect 3985 7361 4019 7395
rect 5457 7361 5491 7395
rect 7481 7361 7515 7395
rect 7205 7293 7239 7327
rect 8033 7293 8067 7327
rect 8585 7293 8619 7327
rect 8852 7293 8886 7327
rect 3893 7225 3927 7259
rect 5365 7225 5399 7259
rect 10793 7361 10827 7395
rect 11805 7361 11839 7395
rect 13185 7361 13219 7395
rect 13369 7361 13403 7395
rect 13737 7361 13771 7395
rect 16773 7361 16807 7395
rect 19257 7361 19291 7395
rect 20361 7361 20395 7395
rect 13093 7293 13127 7327
rect 13645 7293 13679 7327
rect 16589 7293 16623 7327
rect 16681 7293 16715 7327
rect 19073 7293 19107 7327
rect 20085 7293 20119 7327
rect 20729 7293 20763 7327
rect 11713 7225 11747 7259
rect 14004 7225 14038 7259
rect 2513 7157 2547 7191
rect 2605 7157 2639 7191
rect 3433 7157 3467 7191
rect 3801 7157 3835 7191
rect 5273 7157 5307 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 7849 7157 7883 7191
rect 10057 7157 10091 7191
rect 10609 7157 10643 7191
rect 10701 7157 10735 7191
rect 11253 7157 11287 7191
rect 11621 7157 11655 7191
rect 12725 7157 12759 7191
rect 13645 7157 13679 7191
rect 15393 7157 15427 7191
rect 18245 7157 18279 7191
rect 18705 7157 18739 7191
rect 19165 7157 19199 7191
rect 19717 7157 19751 7191
rect 20177 7157 20211 7191
rect 20913 7157 20947 7191
rect 6929 6953 6963 6987
rect 9965 6953 9999 6987
rect 13553 6953 13587 6987
rect 16037 6953 16071 6987
rect 16129 6953 16163 6987
rect 16681 6953 16715 6987
rect 17693 6953 17727 6987
rect 18613 6953 18647 6987
rect 18981 6953 19015 6987
rect 19993 6953 20027 6987
rect 4988 6885 5022 6919
rect 10333 6885 10367 6919
rect 17049 6885 17083 6919
rect 17509 6885 17543 6919
rect 20085 6885 20119 6919
rect 2145 6817 2179 6851
rect 2412 6817 2446 6851
rect 6837 6817 6871 6851
rect 7849 6817 7883 6851
rect 8861 6817 8895 6851
rect 11069 6817 11103 6851
rect 11336 6817 11370 6851
rect 14565 6817 14599 6851
rect 17141 6817 17175 6851
rect 1685 6749 1719 6783
rect 4721 6749 4755 6783
rect 7113 6749 7147 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 8953 6749 8987 6783
rect 9045 6749 9079 6783
rect 10425 6749 10459 6783
rect 10517 6749 10551 6783
rect 12725 6749 12759 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 16313 6749 16347 6783
rect 17325 6749 17359 6783
rect 6469 6681 6503 6715
rect 8493 6681 8527 6715
rect 13185 6681 13219 6715
rect 17877 6817 17911 6851
rect 18061 6817 18095 6851
rect 19073 6817 19107 6851
rect 3525 6613 3559 6647
rect 6101 6613 6135 6647
rect 7481 6613 7515 6647
rect 12449 6613 12483 6647
rect 14197 6613 14231 6647
rect 15669 6613 15703 6647
rect 17509 6613 17543 6647
rect 17601 6749 17635 6783
rect 19257 6749 19291 6783
rect 20177 6749 20211 6783
rect 18245 6681 18279 6715
rect 17601 6613 17635 6647
rect 19625 6613 19659 6647
rect 3341 6409 3375 6443
rect 6837 6409 6871 6443
rect 11253 6409 11287 6443
rect 15761 6409 15795 6443
rect 17601 6409 17635 6443
rect 20177 6409 20211 6443
rect 9597 6341 9631 6375
rect 11989 6341 12023 6375
rect 13829 6341 13863 6375
rect 13921 6341 13955 6375
rect 16037 6341 16071 6375
rect 3893 6273 3927 6307
rect 5457 6273 5491 6307
rect 6285 6273 6319 6307
rect 7481 6273 7515 6307
rect 12449 6273 12483 6307
rect 1685 6205 1719 6239
rect 3709 6205 3743 6239
rect 5365 6205 5399 6239
rect 6101 6205 6135 6239
rect 8217 6205 8251 6239
rect 9873 6205 9907 6239
rect 10129 6205 10163 6239
rect 11805 6205 11839 6239
rect 16681 6273 16715 6307
rect 18705 6273 18739 6307
rect 19717 6273 19751 6307
rect 20729 6273 20763 6307
rect 14289 6205 14323 6239
rect 14381 6205 14415 6239
rect 16497 6205 16531 6239
rect 17417 6205 17451 6239
rect 18429 6205 18463 6239
rect 19533 6205 19567 6239
rect 1952 6137 1986 6171
rect 7205 6137 7239 6171
rect 8462 6137 8496 6171
rect 12694 6137 12728 6171
rect 13921 6137 13955 6171
rect 14648 6137 14682 6171
rect 16405 6137 16439 6171
rect 20637 6137 20671 6171
rect 3065 6069 3099 6103
rect 3801 6069 3835 6103
rect 4905 6069 4939 6103
rect 5273 6069 5307 6103
rect 5917 6069 5951 6103
rect 7297 6069 7331 6103
rect 14105 6069 14139 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 19165 6069 19199 6103
rect 19625 6069 19659 6103
rect 20545 6069 20579 6103
rect 1961 5865 1995 5899
rect 2421 5865 2455 5899
rect 2973 5865 3007 5899
rect 3433 5865 3467 5899
rect 5917 5865 5951 5899
rect 8953 5865 8987 5899
rect 11989 5865 12023 5899
rect 17509 5865 17543 5899
rect 17601 5865 17635 5899
rect 4322 5797 4356 5831
rect 12900 5797 12934 5831
rect 16396 5797 16430 5831
rect 19257 5865 19291 5899
rect 19441 5865 19475 5899
rect 18052 5797 18086 5831
rect 2329 5729 2363 5763
rect 3341 5729 3375 5763
rect 6285 5729 6319 5763
rect 7196 5729 7230 5763
rect 10057 5729 10091 5763
rect 11069 5729 11103 5763
rect 12081 5729 12115 5763
rect 12633 5729 12667 5763
rect 14289 5729 14323 5763
rect 15577 5729 15611 5763
rect 16129 5729 16163 5763
rect 17601 5729 17635 5763
rect 17785 5729 17819 5763
rect 2605 5661 2639 5695
rect 3525 5661 3559 5695
rect 4077 5661 4111 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 6929 5661 6963 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 12265 5661 12299 5695
rect 19809 5729 19843 5763
rect 19901 5661 19935 5695
rect 19993 5661 20027 5695
rect 11621 5593 11655 5627
rect 19165 5593 19199 5627
rect 19257 5593 19291 5627
rect 5457 5525 5491 5559
rect 8309 5525 8343 5559
rect 8585 5525 8619 5559
rect 9689 5525 9723 5559
rect 11253 5525 11287 5559
rect 14013 5525 14047 5559
rect 14473 5525 14507 5559
rect 15761 5525 15795 5559
rect 2053 5321 2087 5355
rect 8585 5321 8619 5355
rect 12909 5321 12943 5355
rect 14289 5321 14323 5355
rect 4721 5253 4755 5287
rect 6561 5253 6595 5287
rect 10057 5253 10091 5287
rect 18429 5253 18463 5287
rect 2605 5185 2639 5219
rect 5273 5185 5307 5219
rect 6285 5185 6319 5219
rect 2421 5117 2455 5151
rect 7481 5185 7515 5219
rect 9045 5185 9079 5219
rect 9137 5185 9171 5219
rect 10701 5185 10735 5219
rect 11713 5185 11747 5219
rect 13461 5185 13495 5219
rect 14749 5185 14783 5219
rect 14933 5185 14967 5219
rect 15301 5185 15335 5219
rect 15761 5185 15795 5219
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 8493 5117 8527 5151
rect 10425 5117 10459 5151
rect 16028 5117 16062 5151
rect 17417 5117 17451 5151
rect 5181 5049 5215 5083
rect 6561 5049 6595 5083
rect 7297 5049 7331 5083
rect 10517 5049 10551 5083
rect 11437 5049 11471 5083
rect 12449 5049 12483 5083
rect 13369 5049 13403 5083
rect 18797 5049 18831 5083
rect 19870 5049 19904 5083
rect 2513 4981 2547 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 6101 4981 6135 5015
rect 6193 4981 6227 5015
rect 6837 4981 6871 5015
rect 7205 4981 7239 5015
rect 8309 4981 8343 5015
rect 8953 4981 8987 5015
rect 11069 4981 11103 5015
rect 11529 4981 11563 5015
rect 13277 4981 13311 5015
rect 14657 4981 14691 5015
rect 17141 4981 17175 5015
rect 17601 4981 17635 5015
rect 18889 4981 18923 5015
rect 21005 4981 21039 5015
rect 3525 4777 3559 4811
rect 9689 4777 9723 4811
rect 11161 4777 11195 4811
rect 12909 4777 12943 4811
rect 16037 4777 16071 4811
rect 18245 4777 18279 4811
rect 19809 4777 19843 4811
rect 4620 4709 4654 4743
rect 6469 4709 6503 4743
rect 7665 4709 7699 4743
rect 11069 4709 11103 4743
rect 12081 4709 12115 4743
rect 12173 4709 12207 4743
rect 13544 4709 13578 4743
rect 16773 4709 16807 4743
rect 2145 4641 2179 4675
rect 2412 4641 2446 4675
rect 6377 4641 6411 4675
rect 8677 4641 8711 4675
rect 10057 4641 10091 4675
rect 12725 4641 12759 4675
rect 15301 4641 15335 4675
rect 15853 4641 15887 4675
rect 16865 4641 16899 4675
rect 17785 4641 17819 4675
rect 18674 4709 18708 4743
rect 20269 4641 20303 4675
rect 4353 4573 4387 4607
rect 6561 4573 6595 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 8769 4573 8803 4607
rect 8861 4573 8895 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11345 4573 11379 4607
rect 12357 4573 12391 4607
rect 13277 4573 13311 4607
rect 16957 4573 16991 4607
rect 17877 4573 17911 4607
rect 18061 4573 18095 4607
rect 18245 4573 18279 4607
rect 18429 4573 18463 4607
rect 7297 4505 7331 4539
rect 16405 4505 16439 4539
rect 5733 4437 5767 4471
rect 6009 4437 6043 4471
rect 8309 4437 8343 4471
rect 10701 4437 10735 4471
rect 11713 4437 11747 4471
rect 14657 4437 14691 4471
rect 15485 4437 15519 4471
rect 17417 4437 17451 4471
rect 20453 4437 20487 4471
rect 3157 4233 3191 4267
rect 4537 4233 4571 4267
rect 5457 4233 5491 4267
rect 8953 4233 8987 4267
rect 1777 4097 1811 4131
rect 3985 4097 4019 4131
rect 5089 4097 5123 4131
rect 6101 4097 6135 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 13001 4097 13035 4131
rect 13829 4097 13863 4131
rect 16497 4097 16531 4131
rect 17509 4097 17543 4131
rect 18797 4097 18831 4131
rect 19809 4097 19843 4131
rect 20821 4097 20855 4131
rect 3893 4029 3927 4063
rect 5457 4029 5491 4063
rect 6009 4029 6043 4063
rect 7021 4029 7055 4063
rect 7573 4029 7607 4063
rect 10333 4029 10367 4063
rect 12817 4029 12851 4063
rect 16221 4029 16255 4063
rect 17233 4029 17267 4063
rect 2044 3961 2078 3995
rect 5917 3961 5951 3995
rect 7840 3961 7874 3995
rect 10600 3961 10634 3995
rect 12909 3961 12943 3995
rect 14096 3961 14130 3995
rect 16313 3961 16347 3995
rect 17325 3961 17359 3995
rect 20729 3961 20763 3995
rect 3433 3893 3467 3927
rect 3801 3893 3835 3927
rect 4905 3893 4939 3927
rect 4997 3893 5031 3927
rect 5549 3893 5583 3927
rect 7205 3893 7239 3927
rect 9321 3893 9355 3927
rect 9689 3893 9723 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 15209 3893 15243 3927
rect 15853 3893 15887 3927
rect 16865 3893 16899 3927
rect 18153 3893 18187 3927
rect 18521 3893 18555 3927
rect 18613 3893 18647 3927
rect 19165 3893 19199 3927
rect 19533 3893 19567 3927
rect 19625 3893 19659 3927
rect 20269 3893 20303 3927
rect 20637 3893 20671 3927
rect 4077 3689 4111 3723
rect 7113 3689 7147 3723
rect 8769 3689 8803 3723
rect 10885 3689 10919 3723
rect 11529 3689 11563 3723
rect 11897 3689 11931 3723
rect 12357 3689 12391 3723
rect 12541 3689 12575 3723
rect 13001 3689 13035 3723
rect 13829 3689 13863 3723
rect 14565 3689 14599 3723
rect 15301 3689 15335 3723
rect 15761 3689 15795 3723
rect 17785 3689 17819 3723
rect 18613 3689 18647 3723
rect 18981 3689 19015 3723
rect 19809 3689 19843 3723
rect 10977 3621 11011 3655
rect 4445 3553 4479 3587
rect 4537 3553 4571 3587
rect 6000 3553 6034 3587
rect 7645 3553 7679 3587
rect 9045 3553 9079 3587
rect 9689 3553 9723 3587
rect 11989 3553 12023 3587
rect 4629 3485 4663 3519
rect 5273 3485 5307 3519
rect 5733 3485 5767 3519
rect 7389 3485 7423 3519
rect 9873 3485 9907 3519
rect 11069 3485 11103 3519
rect 12081 3485 12115 3519
rect 9229 3417 9263 3451
rect 20177 3621 20211 3655
rect 20269 3621 20303 3655
rect 12909 3553 12943 3587
rect 13645 3553 13679 3587
rect 15669 3553 15703 3587
rect 16405 3553 16439 3587
rect 16672 3553 16706 3587
rect 18061 3553 18095 3587
rect 20913 3553 20947 3587
rect 13093 3485 13127 3519
rect 14657 3485 14691 3519
rect 14841 3485 14875 3519
rect 15853 3485 15887 3519
rect 19073 3485 19107 3519
rect 19165 3485 19199 3519
rect 20453 3485 20487 3519
rect 10517 3349 10551 3383
rect 12357 3349 12391 3383
rect 14197 3349 14231 3383
rect 18245 3349 18279 3383
rect 4905 3145 4939 3179
rect 5181 3145 5215 3179
rect 6377 3145 6411 3179
rect 6653 3145 6687 3179
rect 6929 3145 6963 3179
rect 7941 3145 7975 3179
rect 10333 3145 10367 3179
rect 13001 3145 13035 3179
rect 14013 3145 14047 3179
rect 16957 3145 16991 3179
rect 3525 3009 3559 3043
rect 5733 3009 5767 3043
rect 5641 2941 5675 2975
rect 6193 2941 6227 2975
rect 7573 3009 7607 3043
rect 8585 3009 8619 3043
rect 10609 3009 10643 3043
rect 7297 2941 7331 2975
rect 7389 2941 7423 2975
rect 8309 2941 8343 2975
rect 8953 2941 8987 2975
rect 10876 2941 10910 2975
rect 12449 2941 12483 2975
rect 19441 3077 19475 3111
rect 14657 3009 14691 3043
rect 15577 3009 15611 3043
rect 16313 3009 16347 3043
rect 17417 3009 17451 3043
rect 17601 3009 17635 3043
rect 18061 3009 18095 3043
rect 20453 3009 20487 3043
rect 13185 2941 13219 2975
rect 14473 2941 14507 2975
rect 15393 2941 15427 2975
rect 16129 2941 16163 2975
rect 17325 2941 17359 2975
rect 18328 2941 18362 2975
rect 20269 2941 20303 2975
rect 3792 2873 3826 2907
rect 6653 2873 6687 2907
rect 9220 2873 9254 2907
rect 12725 2873 12759 2907
rect 13001 2873 13035 2907
rect 13461 2873 13495 2907
rect 3065 2805 3099 2839
rect 5549 2805 5583 2839
rect 8401 2805 8435 2839
rect 11989 2805 12023 2839
rect 14381 2805 14415 2839
rect 4077 2601 4111 2635
rect 4445 2601 4479 2635
rect 6285 2601 6319 2635
rect 6929 2601 6963 2635
rect 8217 2601 8251 2635
rect 8677 2601 8711 2635
rect 10885 2601 10919 2635
rect 11345 2601 11379 2635
rect 12173 2601 12207 2635
rect 16221 2601 16255 2635
rect 17693 2601 17727 2635
rect 18613 2601 18647 2635
rect 18981 2601 19015 2635
rect 4537 2533 4571 2567
rect 6193 2533 6227 2567
rect 7389 2533 7423 2567
rect 11253 2533 11287 2567
rect 13369 2533 13403 2567
rect 15761 2533 15795 2567
rect 17601 2533 17635 2567
rect 19073 2533 19107 2567
rect 19901 2533 19935 2567
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 9781 2465 9815 2499
rect 10057 2465 10091 2499
rect 11989 2465 12023 2499
rect 13093 2465 13127 2499
rect 13829 2465 13863 2499
rect 14105 2465 14139 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16681 2465 16715 2499
rect 19625 2465 19659 2499
rect 20545 2465 20579 2499
rect 4629 2397 4663 2431
rect 6469 2397 6503 2431
rect 7573 2397 7607 2431
rect 8861 2397 8895 2431
rect 11437 2397 11471 2431
rect 17877 2397 17911 2431
rect 19165 2397 19199 2431
rect 5825 2329 5859 2363
rect 16865 2329 16899 2363
rect 15025 2261 15059 2295
rect 17233 2261 17267 2295
rect 20729 2261 20763 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3878 19456 3884 19508
rect 3936 19496 3942 19508
rect 5813 19499 5871 19505
rect 5813 19496 5825 19499
rect 3936 19468 5825 19496
rect 3936 19456 3942 19468
rect 5813 19465 5825 19468
rect 5859 19465 5871 19499
rect 19150 19496 19156 19508
rect 19111 19468 19156 19496
rect 5813 19459 5871 19465
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 4982 19292 4988 19304
rect 2363 19264 4988 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 1780 19224 1808 19255
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5626 19292 5632 19304
rect 5587 19264 5632 19292
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 18414 19252 18420 19304
rect 18472 19292 18478 19304
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18472 19264 18981 19292
rect 18472 19252 18478 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 18969 19255 19027 19261
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 19760 19264 20545 19292
rect 19760 19252 19766 19264
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 6086 19224 6092 19236
rect 1780 19196 6092 19224
rect 6086 19184 6092 19196
rect 6144 19184 6150 19236
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 5626 18844 5632 18896
rect 5684 18884 5690 18896
rect 6273 18887 6331 18893
rect 6273 18884 6285 18887
rect 5684 18856 6285 18884
rect 5684 18844 5690 18856
rect 6273 18853 6285 18856
rect 6319 18853 6331 18887
rect 18414 18884 18420 18896
rect 18375 18856 18420 18884
rect 6273 18847 6331 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 1486 18776 1492 18828
rect 1544 18816 1550 18828
rect 1765 18819 1823 18825
rect 1765 18816 1777 18819
rect 1544 18788 1777 18816
rect 1544 18776 1550 18788
rect 1765 18785 1777 18788
rect 1811 18785 1823 18819
rect 5994 18816 6000 18828
rect 5955 18788 6000 18816
rect 1765 18779 1823 18785
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18816 18199 18819
rect 19610 18816 19616 18828
rect 18187 18788 19616 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 19610 18776 19616 18788
rect 19668 18776 19674 18828
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 8202 18204 8208 18216
rect 5776 18176 8208 18204
rect 5776 18164 5782 18176
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 20530 18204 20536 18216
rect 20491 18176 20536 18204
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2409 17799 2467 17805
rect 2409 17796 2421 17799
rect 1820 17768 2421 17796
rect 1820 17756 1826 17768
rect 2409 17765 2421 17768
rect 2455 17765 2467 17799
rect 2409 17759 2467 17765
rect 19889 17799 19947 17805
rect 19889 17765 19901 17799
rect 19935 17796 19947 17799
rect 20530 17796 20536 17808
rect 19935 17768 20536 17796
rect 19935 17765 19947 17768
rect 19889 17759 19947 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 6730 17728 6736 17740
rect 2179 17700 6736 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 1596 17660 1624 17691
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 20254 17728 20260 17740
rect 19659 17700 20260 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 7374 17660 7380 17672
rect 1596 17632 7380 17660
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 1728 17564 1777 17592
rect 1728 17552 1734 17564
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 1765 17555 1823 17561
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 7098 17116 7104 17128
rect 1811 17088 7104 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 20530 17116 20536 17128
rect 20491 17088 20536 17116
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1912 16748 1961 16776
rect 1912 16736 1918 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 20438 16776 20444 16788
rect 20399 16748 20444 16776
rect 1949 16739 2007 16745
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 4890 16640 4896 16652
rect 1811 16612 4896 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20622 16640 20628 16652
rect 20303 16612 20628 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 3326 16232 3332 16244
rect 3287 16204 3332 16232
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 17862 16232 17868 16244
rect 13587 16204 17868 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20806 16232 20812 16244
rect 20763 16204 20812 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 7466 16096 7472 16108
rect 2332 16068 7472 16096
rect 2332 16037 2360 16068
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 2323 16031 2381 16037
rect 2323 15997 2335 16031
rect 2369 15997 2381 16031
rect 3142 16028 3148 16040
rect 3103 16000 3148 16028
rect 2323 15991 2381 15997
rect 1780 15960 1808 15991
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 12860 16000 13369 16028
rect 12860 15988 12866 16000
rect 13357 15997 13369 16000
rect 13403 15997 13415 16031
rect 13357 15991 13415 15997
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19392 16000 19993 16028
rect 19392 15988 19398 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 20162 15988 20168 16040
rect 20220 16028 20226 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20220 16000 20545 16028
rect 20220 15988 20226 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 4706 15960 4712 15972
rect 1780 15932 4712 15960
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2464 15660 2513 15688
rect 2464 15648 2470 15660
rect 2501 15657 2513 15660
rect 2547 15657 2559 15691
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 2501 15651 2559 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 3142 15580 3148 15632
rect 3200 15620 3206 15632
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 3200 15592 4353 15620
rect 3200 15580 3206 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 12802 15620 12808 15632
rect 12763 15592 12808 15620
rect 4341 15583 4399 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 2323 15555 2381 15561
rect 2323 15521 2335 15555
rect 2369 15521 2381 15555
rect 2323 15515 2381 15521
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4246 15552 4252 15564
rect 4111 15524 4252 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 1780 15416 1808 15515
rect 2332 15484 2360 15515
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 5074 15484 5080 15496
rect 2332 15456 5080 15484
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 19720 15484 19748 15515
rect 19978 15512 19984 15564
rect 20036 15552 20042 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 20036 15524 20269 15552
rect 20036 15512 20042 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20806 15484 20812 15496
rect 19720 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 5166 15416 5172 15428
rect 1780 15388 5172 15416
rect 5166 15376 5172 15388
rect 5224 15376 5230 15428
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2774 15144 2780 15156
rect 2547 15116 2780 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 20070 15104 20076 15156
rect 20128 15144 20134 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 20128 15116 20177 15144
rect 20128 15104 20134 15116
rect 20165 15113 20177 15116
rect 20211 15113 20223 15147
rect 20165 15107 20223 15113
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20717 15147 20775 15153
rect 20717 15144 20729 15147
rect 20404 15116 20729 15144
rect 20404 15104 20410 15116
rect 20717 15113 20729 15116
rect 20763 15113 20775 15147
rect 20717 15107 20775 15113
rect 1946 15076 1952 15088
rect 1907 15048 1952 15076
rect 1946 15036 1952 15048
rect 2004 15036 2010 15088
rect 19610 15076 19616 15088
rect 19571 15048 19616 15076
rect 19610 15036 19616 15048
rect 19668 15036 19674 15088
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2464 14980 2973 15008
rect 2464 14968 2470 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 16390 14968 16396 15020
rect 16448 15008 16454 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16448 14980 16773 15008
rect 16448 14968 16454 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 17552 14980 20024 15008
rect 17552 14968 17558 14980
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2323 14943 2381 14949
rect 2323 14909 2335 14943
rect 2369 14909 2381 14943
rect 5902 14940 5908 14952
rect 2323 14903 2381 14909
rect 3160 14912 5908 14940
rect 2332 14872 2360 14903
rect 3160 14872 3188 14912
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19996 14949 20024 14980
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 2332 14844 3188 14872
rect 3228 14875 3286 14881
rect 3228 14841 3240 14875
rect 3274 14872 3286 14875
rect 3786 14872 3792 14884
rect 3274 14844 3792 14872
rect 3274 14841 3286 14844
rect 3228 14835 3286 14841
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 12768 14844 16681 14872
rect 12768 14832 12774 14844
rect 16669 14841 16681 14844
rect 16715 14872 16727 14875
rect 20548 14872 20576 14903
rect 16715 14844 20576 14872
rect 16715 14841 16727 14844
rect 16669 14835 16727 14841
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4212 14776 4353 14804
rect 4212 14764 4218 14776
rect 4341 14773 4353 14776
rect 4387 14773 4399 14807
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 4341 14767 4399 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16574 14804 16580 14816
rect 16535 14776 16580 14804
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3476 14572 4261 14600
rect 3476 14560 3482 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 17126 14600 17132 14612
rect 11756 14572 17132 14600
rect 11756 14560 11762 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 19334 14600 19340 14612
rect 19295 14572 19340 14600
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2317 14535 2375 14541
rect 2317 14532 2329 14535
rect 1820 14504 2329 14532
rect 1820 14492 1826 14504
rect 2317 14501 2329 14504
rect 2363 14501 2375 14535
rect 2317 14495 2375 14501
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14532 7619 14535
rect 7742 14532 7748 14544
rect 7607 14504 7748 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 11808 14504 12204 14532
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14464 1547 14467
rect 1854 14464 1860 14476
rect 1535 14436 1860 14464
rect 1535 14433 1547 14436
rect 1489 14427 1547 14433
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1995 14436 2053 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3237 14467 3295 14473
rect 3237 14464 3249 14467
rect 2924 14436 3249 14464
rect 2924 14424 2930 14436
rect 3237 14433 3249 14436
rect 3283 14433 3295 14467
rect 3237 14427 3295 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 5350 14464 5356 14476
rect 4111 14436 5356 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 11808 14473 11836 14504
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 9916 14436 10425 14464
rect 9916 14424 9922 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14433 11851 14467
rect 12049 14467 12107 14473
rect 12049 14464 12061 14467
rect 11793 14427 11851 14433
rect 11900 14436 12061 14464
rect 3326 14396 3332 14408
rect 3287 14368 3332 14396
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14396 3571 14399
rect 4154 14396 4160 14408
rect 3559 14368 4160 14396
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 7650 14396 7656 14408
rect 7611 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 10502 14396 10508 14408
rect 10463 14368 10508 14396
rect 7745 14359 7803 14365
rect 7558 14288 7564 14340
rect 7616 14328 7622 14340
rect 7760 14328 7788 14359
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 11146 14396 11152 14408
rect 10735 14368 11152 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 11900 14396 11928 14436
rect 12049 14433 12061 14436
rect 12095 14433 12107 14467
rect 12176 14464 12204 14504
rect 13096 14504 19288 14532
rect 12434 14464 12440 14476
rect 12176 14436 12440 14464
rect 12049 14427 12107 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 11808 14368 11928 14396
rect 7616 14300 7788 14328
rect 7616 14288 7622 14300
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 11808 14328 11836 14368
rect 8260 14300 11836 14328
rect 8260 14288 8266 14300
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 1995 14232 2881 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 2869 14223 2927 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 10045 14263 10103 14269
rect 10045 14229 10057 14263
rect 10091 14260 10103 14263
rect 13096 14260 13124 14504
rect 14274 14464 14280 14476
rect 14235 14436 14280 14464
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 14369 14467 14427 14473
rect 14369 14433 14381 14467
rect 14415 14464 14427 14467
rect 15286 14464 15292 14476
rect 14415 14436 15292 14464
rect 14415 14433 14427 14436
rect 14369 14427 14427 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 16016 14467 16074 14473
rect 16016 14433 16028 14467
rect 16062 14464 16074 14467
rect 16390 14464 16396 14476
rect 16062 14436 16396 14464
rect 16062 14433 16074 14436
rect 16016 14427 16074 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 18598 14464 18604 14476
rect 18559 14436 18604 14464
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 18748 14436 19165 14464
rect 18748 14424 18754 14436
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 19260 14464 19288 14504
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19981 14535 20039 14541
rect 19981 14532 19993 14535
rect 19484 14504 19993 14532
rect 19484 14492 19490 14504
rect 19981 14501 19993 14504
rect 20027 14501 20039 14535
rect 19981 14495 20039 14501
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 19260 14436 19717 14464
rect 19153 14427 19211 14433
rect 19705 14433 19717 14436
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 14734 14396 14740 14408
rect 14599 14368 14740 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15562 14396 15568 14408
rect 15068 14368 15568 14396
rect 15068 14356 15074 14368
rect 15562 14356 15568 14368
rect 15620 14396 15626 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15620 14368 15761 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 20530 14396 20536 14408
rect 15749 14359 15807 14365
rect 16960 14368 20536 14396
rect 10091 14232 13124 14260
rect 13173 14263 13231 14269
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 13173 14229 13185 14263
rect 13219 14260 13231 14263
rect 13538 14260 13544 14272
rect 13219 14232 13544 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 13909 14263 13967 14269
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 15194 14260 15200 14272
rect 13955 14232 15200 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 16960 14260 16988 14368
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 20622 14328 20628 14340
rect 17092 14300 20628 14328
rect 17092 14288 17098 14300
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 17126 14260 17132 14272
rect 16172 14232 16988 14260
rect 17087 14232 17132 14260
rect 16172 14220 16178 14232
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 18785 14263 18843 14269
rect 18785 14229 18797 14263
rect 18831 14260 18843 14263
rect 18874 14260 18880 14272
rect 18831 14232 18880 14260
rect 18831 14229 18843 14232
rect 18785 14223 18843 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 2464 14028 4016 14056
rect 2464 14016 2470 14028
rect 2130 13920 2136 13932
rect 1688 13892 2136 13920
rect 1688 13861 1716 13892
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2406 13920 2412 13932
rect 2367 13892 2412 13920
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 3988 13920 4016 14028
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 11204 14028 11437 14056
rect 11204 14016 11210 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 11425 14019 11483 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 19242 14056 19248 14068
rect 16132 14028 19248 14056
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 5316 13960 5457 13988
rect 5316 13948 5322 13960
rect 5445 13957 5457 13960
rect 5491 13957 5503 13991
rect 5445 13951 5503 13957
rect 7282 13948 7288 14000
rect 7340 13988 7346 14000
rect 9766 13988 9772 14000
rect 7340 13960 7420 13988
rect 9727 13960 9772 13988
rect 7340 13948 7346 13960
rect 4062 13920 4068 13932
rect 3975 13892 4068 13920
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13821 1731 13855
rect 1673 13815 1731 13821
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 3234 13852 3240 13864
rect 1995 13824 3240 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4321 13855 4379 13861
rect 4321 13852 4333 13855
rect 4212 13824 4333 13852
rect 4212 13812 4218 13824
rect 4321 13821 4333 13824
rect 4367 13821 4379 13855
rect 4321 13815 4379 13821
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 4856 13824 7297 13852
rect 4856 13812 4862 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7392 13852 7420 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 9784 13920 9812 13948
rect 14752 13920 14780 14016
rect 9784 13892 10180 13920
rect 14752 13892 15148 13920
rect 10152 13864 10180 13892
rect 8662 13861 8668 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 7392 13824 8401 13852
rect 7285 13815 7343 13821
rect 8389 13821 8401 13824
rect 8435 13852 8447 13855
rect 8656 13852 8668 13861
rect 8435 13824 8524 13852
rect 8623 13824 8668 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8496 13796 8524 13824
rect 8656 13815 8668 13824
rect 8662 13812 8668 13815
rect 8720 13812 8726 13864
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 8772 13824 10057 13852
rect 2676 13787 2734 13793
rect 2676 13753 2688 13787
rect 2722 13784 2734 13787
rect 3142 13784 3148 13796
rect 2722 13756 3148 13784
rect 2722 13753 2734 13756
rect 2676 13747 2734 13753
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 7193 13787 7251 13793
rect 5132 13756 6960 13784
rect 5132 13744 5138 13756
rect 3786 13716 3792 13728
rect 3747 13688 3792 13716
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 6932 13716 6960 13756
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7239 13756 7849 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 8772 13784 8800 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10134 13812 10140 13864
rect 10192 13852 10198 13864
rect 10301 13855 10359 13861
rect 10301 13852 10313 13855
rect 10192 13824 10313 13852
rect 10192 13812 10198 13824
rect 10301 13821 10313 13824
rect 10347 13821 10359 13855
rect 12434 13852 12440 13864
rect 10301 13815 10359 13821
rect 11072 13824 12440 13852
rect 8536 13756 8800 13784
rect 8536 13744 8542 13756
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 11072 13784 11100 13824
rect 12434 13812 12440 13824
rect 12492 13852 12498 13864
rect 13078 13852 13084 13864
rect 12492 13824 13084 13852
rect 12492 13812 12498 13824
rect 13078 13812 13084 13824
rect 13136 13852 13142 13864
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 13136 13824 13369 13852
rect 13136 13812 13142 13824
rect 13357 13821 13369 13824
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 13624 13855 13682 13861
rect 13624 13821 13636 13855
rect 13670 13852 13682 13855
rect 14458 13852 14464 13864
rect 13670 13824 14464 13852
rect 13670 13821 13682 13824
rect 13624 13815 13682 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15010 13852 15016 13864
rect 14971 13824 15016 13852
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15120 13852 15148 13892
rect 15269 13855 15327 13861
rect 15269 13852 15281 13855
rect 15120 13824 15281 13852
rect 15269 13821 15281 13824
rect 15315 13821 15327 13855
rect 15269 13815 15327 13821
rect 11020 13756 11100 13784
rect 11020 13744 11026 13756
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 16132 13784 16160 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 16669 13991 16727 13997
rect 16669 13957 16681 13991
rect 16715 13988 16727 13991
rect 16715 13960 18092 13988
rect 16715 13957 16727 13960
rect 16669 13951 16727 13957
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17184 13892 17233 13920
rect 17184 13880 17190 13892
rect 17221 13889 17233 13892
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 18064 13861 18092 13960
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 19702 13988 19708 14000
rect 19392 13960 19708 13988
rect 19392 13948 19398 13960
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 18598 13880 18604 13932
rect 18656 13920 18662 13932
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 18656 13892 20085 13920
rect 18656 13880 18662 13892
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20806 13920 20812 13932
rect 20767 13892 20812 13920
rect 20073 13883 20131 13889
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 17037 13855 17095 13861
rect 17037 13852 17049 13855
rect 16264 13824 17049 13852
rect 16264 13812 16270 13824
rect 17037 13821 17049 13824
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18782 13852 18788 13864
rect 18743 13824 18788 13852
rect 18049 13815 18107 13821
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19889 13855 19947 13861
rect 19889 13852 19901 13855
rect 19576 13824 19901 13852
rect 19576 13812 19582 13824
rect 19889 13821 19901 13824
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 11296 13756 16160 13784
rect 11296 13744 11302 13756
rect 16850 13744 16856 13796
rect 16908 13784 16914 13796
rect 17129 13787 17187 13793
rect 17129 13784 17141 13787
rect 16908 13756 17141 13784
rect 16908 13744 16914 13756
rect 17129 13753 17141 13756
rect 17175 13753 17187 13787
rect 17129 13747 17187 13753
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 18325 13787 18383 13793
rect 18325 13784 18337 13787
rect 17276 13756 18337 13784
rect 17276 13744 17282 13756
rect 18325 13753 18337 13756
rect 18371 13753 18383 13787
rect 18325 13747 18383 13753
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18656 13756 19073 13784
rect 18656 13744 18662 13756
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 19702 13744 19708 13796
rect 19760 13784 19766 13796
rect 20640 13784 20668 13815
rect 19760 13756 20668 13784
rect 19760 13744 19766 13756
rect 15746 13716 15752 13728
rect 6932 13688 15752 13716
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 16390 13716 16396 13728
rect 16303 13688 16396 13716
rect 16390 13676 16396 13688
rect 16448 13716 16454 13728
rect 17402 13716 17408 13728
rect 16448 13688 17408 13716
rect 16448 13676 16454 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2866 13512 2872 13524
rect 1995 13484 2872 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 3326 13512 3332 13524
rect 3007 13484 3332 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 3568 13484 4261 13512
rect 3568 13472 3574 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 4249 13475 4307 13481
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6052 13484 6285 13512
rect 6052 13472 6058 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 6822 13512 6828 13524
rect 6687 13484 6828 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8404 13484 8677 13512
rect 6733 13447 6791 13453
rect 6733 13413 6745 13447
rect 6779 13444 6791 13447
rect 7190 13444 7196 13456
rect 6779 13416 7196 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 8404 13444 8432 13484
rect 8665 13481 8677 13484
rect 8711 13512 8723 13515
rect 11698 13512 11704 13524
rect 8711 13484 11704 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 14458 13512 14464 13524
rect 14419 13484 14464 13512
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16574 13512 16580 13524
rect 16439 13484 16580 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 20441 13515 20499 13521
rect 20441 13512 20453 13515
rect 19852 13484 20453 13512
rect 19852 13472 19858 13484
rect 20441 13481 20453 13484
rect 20487 13481 20499 13515
rect 20441 13475 20499 13481
rect 7392 13416 8432 13444
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 3878 13376 3884 13388
rect 3375 13348 3884 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 7282 13376 7288 13388
rect 7243 13348 7288 13376
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2498 13308 2504 13320
rect 2455 13280 2504 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 3418 13308 3424 13320
rect 3379 13280 3424 13308
rect 2593 13271 2651 13277
rect 2608 13240 2636 13271
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 3786 13308 3792 13320
rect 3559 13280 3792 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 3528 13240 3556 13271
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 4764 13280 5181 13308
rect 4764 13268 4770 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 2608 13212 3556 13240
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 5184 13240 5212 13271
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7392 13308 7420 13416
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10410 13444 10416 13456
rect 10008 13416 10416 13444
rect 10008 13404 10014 13416
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 11054 13444 11060 13456
rect 10520 13416 11060 13444
rect 7558 13385 7564 13388
rect 7552 13339 7564 13385
rect 7616 13376 7622 13388
rect 7616 13348 7652 13376
rect 7558 13336 7564 13339
rect 7616 13336 7622 13348
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 10321 13379 10379 13385
rect 7892 13348 10272 13376
rect 7892 13336 7898 13348
rect 6963 13280 7420 13308
rect 9125 13311 9183 13317
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 10134 13308 10140 13320
rect 9171 13280 10140 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10244 13308 10272 13348
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10520 13376 10548 13416
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 11146 13404 11152 13456
rect 11204 13453 11210 13456
rect 11204 13447 11268 13453
rect 11204 13413 11222 13447
rect 11256 13413 11268 13447
rect 11204 13407 11268 13413
rect 11204 13404 11210 13407
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 15620 13416 16344 13444
rect 15620 13404 15626 13416
rect 16316 13388 16344 13416
rect 17126 13404 17132 13456
rect 17184 13453 17190 13456
rect 17184 13447 17248 13453
rect 17184 13413 17202 13447
rect 17236 13413 17248 13447
rect 18506 13444 18512 13456
rect 17184 13407 17248 13413
rect 17328 13416 18512 13444
rect 17184 13404 17190 13407
rect 13078 13376 13084 13388
rect 10367 13348 10548 13376
rect 10612 13348 12940 13376
rect 13039 13348 13084 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10612 13317 10640 13348
rect 10597 13311 10655 13317
rect 10244 13280 10548 13308
rect 7190 13240 7196 13252
rect 4028 13212 4844 13240
rect 5184 13212 7196 13240
rect 4028 13200 4034 13212
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4816 13172 4844 13212
rect 7190 13200 7196 13212
rect 7248 13200 7254 13252
rect 10520 13240 10548 13280
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10686 13308 10692 13320
rect 10643 13280 10692 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10962 13308 10968 13320
rect 10923 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13308 12679 13311
rect 12802 13308 12808 13320
rect 12667 13280 12808 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 12912 13308 12940 13348
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13348 13379 13406 13385
rect 13348 13345 13360 13379
rect 13394 13376 13406 13379
rect 15102 13376 15108 13388
rect 13394 13348 15108 13376
rect 13394 13345 13406 13348
rect 13348 13339 13406 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15436 13348 15669 13376
rect 15436 13336 15442 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16356 13348 16957 13376
rect 16356 13336 16362 13348
rect 16945 13345 16957 13348
rect 16991 13376 17003 13379
rect 17328 13376 17356 13416
rect 18506 13404 18512 13416
rect 18564 13404 18570 13456
rect 18868 13379 18926 13385
rect 18868 13376 18880 13379
rect 16991 13348 17356 13376
rect 18340 13348 18880 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 14734 13308 14740 13320
rect 12912 13280 13124 13308
rect 14695 13280 14740 13308
rect 10778 13240 10784 13252
rect 8220 13212 10456 13240
rect 10520 13212 10784 13240
rect 8220 13172 8248 13212
rect 4816 13144 8248 13172
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10318 13172 10324 13184
rect 9999 13144 10324 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10428 13172 10456 13212
rect 10778 13200 10784 13212
rect 10836 13200 10842 13252
rect 12986 13240 12992 13252
rect 11900 13212 12992 13240
rect 11900 13172 11928 13212
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 12342 13172 12348 13184
rect 10428 13144 11928 13172
rect 12303 13144 12348 13172
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 13096 13172 13124 13280
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 15856 13240 15884 13271
rect 18340 13249 18368 13348
rect 18868 13345 18880 13348
rect 18914 13376 18926 13379
rect 19978 13376 19984 13388
rect 18914 13348 19984 13376
rect 18914 13345 18926 13348
rect 18868 13339 18926 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 18506 13268 18512 13320
rect 18564 13308 18570 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 18564 13280 18613 13308
rect 18564 13268 18570 13280
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20272 13308 20300 13339
rect 19852 13280 20300 13308
rect 19852 13268 19858 13280
rect 14516 13212 15884 13240
rect 18325 13243 18383 13249
rect 14516 13200 14522 13212
rect 18325 13209 18337 13243
rect 18371 13209 18383 13243
rect 18325 13203 18383 13209
rect 16666 13172 16672 13184
rect 13096 13144 16672 13172
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 19886 13132 19892 13184
rect 19944 13172 19950 13184
rect 19981 13175 20039 13181
rect 19981 13172 19993 13175
rect 19944 13144 19993 13172
rect 19944 13132 19950 13144
rect 19981 13141 19993 13144
rect 20027 13141 20039 13175
rect 19981 13135 20039 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2498 12968 2504 12980
rect 2459 12940 2504 12968
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 3789 12971 3847 12977
rect 3789 12968 3801 12971
rect 3476 12940 3801 12968
rect 3476 12928 3482 12940
rect 3789 12937 3801 12940
rect 3835 12937 3847 12971
rect 3789 12931 3847 12937
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 3936 12940 6837 12968
rect 3936 12928 3942 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12968 9183 12971
rect 10502 12968 10508 12980
rect 9171 12940 10508 12968
rect 9171 12937 9183 12940
rect 9125 12931 9183 12937
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 10652 12940 13829 12968
rect 10652 12928 10658 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 14274 12968 14280 12980
rect 13955 12940 14280 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18782 12968 18788 12980
rect 18371 12940 18788 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 4062 12900 4068 12912
rect 2056 12872 4068 12900
rect 2056 12841 2084 12872
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 4154 12860 4160 12912
rect 4212 12900 4218 12912
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4212 12872 4629 12900
rect 4212 12860 4218 12872
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 6181 12903 6239 12909
rect 6181 12869 6193 12903
rect 6227 12869 6239 12903
rect 6181 12863 6239 12869
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 7837 12903 7895 12909
rect 6687 12872 7512 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2041 12795 2099 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 4430 12832 4436 12844
rect 4343 12804 4436 12832
rect 4430 12792 4436 12804
rect 4488 12832 4494 12844
rect 6196 12832 6224 12863
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 4488 12804 4936 12832
rect 4488 12792 4494 12804
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 3694 12764 3700 12776
rect 1811 12736 3700 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4663 12736 4813 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 4908 12764 4936 12804
rect 6196 12804 7389 12832
rect 6196 12764 6224 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7484 12832 7512 12872
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 8662 12900 8668 12912
rect 7883 12872 8432 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7484 12804 8309 12832
rect 7377 12795 7435 12801
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 4908 12736 6224 12764
rect 4801 12727 4859 12733
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 8404 12764 8432 12872
rect 8496 12872 8668 12900
rect 8496 12841 8524 12872
rect 8662 12860 8668 12872
rect 8720 12900 8726 12912
rect 8720 12872 10732 12900
rect 8720 12860 8726 12872
rect 10704 12844 10732 12872
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 12158 12900 12164 12912
rect 10836 12872 12164 12900
rect 10836 12860 10842 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 12437 12903 12495 12909
rect 12437 12869 12449 12903
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 10042 12832 10048 12844
rect 9815 12804 10048 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10502 12832 10508 12844
rect 10192 12804 10508 12832
rect 10192 12792 10198 12804
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10686 12832 10692 12844
rect 10647 12804 10692 12832
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 11882 12832 11888 12844
rect 11843 12804 11888 12832
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12452 12832 12480 12863
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 20254 12900 20260 12912
rect 15988 12872 20260 12900
rect 15988 12860 15994 12872
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 12032 12804 12480 12832
rect 12032 12792 12038 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12768 12804 12909 12832
rect 12768 12792 12774 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 12989 12795 13047 12801
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 7064 12736 7328 12764
rect 8404 12736 9505 12764
rect 7064 12724 7070 12736
rect 2869 12699 2927 12705
rect 2869 12665 2881 12699
rect 2915 12696 2927 12699
rect 3050 12696 3056 12708
rect 2915 12668 3056 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4706 12696 4712 12708
rect 4203 12668 4712 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4706 12656 4712 12668
rect 4764 12696 4770 12708
rect 5068 12699 5126 12705
rect 4764 12668 5028 12696
rect 4764 12656 4770 12668
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3786 12628 3792 12640
rect 3016 12600 3792 12628
rect 3016 12588 3022 12600
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 4614 12628 4620 12640
rect 4295 12600 4620 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5000 12628 5028 12668
rect 5068 12665 5080 12699
rect 5114 12696 5126 12699
rect 5442 12696 5448 12708
rect 5114 12668 5448 12696
rect 5114 12665 5126 12668
rect 5068 12659 5126 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7300 12705 7328 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 13004 12764 13032 12795
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 16080 12804 16313 12832
rect 16080 12792 16086 12804
rect 16301 12801 16313 12804
rect 16347 12832 16359 12835
rect 16390 12832 16396 12844
rect 16347 12804 16396 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16850 12832 16856 12844
rect 16531 12804 16856 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17402 12832 17408 12844
rect 17363 12804 17408 12832
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19886 12832 19892 12844
rect 19847 12804 19892 12832
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 19978 12792 19984 12844
rect 20036 12832 20042 12844
rect 20901 12835 20959 12841
rect 20901 12832 20913 12835
rect 20036 12804 20913 12832
rect 20036 12792 20042 12804
rect 20901 12801 20913 12804
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 12400 12736 13032 12764
rect 14277 12767 14335 12773
rect 12400 12724 12406 12736
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 14734 12764 14740 12776
rect 14323 12736 14740 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 20806 12764 20812 12776
rect 15620 12736 20812 12764
rect 15620 12724 15626 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 8205 12699 8263 12705
rect 8205 12696 8217 12699
rect 7331 12668 8217 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 8205 12665 8217 12668
rect 8251 12665 8263 12699
rect 8205 12659 8263 12665
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10502 12696 10508 12708
rect 9640 12668 10272 12696
rect 10463 12668 10508 12696
rect 9640 12656 9646 12668
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 5000 12600 6653 12628
rect 6641 12597 6653 12600
rect 6687 12597 6699 12631
rect 6641 12591 6699 12597
rect 7193 12631 7251 12637
rect 7193 12597 7205 12631
rect 7239 12628 7251 12631
rect 9950 12628 9956 12640
rect 7239 12600 9956 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10134 12628 10140 12640
rect 10095 12600 10140 12628
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10244 12628 10272 12668
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 11698 12696 11704 12708
rect 11659 12668 11704 12696
rect 11698 12656 11704 12668
rect 11756 12656 11762 12708
rect 12802 12696 12808 12708
rect 12763 12668 12808 12696
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12696 14427 12699
rect 17494 12696 17500 12708
rect 14415 12668 17500 12696
rect 14415 12665 14427 12668
rect 14369 12659 14427 12665
rect 10594 12628 10600 12640
rect 10244 12600 10600 12628
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 11333 12631 11391 12637
rect 11333 12597 11345 12631
rect 11379 12628 11391 12631
rect 11606 12628 11612 12640
rect 11379 12600 11612 12628
rect 11379 12597 11391 12600
rect 11333 12591 11391 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12066 12628 12072 12640
rect 11839 12600 12072 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14384 12628 14412 12659
rect 17494 12656 17500 12668
rect 17552 12656 17558 12708
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12696 18751 12699
rect 19705 12699 19763 12705
rect 18739 12668 19380 12696
rect 18739 12665 18751 12668
rect 18693 12659 18751 12665
rect 15838 12628 15844 12640
rect 13863 12600 14412 12628
rect 15799 12600 15844 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 16540 12600 17233 12628
rect 16540 12588 16546 12600
rect 17221 12597 17233 12600
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 17586 12628 17592 12640
rect 17359 12600 17592 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 18782 12628 18788 12640
rect 18743 12600 18788 12628
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 19352 12637 19380 12668
rect 19705 12665 19717 12699
rect 19751 12696 19763 12699
rect 20530 12696 20536 12708
rect 19751 12668 20536 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 20530 12656 20536 12668
rect 20588 12656 20594 12708
rect 20714 12696 20720 12708
rect 20675 12668 20720 12696
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12597 19395 12631
rect 19794 12628 19800 12640
rect 19755 12600 19800 12628
rect 19337 12591 19395 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 20346 12628 20352 12640
rect 20307 12600 20352 12628
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2372 12396 2421 12424
rect 2372 12384 2378 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 3602 12424 3608 12436
rect 3563 12396 3608 12424
rect 2409 12387 2467 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 7558 12424 7564 12436
rect 7515 12396 7564 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 7800 12396 8125 12424
rect 7800 12384 7806 12396
rect 8113 12393 8125 12396
rect 8159 12393 8171 12427
rect 8113 12387 8171 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9306 12424 9312 12436
rect 8619 12396 9312 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9858 12424 9864 12436
rect 9819 12396 9864 12424
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10318 12424 10324 12436
rect 10279 12396 10324 12424
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 12802 12424 12808 12436
rect 10428 12396 12808 12424
rect 1394 12316 1400 12368
rect 1452 12356 1458 12368
rect 1949 12359 2007 12365
rect 1949 12356 1961 12359
rect 1452 12328 1961 12356
rect 1452 12316 1458 12328
rect 1949 12325 1961 12328
rect 1995 12325 2007 12359
rect 1949 12319 2007 12325
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 4028 12328 8616 12356
rect 4028 12316 4034 12328
rect 1670 12288 1676 12300
rect 1631 12260 1676 12288
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 3234 12248 3240 12300
rect 3292 12288 3298 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3292 12260 3433 12288
rect 3292 12248 3298 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 4321 12291 4379 12297
rect 4321 12288 4333 12291
rect 3568 12260 4333 12288
rect 3568 12248 3574 12260
rect 4321 12257 4333 12260
rect 4367 12257 4379 12291
rect 4321 12251 4379 12257
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5442 12288 5448 12300
rect 4948 12260 5448 12288
rect 4948 12248 4954 12260
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6356 12291 6414 12297
rect 6356 12257 6368 12291
rect 6402 12288 6414 12291
rect 6914 12288 6920 12300
rect 6402 12260 6920 12288
rect 6402 12257 6414 12260
rect 6356 12251 6414 12257
rect 6914 12248 6920 12260
rect 6972 12288 6978 12300
rect 8018 12288 8024 12300
rect 6972 12260 8024 12288
rect 6972 12248 6978 12260
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12257 8539 12291
rect 8588 12288 8616 12328
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 10192 12328 10241 12356
rect 10192 12316 10198 12328
rect 10229 12325 10241 12328
rect 10275 12325 10287 12359
rect 10229 12319 10287 12325
rect 10428 12288 10456 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 12986 12424 12992 12436
rect 12947 12396 12992 12424
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 15896 12396 17601 12424
rect 15896 12384 15902 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 17589 12387 17647 12393
rect 18506 12384 18512 12436
rect 18564 12384 18570 12436
rect 18966 12384 18972 12436
rect 19024 12424 19030 12436
rect 19334 12424 19340 12436
rect 19024 12396 19340 12424
rect 19024 12384 19030 12396
rect 19334 12384 19340 12396
rect 19392 12424 19398 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19392 12396 19717 12424
rect 19392 12384 19398 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 20530 12384 20536 12436
rect 20588 12424 20594 12436
rect 20901 12427 20959 12433
rect 20901 12424 20913 12427
rect 20588 12396 20913 12424
rect 20588 12384 20594 12396
rect 20901 12393 20913 12396
rect 20947 12393 20959 12427
rect 20901 12387 20959 12393
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 17494 12356 17500 12368
rect 10652 12328 17500 12356
rect 10652 12316 10658 12328
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 8588 12260 10456 12288
rect 10873 12291 10931 12297
rect 8481 12251 8539 12257
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 10962 12288 10968 12300
rect 10919 12260 10968 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3142 12220 3148 12232
rect 3099 12192 3148 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 2884 12152 2912 12183
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 4062 12220 4068 12232
rect 4023 12192 4068 12220
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 6052 12192 6101 12220
rect 6052 12180 6058 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 8496 12220 8524 12251
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11140 12291 11198 12297
rect 11140 12257 11152 12291
rect 11186 12288 11198 12291
rect 11882 12288 11888 12300
rect 11186 12260 11888 12288
rect 11186 12257 11198 12260
rect 11140 12251 11198 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 12943 12260 13553 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 15832 12291 15890 12297
rect 15832 12288 15844 12291
rect 15712 12260 15844 12288
rect 15712 12248 15718 12260
rect 15832 12257 15844 12260
rect 15878 12288 15890 12291
rect 18325 12291 18383 12297
rect 15878 12260 17908 12288
rect 15878 12257 15890 12260
rect 15832 12251 15890 12257
rect 17880 12232 17908 12260
rect 18325 12257 18337 12291
rect 18371 12288 18383 12291
rect 18524 12288 18552 12384
rect 18592 12359 18650 12365
rect 18592 12325 18604 12359
rect 18638 12356 18650 12359
rect 18874 12356 18880 12368
rect 18638 12328 18880 12356
rect 18638 12325 18650 12328
rect 18592 12319 18650 12325
rect 18874 12316 18880 12328
rect 18932 12356 18938 12368
rect 19886 12356 19892 12368
rect 18932 12328 19892 12356
rect 18932 12316 18938 12328
rect 19886 12316 19892 12328
rect 19944 12316 19950 12368
rect 19058 12288 19064 12300
rect 18371 12260 19064 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19978 12288 19984 12300
rect 19939 12260 19984 12288
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 8662 12220 8668 12232
rect 8496 12192 8668 12220
rect 6089 12183 6147 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 3234 12152 3240 12164
rect 2884 12124 3240 12152
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 7282 12152 7288 12164
rect 7024 12124 7288 12152
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 7024 12084 7052 12124
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 7374 12112 7380 12164
rect 7432 12152 7438 12164
rect 7926 12152 7932 12164
rect 7432 12124 7932 12152
rect 7432 12112 7438 12124
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 8018 12112 8024 12164
rect 8076 12152 8082 12164
rect 8772 12152 8800 12183
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10413 12223 10471 12229
rect 10413 12220 10425 12223
rect 9824 12192 10425 12220
rect 9824 12180 9830 12192
rect 10413 12189 10425 12192
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12986 12220 12992 12232
rect 12124 12192 12992 12220
rect 12124 12180 12130 12192
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12189 15623 12223
rect 15565 12183 15623 12189
rect 8076 12124 8800 12152
rect 8076 12112 8082 12124
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 10686 12152 10692 12164
rect 8904 12124 10692 12152
rect 8904 12112 8910 12124
rect 10686 12112 10692 12124
rect 10744 12112 10750 12164
rect 12250 12152 12256 12164
rect 12163 12124 12256 12152
rect 12250 12112 12256 12124
rect 12308 12152 12314 12164
rect 13096 12152 13124 12183
rect 12308 12124 13124 12152
rect 12308 12112 12314 12124
rect 1912 12056 7052 12084
rect 1912 12044 1918 12056
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7742 12084 7748 12096
rect 7156 12056 7748 12084
rect 7156 12044 7162 12056
rect 7742 12044 7748 12056
rect 7800 12084 7806 12096
rect 11790 12084 11796 12096
rect 7800 12056 11796 12084
rect 7800 12044 7806 12056
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12802 12084 12808 12096
rect 12575 12056 12808 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 15580 12084 15608 12183
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 16632 12192 17693 12220
rect 16632 12180 16638 12192
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 17862 12220 17868 12232
rect 17823 12192 17868 12220
rect 17681 12183 17739 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17954 12180 17960 12232
rect 18012 12180 18018 12232
rect 20254 12220 20260 12232
rect 20215 12192 20260 12220
rect 20254 12180 20260 12192
rect 20312 12180 20318 12232
rect 16945 12155 17003 12161
rect 16945 12121 16957 12155
rect 16991 12152 17003 12155
rect 17310 12152 17316 12164
rect 16991 12124 17316 12152
rect 16991 12121 17003 12124
rect 16945 12115 17003 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 17402 12112 17408 12164
rect 17460 12152 17466 12164
rect 17972 12152 18000 12180
rect 17460 12124 18000 12152
rect 17460 12112 17466 12124
rect 16298 12084 16304 12096
rect 15580 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 17954 12084 17960 12096
rect 17267 12056 17960 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 7469 11883 7527 11889
rect 5408 11852 6316 11880
rect 5408 11840 5414 11852
rect 4985 11815 5043 11821
rect 4985 11781 4997 11815
rect 5031 11812 5043 11815
rect 6178 11812 6184 11824
rect 5031 11784 6184 11812
rect 5031 11781 5043 11784
rect 4985 11775 5043 11781
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 6288 11812 6316 11852
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7650 11880 7656 11892
rect 7515 11852 7656 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 10594 11880 10600 11892
rect 7760 11852 10600 11880
rect 7760 11812 7788 11852
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 11793 11883 11851 11889
rect 10744 11852 11744 11880
rect 10744 11840 10750 11852
rect 11716 11824 11744 11852
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 11882 11880 11888 11892
rect 11839 11852 11888 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 14090 11880 14096 11892
rect 11992 11852 14096 11880
rect 8478 11812 8484 11824
rect 6288 11784 7788 11812
rect 7852 11784 8156 11812
rect 8439 11784 8484 11812
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3418 11744 3424 11756
rect 2547 11716 3424 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 4448 11676 4476 11707
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5316 11716 5549 11744
rect 5316 11704 5322 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 6546 11744 6552 11756
rect 5868 11716 6552 11744
rect 5868 11704 5874 11716
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 7852 11744 7880 11784
rect 8018 11744 8024 11756
rect 7668 11716 7880 11744
rect 7979 11716 8024 11744
rect 5350 11676 5356 11688
rect 2464 11648 4476 11676
rect 5311 11648 5356 11676
rect 2464 11636 2470 11648
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 7668 11676 7696 11716
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8128 11676 8156 11784
rect 8478 11772 8484 11784
rect 8536 11812 8542 11824
rect 8536 11784 8800 11812
rect 8536 11772 8542 11784
rect 8772 11753 8800 11784
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 11992 11812 12020 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 15654 11880 15660 11892
rect 14292 11852 15516 11880
rect 15615 11852 15660 11880
rect 12342 11812 12348 11824
rect 11756 11784 12020 11812
rect 12176 11784 12348 11812
rect 11756 11772 11762 11784
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 9784 11716 10548 11744
rect 8202 11676 8208 11688
rect 6227 11648 7696 11676
rect 8115 11648 8208 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 8202 11636 8208 11648
rect 8260 11676 8266 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8260 11648 8677 11676
rect 8260 11636 8266 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 9784 11676 9812 11716
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 8665 11639 8723 11645
rect 8956 11648 9812 11676
rect 9876 11648 10425 11676
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 3237 11611 3295 11617
rect 3237 11608 3249 11611
rect 3016 11580 3249 11608
rect 3016 11568 3022 11580
rect 3237 11577 3249 11580
rect 3283 11577 3295 11611
rect 3237 11571 3295 11577
rect 4154 11568 4160 11620
rect 4212 11608 4218 11620
rect 4341 11611 4399 11617
rect 4341 11608 4353 11611
rect 4212 11580 4353 11608
rect 4212 11568 4218 11580
rect 4341 11577 4353 11580
rect 4387 11577 4399 11611
rect 4341 11571 4399 11577
rect 4890 11568 4896 11620
rect 4948 11608 4954 11620
rect 5166 11608 5172 11620
rect 4948 11580 5172 11608
rect 4948 11568 4954 11580
rect 5166 11568 5172 11580
rect 5224 11568 5230 11620
rect 5442 11608 5448 11620
rect 5355 11580 5448 11608
rect 5442 11568 5448 11580
rect 5500 11608 5506 11620
rect 5500 11580 7328 11608
rect 5500 11568 5506 11580
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2866 11540 2872 11552
rect 2372 11512 2417 11540
rect 2827 11512 2872 11540
rect 2372 11500 2378 11512
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 5810 11540 5816 11552
rect 4295 11512 5816 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 5994 11540 6000 11552
rect 5955 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 7300 11540 7328 11580
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 7432 11580 7849 11608
rect 7432 11568 7438 11580
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7837 11571 7895 11577
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8956 11608 8984 11648
rect 7984 11580 8984 11608
rect 9024 11611 9082 11617
rect 7984 11568 7990 11580
rect 9024 11577 9036 11611
rect 9070 11608 9082 11611
rect 9582 11608 9588 11620
rect 9070 11580 9588 11608
rect 9070 11577 9082 11580
rect 9024 11571 9082 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 8294 11540 8300 11552
rect 7300 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9876 11540 9904 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10520 11676 10548 11716
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12176 11744 12204 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 12437 11815 12495 11821
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 12483 11784 13492 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 12986 11744 12992 11756
rect 11940 11716 12204 11744
rect 12360 11716 12664 11744
rect 12947 11716 12992 11744
rect 11940 11704 11946 11716
rect 12158 11676 12164 11688
rect 10520 11648 12164 11676
rect 10413 11639 10471 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12360 11676 12388 11716
rect 12299 11648 12388 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 10658 11611 10716 11617
rect 10658 11608 10670 11611
rect 10244 11580 10670 11608
rect 10244 11552 10272 11580
rect 10658 11577 10670 11580
rect 10704 11577 10716 11611
rect 12636 11608 12664 11716
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13464 11685 13492 11784
rect 14292 11753 14320 11852
rect 15488 11812 15516 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 18049 11883 18107 11889
rect 15896 11852 17264 11880
rect 15896 11840 15902 11852
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 15488 11784 16037 11812
rect 16025 11781 16037 11784
rect 16071 11781 16083 11815
rect 17236 11812 17264 11852
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 19978 11880 19984 11892
rect 18095 11852 19984 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 20990 11880 20996 11892
rect 20947 11852 20996 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 18690 11812 18696 11824
rect 17236 11784 18696 11812
rect 16025 11775 16083 11781
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 16040 11744 16068 11775
rect 18690 11772 18696 11784
rect 18748 11772 18754 11824
rect 16298 11744 16304 11756
rect 16040 11716 16304 11744
rect 14277 11707 14335 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17368 11716 18613 11744
rect 17368 11704 17374 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 15286 11676 15292 11688
rect 13449 11639 13507 11645
rect 13617 11648 15292 11676
rect 13617 11608 13645 11648
rect 15286 11636 15292 11648
rect 15344 11676 15350 11688
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 15344 11648 16221 11676
rect 15344 11636 15350 11648
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16568 11679 16626 11685
rect 16568 11645 16580 11679
rect 16614 11676 16626 11679
rect 17328 11676 17356 11704
rect 16614 11648 17356 11676
rect 16614 11645 16626 11648
rect 16568 11639 16626 11645
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 18012 11648 18429 11676
rect 18012 11636 18018 11648
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 19058 11676 19064 11688
rect 19019 11648 19064 11676
rect 18417 11639 18475 11645
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 19334 11685 19340 11688
rect 19328 11676 19340 11685
rect 19295 11648 19340 11676
rect 19328 11639 19340 11648
rect 19334 11636 19340 11639
rect 19392 11636 19398 11688
rect 20714 11676 20720 11688
rect 20675 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 13722 11608 13728 11620
rect 12636 11580 13645 11608
rect 13683 11580 13728 11608
rect 10658 11571 10716 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 14550 11617 14556 11620
rect 14544 11608 14556 11617
rect 14511 11580 14556 11608
rect 14544 11571 14556 11580
rect 14550 11568 14556 11571
rect 14608 11568 14614 11620
rect 17696 11580 19380 11608
rect 8536 11512 9904 11540
rect 10137 11543 10195 11549
rect 8536 11500 8542 11512
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10226 11540 10232 11552
rect 10183 11512 10232 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 11020 11512 12081 11540
rect 11020 11500 11026 11512
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 12069 11503 12127 11509
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12400 11512 12909 11540
rect 12400 11500 12406 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 17586 11540 17592 11552
rect 13136 11512 17592 11540
rect 13136 11500 13142 11512
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 17696 11549 17724 11580
rect 19352 11552 19380 11580
rect 17681 11543 17739 11549
rect 17681 11509 17693 11543
rect 17727 11509 17739 11543
rect 18506 11540 18512 11552
rect 18467 11512 18512 11540
rect 17681 11503 17739 11509
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19334 11500 19340 11552
rect 19392 11500 19398 11552
rect 20438 11540 20444 11552
rect 20399 11512 20444 11540
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 2832 11308 3525 11336
rect 2832 11296 2838 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 3513 11299 3571 11305
rect 4356 11308 5917 11336
rect 1872 11240 4108 11268
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 1872 11209 1900 11240
rect 4080 11212 4108 11240
rect 1857 11203 1915 11209
rect 1857 11200 1869 11203
rect 1820 11172 1869 11200
rect 1820 11160 1826 11172
rect 1857 11169 1869 11172
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 2124 11203 2182 11209
rect 2124 11169 2136 11203
rect 2170 11200 2182 11203
rect 2406 11200 2412 11212
rect 2170 11172 2412 11200
rect 2170 11169 2182 11172
rect 2124 11163 2182 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 4356 11209 4384 11308
rect 5905 11305 5917 11308
rect 5951 11336 5963 11339
rect 5994 11336 6000 11348
rect 5951 11308 6000 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 6880 11308 7389 11336
rect 6880 11296 6886 11308
rect 7377 11305 7389 11308
rect 7423 11336 7435 11339
rect 7561 11339 7619 11345
rect 7561 11336 7573 11339
rect 7423 11308 7573 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7561 11305 7573 11308
rect 7607 11305 7619 11339
rect 7561 11299 7619 11305
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7800 11308 8125 11336
rect 7800 11296 7806 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 12897 11339 12955 11345
rect 8113 11299 8171 11305
rect 8220 11308 12848 11336
rect 8220 11268 8248 11308
rect 4448 11240 8248 11268
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 4120 11172 4353 11200
rect 4120 11160 4126 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 4448 11132 4476 11240
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 10778 11268 10784 11280
rect 8352 11240 10784 11268
rect 8352 11228 8358 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 11784 11271 11842 11277
rect 11784 11237 11796 11271
rect 11830 11268 11842 11271
rect 12250 11268 12256 11280
rect 11830 11240 12256 11268
rect 11830 11237 11842 11240
rect 11784 11231 11842 11237
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12434 11228 12440 11280
rect 12492 11228 12498 11280
rect 12820 11268 12848 11308
rect 12897 11305 12909 11339
rect 12943 11336 12955 11339
rect 12986 11336 12992 11348
rect 12943 11308 12992 11336
rect 12943 11305 12955 11308
rect 12897 11299 12955 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13096 11308 14044 11336
rect 13096 11268 13124 11308
rect 12820 11240 13124 11268
rect 13538 11228 13544 11280
rect 13596 11277 13602 11280
rect 13596 11271 13660 11277
rect 13596 11237 13614 11271
rect 13648 11237 13660 11271
rect 14016 11268 14044 11308
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 14148 11308 15761 11336
rect 14148 11296 14154 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 16347 11308 17785 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 17773 11305 17785 11308
rect 17819 11305 17831 11339
rect 17773 11299 17831 11305
rect 18417 11339 18475 11345
rect 18417 11305 18429 11339
rect 18463 11336 18475 11339
rect 18782 11336 18788 11348
rect 18463 11308 18788 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 20346 11336 20352 11348
rect 18923 11308 20352 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 15470 11268 15476 11280
rect 14016 11240 15476 11268
rect 13596 11231 13660 11237
rect 13596 11228 13602 11231
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 15657 11271 15715 11277
rect 15657 11237 15669 11271
rect 15703 11268 15715 11271
rect 15838 11268 15844 11280
rect 15703 11240 15844 11268
rect 15703 11237 15715 11240
rect 15657 11231 15715 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 16850 11268 16856 11280
rect 16040 11240 16856 11268
rect 4608 11203 4666 11209
rect 4608 11169 4620 11203
rect 4654 11200 4666 11203
rect 5442 11200 5448 11212
rect 4654 11172 5448 11200
rect 4654 11169 4666 11172
rect 4608 11163 4666 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6253 11203 6311 11209
rect 6253 11200 6265 11203
rect 5736 11172 6265 11200
rect 3660 11104 4476 11132
rect 3660 11092 3666 11104
rect 3237 11067 3295 11073
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3510 11064 3516 11076
rect 3283 11036 3516 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5736 11073 5764 11172
rect 6253 11169 6265 11172
rect 6299 11169 6311 11203
rect 6253 11163 6311 11169
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7524 11172 8033 11200
rect 7524 11160 7530 11172
rect 8021 11169 8033 11172
rect 8067 11200 8079 11203
rect 8067 11172 9352 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5951 11104 6009 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 7607 11104 8217 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5592 11036 5733 11064
rect 5592 11024 5598 11036
rect 5721 11033 5733 11036
rect 5767 11033 5779 11067
rect 7650 11064 7656 11076
rect 7611 11036 7656 11064
rect 5721 11027 5779 11033
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 9324 11064 9352 11172
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9824 11172 10057 11200
rect 9824 11160 9830 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11020 11172 11529 11200
rect 11020 11160 11026 11172
rect 11517 11169 11529 11172
rect 11563 11200 11575 11203
rect 12452 11200 12480 11228
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 11563 11172 13369 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 15562 11200 15568 11212
rect 13357 11163 13415 11169
rect 13464 11172 15568 11200
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 13464 11132 13492 11172
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 10284 11104 10329 11132
rect 13372 11104 13492 11132
rect 10284 11092 10290 11104
rect 13372 11064 13400 11104
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 14608 11104 15945 11132
rect 14608 11092 14614 11104
rect 14752 11073 14780 11104
rect 15933 11101 15945 11104
rect 15979 11132 15991 11135
rect 16040 11132 16068 11240
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 16942 11200 16948 11212
rect 16715 11172 16948 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17678 11200 17684 11212
rect 17639 11172 17684 11200
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 18785 11203 18843 11209
rect 18785 11200 18797 11203
rect 17828 11172 18797 11200
rect 17828 11160 17834 11172
rect 18785 11169 18797 11172
rect 18831 11169 18843 11203
rect 20162 11200 20168 11212
rect 20123 11172 20168 11200
rect 18785 11163 18843 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 16758 11132 16764 11144
rect 15979 11104 16068 11132
rect 16719 11104 16764 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17862 11132 17868 11144
rect 16908 11104 16953 11132
rect 17823 11104 17868 11132
rect 16908 11092 16914 11104
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 18969 11135 19027 11141
rect 18969 11132 18981 11135
rect 18932 11104 18981 11132
rect 18932 11092 18938 11104
rect 18969 11101 18981 11104
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 19058 11092 19064 11144
rect 19116 11132 19122 11144
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19116 11104 20269 11132
rect 19116 11092 19122 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20404 11104 20449 11132
rect 20404 11092 20410 11104
rect 9324 11036 11560 11064
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 4154 10996 4160 11008
rect 3200 10968 4160 10996
rect 3200 10956 3206 10968
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 7834 10996 7840 11008
rect 5040 10968 7840 10996
rect 5040 10956 5046 10968
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 9674 10996 9680 11008
rect 9635 10968 9680 10996
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 11532 10996 11560 11036
rect 12452 11036 13400 11064
rect 14737 11067 14795 11073
rect 12452 10996 12480 11036
rect 14737 11033 14749 11067
rect 14783 11033 14795 11067
rect 14737 11027 14795 11033
rect 15289 11067 15347 11073
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 16574 11064 16580 11076
rect 15335 11036 16580 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 18506 11064 18512 11076
rect 17359 11036 18512 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 11532 10968 12480 10996
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 17034 10996 17040 11008
rect 12952 10968 17040 10996
rect 12952 10956 12958 10968
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 19797 10999 19855 11005
rect 19797 10965 19809 10999
rect 19843 10996 19855 10999
rect 20070 10996 20076 11008
rect 19843 10968 20076 10996
rect 19843 10965 19855 10968
rect 19797 10959 19855 10965
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1728 10764 2053 10792
rect 1728 10752 1734 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3142 10792 3148 10804
rect 3099 10764 3148 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 8478 10792 8484 10804
rect 6840 10764 8484 10792
rect 5460 10724 5488 10752
rect 5460 10696 6316 10724
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3510 10656 3516 10668
rect 2731 10628 3516 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3660 10628 3705 10656
rect 3660 10616 3666 10628
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 6178 10656 6184 10668
rect 4028 10628 4200 10656
rect 6139 10628 6184 10656
rect 4028 10616 4034 10628
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3878 10588 3884 10600
rect 2547 10560 3884 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4172 10588 4200 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6288 10665 6316 10696
rect 6840 10665 6868 10764
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9766 10792 9772 10804
rect 9079 10764 9772 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 12158 10792 12164 10804
rect 10244 10764 12164 10792
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 10244 10724 10272 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 18693 10795 18751 10801
rect 12299 10764 17172 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 7892 10696 10272 10724
rect 11333 10727 11391 10733
rect 7892 10684 7898 10696
rect 11333 10693 11345 10727
rect 11379 10724 11391 10727
rect 12342 10724 12348 10736
rect 11379 10696 12348 10724
rect 11379 10693 11391 10696
rect 11333 10687 11391 10693
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 15286 10724 15292 10736
rect 13872 10696 14964 10724
rect 15247 10696 15292 10724
rect 13872 10684 13878 10696
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 6825 10619 6883 10625
rect 9582 10616 9588 10628
rect 9640 10656 9646 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9640 10628 10609 10656
rect 9640 10616 9646 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11664 10628 11805 10656
rect 11664 10616 11670 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12250 10656 12256 10668
rect 12023 10628 12256 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 14366 10656 14372 10668
rect 13596 10628 14372 10656
rect 13596 10616 13602 10628
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14424 10628 14841 10656
rect 14424 10616 14430 10628
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 14936 10656 14964 10696
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 16390 10724 16396 10736
rect 16351 10696 16396 10724
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 15010 10656 15016 10668
rect 14923 10628 15016 10656
rect 14829 10619 14887 10625
rect 15010 10616 15016 10628
rect 15068 10656 15074 10668
rect 15933 10659 15991 10665
rect 15068 10628 15516 10656
rect 15068 10616 15074 10628
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 4172 10560 6224 10588
rect 3421 10523 3479 10529
rect 3421 10489 3433 10523
rect 3467 10520 3479 10523
rect 4154 10520 4160 10532
rect 3467 10492 4160 10520
rect 3467 10489 3479 10492
rect 3421 10483 3479 10489
rect 4154 10480 4160 10492
rect 4212 10480 4218 10532
rect 4332 10523 4390 10529
rect 4332 10489 4344 10523
rect 4378 10520 4390 10523
rect 5166 10520 5172 10532
rect 4378 10492 5172 10520
rect 4378 10489 4390 10492
rect 4332 10483 4390 10489
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 6089 10523 6147 10529
rect 6089 10520 6101 10523
rect 5316 10492 6101 10520
rect 5316 10480 5322 10492
rect 6089 10489 6101 10492
rect 6135 10489 6147 10523
rect 6196 10520 6224 10560
rect 6932 10560 9505 10588
rect 6932 10520 6960 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12704 10591 12762 10597
rect 12492 10560 12537 10588
rect 12492 10548 12498 10560
rect 12704 10557 12716 10591
rect 12750 10588 12762 10591
rect 12986 10588 12992 10600
rect 12750 10560 12992 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 15488 10597 15516 10628
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16206 10656 16212 10668
rect 15979 10628 16212 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16724 10628 16957 10656
rect 16724 10616 16730 10628
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10557 15531 10591
rect 17144 10588 17172 10764
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 19058 10792 19064 10804
rect 18739 10764 19064 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19150 10656 19156 10668
rect 19111 10628 19156 10656
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19337 10659 19395 10665
rect 19337 10625 19349 10659
rect 19383 10656 19395 10659
rect 19383 10628 19840 10656
rect 19383 10625 19395 10628
rect 19337 10619 19395 10625
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 17144 10560 19073 10588
rect 15473 10551 15531 10557
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 19484 10560 19717 10588
rect 19484 10548 19490 10560
rect 19705 10557 19717 10560
rect 19751 10557 19763 10591
rect 19812 10588 19840 10628
rect 19972 10591 20030 10597
rect 19972 10588 19984 10591
rect 19812 10560 19984 10588
rect 19705 10551 19763 10557
rect 19972 10557 19984 10560
rect 20018 10588 20030 10591
rect 20438 10588 20444 10600
rect 20018 10560 20444 10588
rect 20018 10557 20030 10560
rect 19972 10551 20030 10557
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 6196 10492 6960 10520
rect 7092 10523 7150 10529
rect 6089 10483 6147 10489
rect 7092 10489 7104 10523
rect 7138 10520 7150 10523
rect 7742 10520 7748 10532
rect 7138 10492 7748 10520
rect 7138 10489 7150 10492
rect 7092 10483 7150 10489
rect 7742 10480 7748 10492
rect 7800 10480 7806 10532
rect 8573 10523 8631 10529
rect 8573 10489 8585 10523
rect 8619 10520 8631 10523
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 8619 10492 9413 10520
rect 8619 10489 8631 10492
rect 8573 10483 8631 10489
rect 9401 10489 9413 10492
rect 9447 10489 9459 10523
rect 9401 10483 9459 10489
rect 10413 10523 10471 10529
rect 10413 10489 10425 10523
rect 10459 10520 10471 10523
rect 10962 10520 10968 10532
rect 10459 10492 10968 10520
rect 10459 10489 10471 10492
rect 10413 10483 10471 10489
rect 10962 10480 10968 10492
rect 11020 10520 11026 10532
rect 11020 10492 12572 10520
rect 11020 10480 11026 10492
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 5718 10452 5724 10464
rect 3568 10424 3613 10452
rect 5679 10424 5724 10452
rect 3568 10412 3574 10424
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 6972 10424 8217 10452
rect 6972 10412 6978 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 10318 10452 10324 10464
rect 9364 10424 10324 10452
rect 9364 10412 9370 10424
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11698 10452 11704 10464
rect 10560 10424 10605 10452
rect 11659 10424 11704 10452
rect 10560 10412 10566 10424
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 11848 10424 12265 10452
rect 11848 10412 11854 10424
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12544 10452 12572 10492
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 14645 10523 14703 10529
rect 14645 10520 14657 10523
rect 12676 10492 14657 10520
rect 12676 10480 12682 10492
rect 14645 10489 14657 10492
rect 14691 10489 14703 10523
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 14645 10483 14703 10489
rect 15212 10492 16773 10520
rect 12894 10452 12900 10464
rect 12544 10424 12900 10452
rect 12253 10415 12311 10421
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13044 10424 13829 10452
rect 13044 10412 13050 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 14458 10452 14464 10464
rect 14323 10424 14464 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14737 10455 14795 10461
rect 14737 10421 14749 10455
rect 14783 10452 14795 10455
rect 15212 10452 15240 10492
rect 16761 10489 16773 10492
rect 16807 10520 16819 10523
rect 17126 10520 17132 10532
rect 16807 10492 17132 10520
rect 16807 10489 16819 10492
rect 16761 10483 16819 10489
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 14783 10424 15240 10452
rect 14783 10421 14795 10424
rect 14737 10415 14795 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 16022 10452 16028 10464
rect 15344 10424 16028 10452
rect 15344 10412 15350 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 17954 10452 17960 10464
rect 16899 10424 17960 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 21085 10455 21143 10461
rect 21085 10452 21097 10455
rect 20404 10424 21097 10452
rect 20404 10412 20410 10424
rect 21085 10421 21097 10424
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2096 10220 2268 10248
rect 2096 10208 2102 10220
rect 2240 10180 2268 10220
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 2556 10220 3157 10248
rect 2556 10208 2562 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 3145 10211 3203 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4663 10220 5273 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5408 10220 5856 10248
rect 5408 10208 5414 10220
rect 2590 10180 2596 10192
rect 2240 10152 2596 10180
rect 2590 10140 2596 10152
rect 2648 10180 2654 10192
rect 3602 10180 3608 10192
rect 2648 10152 3608 10180
rect 2648 10140 2654 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 4709 10183 4767 10189
rect 4709 10149 4721 10183
rect 4755 10180 4767 10183
rect 5718 10180 5724 10192
rect 4755 10152 5724 10180
rect 4755 10149 4767 10152
rect 4709 10143 4767 10149
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 1762 10112 1768 10124
rect 1723 10084 1768 10112
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 2038 10121 2044 10124
rect 2032 10112 2044 10121
rect 1999 10084 2044 10112
rect 2032 10075 2044 10084
rect 2038 10072 2044 10075
rect 2096 10072 2102 10124
rect 5626 10112 5632 10124
rect 5587 10084 5632 10112
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5828 10112 5856 10220
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7466 10248 7472 10260
rect 7064 10220 7472 10248
rect 7064 10208 7070 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8113 10251 8171 10257
rect 8113 10217 8125 10251
rect 8159 10248 8171 10251
rect 8202 10248 8208 10260
rect 8159 10220 8208 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 9640 10220 11069 10248
rect 9640 10208 9646 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10217 11667 10251
rect 11974 10248 11980 10260
rect 11935 10220 11980 10248
rect 11609 10211 11667 10217
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7374 10180 7380 10192
rect 7156 10152 7380 10180
rect 7156 10140 7162 10152
rect 7374 10140 7380 10152
rect 7432 10140 7438 10192
rect 9674 10180 9680 10192
rect 8864 10152 9680 10180
rect 5736 10084 5856 10112
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5534 10044 5540 10056
rect 4939 10016 5540 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5736 10053 5764 10084
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6178 10112 6184 10124
rect 6052 10084 6184 10112
rect 6052 10072 6058 10084
rect 6178 10072 6184 10084
rect 6236 10112 6242 10124
rect 6457 10115 6515 10121
rect 6457 10112 6469 10115
rect 6236 10084 6469 10112
rect 6236 10072 6242 10084
rect 6457 10081 6469 10084
rect 6503 10081 6515 10115
rect 6457 10075 6515 10081
rect 6724 10115 6782 10121
rect 6724 10081 6736 10115
rect 6770 10112 6782 10115
rect 7558 10112 7564 10124
rect 6770 10084 7564 10112
rect 6770 10081 6782 10084
rect 6724 10075 6782 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8864 10121 8892 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 8260 10084 8309 10112
rect 8260 10072 8266 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8849 10115 8907 10121
rect 8849 10081 8861 10115
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 9944 10115 10002 10121
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10226 10112 10232 10124
rect 9990 10084 10232 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11624 10112 11652 10211
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13814 10248 13820 10260
rect 13679 10220 13820 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10217 14059 10251
rect 14458 10248 14464 10260
rect 14419 10220 14464 10248
rect 14001 10211 14059 10217
rect 14016 10180 14044 10211
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15930 10248 15936 10260
rect 15335 10220 15936 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 16724 10220 18337 10248
rect 16724 10208 16730 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20220 10220 20913 10248
rect 20220 10208 20226 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 17678 10180 17684 10192
rect 14016 10152 17684 10180
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 18417 10183 18475 10189
rect 18417 10149 18429 10183
rect 18463 10180 18475 10183
rect 19426 10180 19432 10192
rect 18463 10152 19432 10180
rect 18463 10149 18475 10152
rect 18417 10143 18475 10149
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 11624 10084 13001 10112
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 12989 10075 13047 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 13964 10084 14381 10112
rect 13964 10072 13970 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 14369 10075 14427 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 18616 10121 18644 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 17212 10115 17270 10121
rect 17212 10081 17224 10115
rect 17258 10112 17270 10115
rect 18601 10115 18659 10121
rect 17258 10084 18552 10112
rect 17258 10081 17270 10084
rect 17212 10075 17270 10081
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 5813 10007 5871 10013
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 5828 9976 5856 10007
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 5500 9948 5856 9976
rect 5500 9936 5506 9948
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9692 9976 9720 10007
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11790 10044 11796 10056
rect 11112 10016 11796 10044
rect 11112 10004 11118 10016
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12250 10044 12256 10056
rect 12211 10016 12256 10044
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12492 10016 13093 10044
rect 12492 10004 12498 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 14550 10044 14556 10056
rect 13228 10016 13273 10044
rect 14511 10016 14556 10044
rect 13228 10004 13234 10016
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 8536 9948 9720 9976
rect 8536 9936 8542 9948
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 10870 9908 10876 9920
rect 4120 9880 10876 9908
rect 4120 9868 4126 9880
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 16114 9908 16120 9920
rect 11848 9880 16120 9908
rect 11848 9868 11854 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16960 9908 16988 10007
rect 18417 9911 18475 9917
rect 18417 9908 18429 9911
rect 16960 9880 18429 9908
rect 18417 9877 18429 9880
rect 18463 9877 18475 9911
rect 18524 9908 18552 10084
rect 18601 10081 18613 10115
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18868 10115 18926 10121
rect 18868 10081 18880 10115
rect 18914 10112 18926 10115
rect 19794 10112 19800 10124
rect 18914 10084 19800 10112
rect 18914 10081 18926 10084
rect 18868 10075 18926 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 20254 10112 20260 10124
rect 20215 10084 20260 10112
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9976 20499 9979
rect 20622 9976 20628 9988
rect 20487 9948 20628 9976
rect 20487 9945 20499 9948
rect 20441 9939 20499 9945
rect 20622 9936 20628 9948
rect 20680 9936 20686 9988
rect 18782 9908 18788 9920
rect 18524 9880 18788 9908
rect 18417 9871 18475 9877
rect 18782 9868 18788 9880
rect 18840 9908 18846 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 18840 9880 19993 9908
rect 18840 9868 18846 9880
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2406 9704 2412 9716
rect 1903 9676 2412 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 10042 9704 10048 9716
rect 4028 9676 10048 9704
rect 4028 9664 4034 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10502 9704 10508 9716
rect 10463 9676 10508 9704
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 10836 9676 11008 9704
rect 10836 9664 10842 9676
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3326 9636 3332 9648
rect 2915 9608 3332 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 4798 9636 4804 9648
rect 4759 9608 4804 9636
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6788 9608 6837 9636
rect 6788 9596 6794 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 7616 9608 7880 9636
rect 7616 9596 7622 9608
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1912 9540 2329 9568
rect 1912 9528 1918 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2317 9531 2375 9537
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2740 9540 3433 9568
rect 2740 9528 2746 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5132 9540 5273 9568
rect 5132 9528 5138 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 6914 9568 6920 9580
rect 5491 9540 6920 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7742 9568 7748 9580
rect 7515 9540 7748 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 7852 9568 7880 9608
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 7852 9540 8401 9568
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8536 9540 8861 9568
rect 8536 9528 8542 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 10244 9568 10272 9664
rect 10980 9636 11008 9676
rect 12452 9676 13400 9704
rect 10980 9608 11192 9636
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10244 9540 11069 9568
rect 8849 9531 8907 9537
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2866 9500 2872 9512
rect 2271 9472 2872 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 7190 9500 7196 9512
rect 3660 9472 7196 9500
rect 3660 9460 3666 9472
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 7708 9472 8309 9500
rect 7708 9460 7714 9472
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 10686 9500 10692 9512
rect 8297 9463 8355 9469
rect 8404 9472 10692 9500
rect 1397 9435 1455 9441
rect 1397 9401 1409 9435
rect 1443 9432 1455 9435
rect 1443 9404 2452 9432
rect 1443 9401 1455 9404
rect 1397 9395 1455 9401
rect 2424 9364 2452 9404
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 8404 9432 8432 9472
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11164 9500 11192 9608
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 12452 9636 12480 9676
rect 11388 9608 12480 9636
rect 13372 9636 13400 9676
rect 14108 9676 16712 9704
rect 14108 9636 14136 9676
rect 13372 9608 14136 9636
rect 14185 9639 14243 9645
rect 11388 9596 11394 9608
rect 14185 9605 14197 9639
rect 14231 9636 14243 9639
rect 15654 9636 15660 9648
rect 14231 9608 15660 9636
rect 14231 9605 14243 9608
rect 14185 9599 14243 9605
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 16684 9636 16712 9676
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 16945 9707 17003 9713
rect 16945 9704 16957 9707
rect 16816 9676 16957 9704
rect 16816 9664 16822 9676
rect 16945 9673 16957 9676
rect 16991 9673 17003 9707
rect 16945 9667 17003 9673
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18049 9707 18107 9713
rect 18049 9704 18061 9707
rect 18012 9676 18061 9704
rect 18012 9664 18018 9676
rect 18049 9673 18061 9676
rect 18095 9673 18107 9707
rect 18049 9667 18107 9673
rect 17770 9636 17776 9648
rect 16684 9608 17776 9636
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 14608 9540 14749 9568
rect 14608 9528 14614 9540
rect 14737 9537 14749 9540
rect 14783 9537 14795 9571
rect 15841 9571 15899 9577
rect 15841 9568 15853 9571
rect 14737 9531 14795 9537
rect 15396 9540 15853 9568
rect 11238 9500 11244 9512
rect 11011 9472 11244 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12526 9500 12532 9512
rect 12483 9472 12532 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 15396 9500 15424 9540
rect 15841 9537 15853 9540
rect 15887 9568 15899 9571
rect 16390 9568 16396 9580
rect 15887 9540 16396 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 17494 9568 17500 9580
rect 17455 9540 17500 9568
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18782 9568 18788 9580
rect 18739 9540 18788 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 19484 9540 19717 9568
rect 19484 9528 19490 9540
rect 19705 9537 19717 9540
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 14016 9472 15424 9500
rect 14016 9444 14044 9472
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 15528 9472 15669 9500
rect 15528 9460 15534 9472
rect 15657 9469 15669 9472
rect 15703 9469 15715 9503
rect 15657 9463 15715 9469
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18598 9500 18604 9512
rect 17828 9472 18604 9500
rect 17828 9460 17834 9472
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19972 9503 20030 9509
rect 19972 9469 19984 9503
rect 20018 9500 20030 9503
rect 20346 9500 20352 9512
rect 20018 9472 20352 9500
rect 20018 9469 20030 9472
rect 19972 9463 20030 9469
rect 20346 9460 20352 9472
rect 20404 9460 20410 9512
rect 4120 9404 8432 9432
rect 9116 9435 9174 9441
rect 4120 9392 4126 9404
rect 9116 9401 9128 9435
rect 9162 9432 9174 9435
rect 9858 9432 9864 9444
rect 9162 9404 9864 9432
rect 9162 9401 9174 9404
rect 9116 9395 9174 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 12704 9435 12762 9441
rect 10928 9404 10973 9432
rect 10928 9392 10934 9404
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 13078 9432 13084 9444
rect 12750 9404 13084 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 13998 9432 14004 9444
rect 13832 9404 14004 9432
rect 2958 9364 2964 9376
rect 2424 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3108 9336 3341 9364
rect 3108 9324 3114 9336
rect 3329 9333 3341 9336
rect 3375 9364 3387 9367
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 3375 9336 5181 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6972 9336 7205 9364
rect 6972 9324 6978 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7331 9336 7849 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9364 8263 9367
rect 8294 9364 8300 9376
rect 8251 9336 8300 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 13832 9373 13860 9404
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 14553 9435 14611 9441
rect 14553 9401 14565 9435
rect 14599 9432 14611 9435
rect 15565 9435 15623 9441
rect 14599 9404 15240 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 8536 9336 13829 9364
rect 8536 9324 8542 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 15212 9373 15240 9404
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 15611 9404 16221 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 17402 9432 17408 9444
rect 17315 9404 17408 9432
rect 16209 9395 16267 9401
rect 17402 9392 17408 9404
rect 17460 9432 17466 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 17460 9404 18521 9432
rect 17460 9392 17466 9404
rect 18509 9401 18521 9404
rect 18555 9432 18567 9435
rect 20438 9432 20444 9444
rect 18555 9404 20444 9432
rect 18555 9401 18567 9404
rect 18509 9395 18567 9401
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13964 9336 14657 9364
rect 13964 9324 13970 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14645 9327 14703 9333
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9333 15255 9367
rect 15197 9327 15255 9333
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 16356 9336 17325 9364
rect 16356 9324 16362 9336
rect 17313 9333 17325 9336
rect 17359 9333 17371 9367
rect 18414 9364 18420 9376
rect 18375 9336 18420 9364
rect 17313 9327 17371 9333
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 21085 9367 21143 9373
rect 21085 9364 21097 9367
rect 18656 9336 21097 9364
rect 18656 9324 18662 9336
rect 21085 9333 21097 9336
rect 21131 9333 21143 9367
rect 21085 9327 21143 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2314 9160 2320 9172
rect 2087 9132 2320 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5626 9160 5632 9172
rect 4571 9132 5632 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 7558 9160 7564 9172
rect 7519 9132 7564 9160
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 7668 9132 10824 9160
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 7668 9092 7696 9132
rect 4120 9064 7696 9092
rect 7745 9095 7803 9101
rect 4120 9052 4126 9064
rect 7745 9061 7757 9095
rect 7791 9092 7803 9095
rect 9766 9092 9772 9104
rect 7791 9064 9772 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 9968 9064 10057 9092
rect 9968 9036 9996 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 10134 9052 10140 9104
rect 10192 9092 10198 9104
rect 10796 9092 10824 9132
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11330 9160 11336 9172
rect 10928 9132 11336 9160
rect 10928 9120 10934 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12584 9132 12664 9160
rect 12584 9120 12590 9132
rect 12342 9092 12348 9104
rect 10192 9064 10237 9092
rect 10796 9064 12348 9092
rect 10192 9052 10198 9064
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 3142 9024 3148 9036
rect 2455 8996 3148 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 4939 8996 5549 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 6178 9024 6184 9036
rect 6139 8996 6184 9024
rect 5537 8987 5595 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6448 9027 6506 9033
rect 6448 8993 6460 9027
rect 6494 9024 6506 9027
rect 6730 9024 6736 9036
rect 6494 8996 6736 9024
rect 6494 8993 6506 8996
rect 6448 8987 6506 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7650 9024 7656 9036
rect 7248 8996 7656 9024
rect 7248 8984 7254 8996
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8386 9024 8392 9036
rect 8343 8996 8392 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 2501 8919 2559 8925
rect 2516 8888 2544 8919
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 2924 8928 4997 8956
rect 2924 8916 2930 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 5166 8956 5172 8968
rect 5127 8928 5172 8956
rect 4985 8919 5043 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 8220 8956 8248 8987
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 9088 8996 9137 9024
rect 9088 8984 9094 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9950 8984 9956 9036
rect 10008 8984 10014 9036
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10778 9024 10784 9036
rect 10735 8996 10784 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 8478 8956 8484 8968
rect 7208 8928 8248 8956
rect 8439 8928 8484 8956
rect 5074 8888 5080 8900
rect 2516 8860 5080 8888
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 7208 8820 7236 8928
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8720 8928 9229 8956
rect 8720 8916 8726 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9398 8956 9404 8968
rect 9359 8928 9404 8956
rect 9217 8919 9275 8925
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 12536 8959 12594 8965
rect 12536 8925 12548 8959
rect 12582 8956 12594 8959
rect 12636 8956 12664 9132
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13136 9132 13921 9160
rect 13136 9120 13142 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 15746 9160 15752 9172
rect 14231 9132 15752 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 15988 9132 16681 9160
rect 15988 9120 15994 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 16669 9123 16727 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 17405 9163 17463 9169
rect 17405 9129 17417 9163
rect 17451 9160 17463 9163
rect 18414 9160 18420 9172
rect 17451 9132 18420 9160
rect 17451 9129 17463 9132
rect 17405 9123 17463 9129
rect 12710 9052 12716 9104
rect 12768 9101 12774 9104
rect 12768 9095 12832 9101
rect 12768 9061 12786 9095
rect 12820 9061 12832 9095
rect 12768 9055 12832 9061
rect 12768 9052 12774 9055
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 14553 9095 14611 9101
rect 14553 9092 14565 9095
rect 12952 9064 14565 9092
rect 12952 9052 12958 9064
rect 14553 9061 14565 9064
rect 14599 9061 14611 9095
rect 15286 9092 15292 9104
rect 14553 9055 14611 9061
rect 14660 9064 15292 9092
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 14660 9024 14688 9064
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 16298 9052 16304 9104
rect 16356 9092 16362 9104
rect 17420 9092 17448 9123
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 19794 9160 19800 9172
rect 19755 9132 19800 9160
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 16356 9064 17448 9092
rect 16356 9052 16362 9064
rect 15545 9027 15603 9033
rect 15545 9024 15557 9027
rect 13136 8996 14688 9024
rect 14752 8996 15557 9024
rect 13136 8984 13142 8996
rect 14642 8956 14648 8968
rect 12582 8928 12664 8956
rect 14603 8928 14648 8956
rect 12582 8925 12594 8928
rect 12536 8919 12594 8925
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7791 8860 7849 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8168 8860 9628 8888
rect 8168 8848 8174 8860
rect 6420 8792 7236 8820
rect 6420 8780 6426 8792
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 8294 8820 8300 8832
rect 7340 8792 8300 8820
rect 7340 8780 7346 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9490 8820 9496 8832
rect 8803 8792 9496 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9600 8820 9628 8860
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 9732 8860 9777 8888
rect 9732 8848 9738 8860
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10244 8888 10272 8919
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 14752 8965 14780 8996
rect 15545 8993 15557 8996
rect 15591 8993 15603 9027
rect 15545 8987 15603 8993
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 17678 9024 17684 9036
rect 17359 8996 17684 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18684 9027 18742 9033
rect 18684 8993 18696 9027
rect 18730 9024 18742 9027
rect 19426 9024 19432 9036
rect 18730 8996 19432 9024
rect 18730 8993 18742 8996
rect 18684 8987 18742 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 19886 8984 19892 9036
rect 19944 9024 19950 9036
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 19944 8996 20269 9024
rect 19944 8984 19950 8996
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8925 14795 8959
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 14737 8919 14795 8925
rect 9916 8860 10272 8888
rect 9916 8848 9922 8860
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 14752 8888 14780 8919
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 17552 8928 17645 8956
rect 17552 8916 17558 8928
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 18012 8928 18429 8956
rect 18012 8916 18018 8928
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 14826 8888 14832 8900
rect 14608 8860 14832 8888
rect 14608 8848 14614 8860
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 11977 8823 12035 8829
rect 11977 8820 11989 8823
rect 9600 8792 11989 8820
rect 11977 8789 11989 8792
rect 12023 8820 12035 8823
rect 13814 8820 13820 8832
rect 12023 8792 13820 8820
rect 12023 8789 12035 8792
rect 11977 8783 12035 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 17512 8820 17540 8916
rect 19610 8848 19616 8900
rect 19668 8888 19674 8900
rect 20441 8891 20499 8897
rect 20441 8888 20453 8891
rect 19668 8860 20453 8888
rect 19668 8848 19674 8860
rect 20441 8857 20453 8860
rect 20487 8857 20499 8891
rect 20441 8851 20499 8857
rect 14424 8792 17540 8820
rect 14424 8780 14430 8792
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 2648 8588 3249 8616
rect 2648 8576 2654 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3568 8588 4077 8616
rect 3568 8576 3574 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 7834 8616 7840 8628
rect 4948 8588 7840 8616
rect 4948 8576 4954 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8202 8616 8208 8628
rect 7975 8588 8208 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 12069 8619 12127 8625
rect 10744 8588 12020 8616
rect 10744 8576 10750 8588
rect 4430 8508 4436 8560
rect 4488 8548 4494 8560
rect 4982 8548 4988 8560
rect 4488 8520 4988 8548
rect 4488 8508 4494 8520
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 5077 8551 5135 8557
rect 5077 8517 5089 8551
rect 5123 8548 5135 8551
rect 6825 8551 6883 8557
rect 5123 8520 6684 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 4522 8480 4528 8492
rect 3660 8452 4528 8480
rect 3660 8440 3666 8452
rect 4522 8440 4528 8452
rect 4580 8480 4586 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4580 8452 4629 8480
rect 4580 8440 4586 8452
rect 4617 8449 4629 8452
rect 4663 8480 4675 8483
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 4663 8452 5641 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 6656 8480 6684 8520
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 6914 8548 6920 8560
rect 6871 8520 6920 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 10318 8548 10324 8560
rect 9640 8520 10324 8548
rect 9640 8508 9646 8520
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 11992 8548 12020 8588
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12250 8616 12256 8628
rect 12115 8588 12256 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12492 8588 12537 8616
rect 12492 8576 12498 8588
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 14700 8588 15853 8616
rect 14700 8576 14706 8588
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 18966 8616 18972 8628
rect 16899 8588 18972 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 12526 8548 12532 8560
rect 11992 8520 12532 8548
rect 12526 8508 12532 8520
rect 12584 8548 12590 8560
rect 14826 8548 14832 8560
rect 12584 8520 13492 8548
rect 14787 8520 14832 8548
rect 12584 8508 12590 8520
rect 13464 8492 13492 8520
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 19610 8508 19616 8560
rect 19668 8548 19674 8560
rect 19978 8548 19984 8560
rect 19668 8520 19984 8548
rect 19668 8508 19674 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 7374 8480 7380 8492
rect 6656 8452 7380 8480
rect 5629 8443 5687 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7558 8480 7564 8492
rect 7515 8452 7564 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9548 8452 10824 8480
rect 9548 8440 9554 8452
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 5445 8415 5503 8421
rect 5445 8412 5457 8415
rect 3936 8384 5457 8412
rect 3936 8372 3942 8384
rect 5445 8381 5457 8384
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5592 8384 5637 8412
rect 5592 8372 5598 8384
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6788 8384 7297 8412
rect 6788 8372 6794 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 8110 8412 8116 8424
rect 8071 8384 8116 8412
rect 7285 8375 7343 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8570 8412 8576 8424
rect 8527 8384 8576 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 10226 8412 10232 8424
rect 8680 8384 10232 8412
rect 2124 8347 2182 8353
rect 2124 8313 2136 8347
rect 2170 8344 2182 8347
rect 2590 8344 2596 8356
rect 2170 8316 2596 8344
rect 2170 8313 2182 8316
rect 2124 8307 2182 8313
rect 2590 8304 2596 8316
rect 2648 8304 2654 8356
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6512 8316 7205 8344
rect 6512 8304 6518 8316
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 7193 8307 7251 8313
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8680 8344 8708 8384
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10686 8412 10692 8424
rect 10647 8384 10692 8412
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10796 8412 10824 8452
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12710 8480 12716 8492
rect 12308 8452 12716 8480
rect 12308 8440 12314 8452
rect 12710 8440 12716 8452
rect 12768 8480 12774 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12768 8452 13001 8480
rect 12768 8440 12774 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 13446 8480 13452 8492
rect 13359 8452 13452 8480
rect 12989 8443 13047 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 16390 8480 16396 8492
rect 16351 8452 16396 8480
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17543 8452 18184 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 10796 8384 12817 8412
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13648 8384 16160 8412
rect 8251 8316 8708 8344
rect 8748 8347 8806 8353
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8748 8313 8760 8347
rect 8794 8344 8806 8347
rect 9214 8344 9220 8356
rect 8794 8316 9220 8344
rect 8794 8313 8806 8316
rect 8748 8307 8806 8313
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 10956 8347 11014 8353
rect 10956 8344 10968 8347
rect 9456 8316 10968 8344
rect 9456 8304 9462 8316
rect 10956 8313 10968 8316
rect 11002 8344 11014 8347
rect 11330 8344 11336 8356
rect 11002 8316 11336 8344
rect 11002 8313 11014 8316
rect 10956 8307 11014 8313
rect 11330 8304 11336 8316
rect 11388 8344 11394 8356
rect 11882 8344 11888 8356
rect 11388 8316 11888 8344
rect 11388 8304 11394 8316
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 13648 8344 13676 8384
rect 11992 8316 13676 8344
rect 13716 8347 13774 8353
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4525 8279 4583 8285
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 4890 8276 4896 8288
rect 4571 8248 4896 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 6270 8276 6276 8288
rect 6231 8248 6276 8276
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 11992 8276 12020 8316
rect 13716 8313 13728 8347
rect 13762 8344 13774 8347
rect 13998 8344 14004 8356
rect 13762 8316 14004 8344
rect 13762 8313 13774 8316
rect 13716 8307 13774 8313
rect 13998 8304 14004 8316
rect 14056 8344 14062 8356
rect 14274 8344 14280 8356
rect 14056 8316 14280 8344
rect 14056 8304 14062 8316
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 16132 8344 16160 8384
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 16264 8384 16313 8412
rect 16264 8372 16270 8384
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16669 8415 16727 8421
rect 16669 8381 16681 8415
rect 16715 8412 16727 8415
rect 17678 8412 17684 8424
rect 16715 8384 17684 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 18012 8384 18061 8412
rect 18012 8372 18018 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18156 8412 18184 8452
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 19852 8452 20269 8480
rect 19852 8440 19858 8452
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 18305 8415 18363 8421
rect 18305 8412 18317 8415
rect 18156 8384 18317 8412
rect 18049 8375 18107 8381
rect 18305 8381 18317 8384
rect 18351 8412 18363 8415
rect 18690 8412 18696 8424
rect 18351 8384 18696 8412
rect 18351 8381 18363 8384
rect 18305 8375 18363 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 20165 8415 20223 8421
rect 20165 8412 20177 8415
rect 19300 8384 20177 8412
rect 19300 8372 19306 8384
rect 20165 8381 20177 8384
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8412 20775 8415
rect 20806 8412 20812 8424
rect 20763 8384 20812 8412
rect 20763 8381 20775 8384
rect 20717 8375 20775 8381
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 18506 8344 18512 8356
rect 16132 8316 18512 8344
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 18656 8316 20085 8344
rect 18656 8304 18662 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 7524 8248 12020 8276
rect 7524 8236 7530 8248
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 12952 8248 12997 8276
rect 12952 8236 12958 8248
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13630 8276 13636 8288
rect 13320 8248 13636 8276
rect 13320 8236 13326 8248
rect 13630 8236 13636 8248
rect 13688 8276 13694 8288
rect 16114 8276 16120 8288
rect 13688 8248 16120 8276
rect 13688 8236 13694 8248
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 16209 8279 16267 8285
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16669 8279 16727 8285
rect 16669 8276 16681 8279
rect 16255 8248 16681 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16669 8245 16681 8248
rect 16715 8245 16727 8279
rect 17218 8276 17224 8288
rect 17179 8248 17224 8276
rect 16669 8239 16727 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 17368 8248 17413 8276
rect 17368 8236 17374 8248
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20901 8279 20959 8285
rect 20901 8276 20913 8279
rect 20036 8248 20913 8276
rect 20036 8236 20042 8248
rect 20901 8245 20913 8248
rect 20947 8245 20959 8279
rect 20901 8239 20959 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2222 8072 2228 8084
rect 1995 8044 2228 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3786 8072 3792 8084
rect 3375 8044 3792 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4212 8044 4261 8072
rect 4212 8032 4218 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4982 8072 4988 8084
rect 4249 8035 4307 8041
rect 4356 8044 4988 8072
rect 3421 8007 3479 8013
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 4356 8004 4384 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6656 8044 6837 8072
rect 3467 7976 4384 8004
rect 4617 8007 4675 8013
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 4798 8004 4804 8016
rect 4663 7976 4804 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 5166 7964 5172 8016
rect 5224 8004 5230 8016
rect 5224 7976 5856 8004
rect 5224 7964 5230 7976
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2682 7936 2688 7948
rect 2363 7908 2688 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 5626 7936 5632 7948
rect 4580 7908 4844 7936
rect 5587 7908 5632 7936
rect 4580 7896 4586 7908
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2280 7840 2421 7868
rect 2280 7828 2286 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2590 7868 2596 7880
rect 2503 7840 2596 7868
rect 2409 7831 2467 7837
rect 2424 7800 2452 7831
rect 2590 7828 2596 7840
rect 2648 7868 2654 7880
rect 3602 7868 3608 7880
rect 2648 7840 3608 7868
rect 2648 7828 2654 7840
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4614 7868 4620 7880
rect 4212 7840 4620 7868
rect 4212 7828 4218 7840
rect 4614 7828 4620 7840
rect 4672 7868 4678 7880
rect 4816 7877 4844 7908
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4672 7840 4721 7868
rect 4672 7828 4678 7840
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 4801 7831 4859 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5828 7877 5856 7976
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 6656 8004 6684 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7432 8044 7941 8072
rect 7432 8032 7438 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 8987 8044 9873 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 10226 8072 10232 8084
rect 10187 8044 10232 8072
rect 9861 8035 9919 8041
rect 6328 7976 6684 8004
rect 8588 8004 8616 8035
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 11149 8075 11207 8081
rect 10376 8044 10421 8072
rect 10376 8032 10382 8044
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11422 8072 11428 8084
rect 11195 8044 11428 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 12066 8072 12072 8084
rect 11563 8044 12072 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12621 8075 12679 8081
rect 12621 8041 12633 8075
rect 12667 8072 12679 8075
rect 12894 8072 12900 8084
rect 12667 8044 12900 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13081 8075 13139 8081
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13127 8044 13553 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13906 8072 13912 8084
rect 13679 8044 13912 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 13998 8032 14004 8084
rect 14056 8072 14062 8084
rect 16482 8072 16488 8084
rect 14056 8044 14101 8072
rect 14660 8044 16488 8072
rect 14056 8032 14062 8044
rect 9950 8004 9956 8016
rect 8588 7976 9956 8004
rect 6328 7964 6334 7976
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 10962 7964 10968 8016
rect 11020 8004 11026 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 11020 7976 11897 8004
rect 11020 7964 11026 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 14660 8004 14688 8044
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 18690 8072 18696 8084
rect 18651 8044 18696 8072
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 15746 8004 15752 8016
rect 12400 7976 14688 8004
rect 14752 7976 15752 8004
rect 12400 7964 12406 7976
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 5920 7908 7849 7936
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 2866 7800 2872 7812
rect 2424 7772 2872 7800
rect 2866 7760 2872 7772
rect 2924 7760 2930 7812
rect 2961 7803 3019 7809
rect 2961 7769 2973 7803
rect 3007 7800 3019 7803
rect 5920 7800 5948 7908
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 10042 7936 10048 7948
rect 8536 7908 10048 7936
rect 8536 7896 8542 7908
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 11054 7936 11060 7948
rect 11015 7908 11060 7936
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 12989 7939 13047 7945
rect 11388 7908 12204 7936
rect 11388 7896 11394 7908
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 3007 7772 5948 7800
rect 6003 7840 6929 7868
rect 3007 7769 3019 7772
rect 2961 7763 3019 7769
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 6003 7732 6031 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 6454 7800 6460 7812
rect 6415 7772 6460 7800
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7024 7800 7052 7831
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7708 7840 8033 7868
rect 7708 7828 7714 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7837 9091 7871
rect 9214 7868 9220 7880
rect 9175 7840 9220 7868
rect 9033 7831 9091 7837
rect 6880 7772 7052 7800
rect 6880 7760 6886 7772
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 9048 7800 9076 7831
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 10226 7868 10232 7880
rect 9539 7840 10232 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10410 7868 10416 7880
rect 10371 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7868 10474 7880
rect 12176 7877 12204 7908
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 14752 7936 14780 7976
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 15930 8013 15936 8016
rect 15924 8004 15936 8013
rect 15891 7976 15936 8004
rect 15924 7967 15936 7976
rect 15930 7964 15936 7967
rect 15988 7964 15994 8016
rect 16758 7964 16764 8016
rect 16816 8004 16822 8016
rect 17558 8007 17616 8013
rect 17558 8004 17570 8007
rect 16816 7976 17570 8004
rect 16816 7964 16822 7976
rect 17558 7973 17570 7976
rect 17604 7973 17616 8007
rect 17558 7967 17616 7973
rect 13035 7908 14780 7936
rect 14829 7939 14887 7945
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 14829 7905 14841 7939
rect 14875 7936 14887 7939
rect 15010 7936 15016 7948
rect 14875 7908 15016 7936
rect 14875 7905 14887 7908
rect 14829 7899 14887 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15344 7908 15669 7936
rect 15344 7896 15350 7908
rect 15657 7905 15669 7908
rect 15703 7936 15715 7939
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 15703 7908 17325 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 17313 7905 17325 7908
rect 17359 7936 17371 7939
rect 17954 7936 17960 7948
rect 17359 7908 17960 7936
rect 17359 7905 17371 7908
rect 17313 7899 17371 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 20070 7936 20076 7948
rect 20031 7908 20076 7936
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 10468 7840 11253 7868
rect 10468 7828 10474 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11241 7831 11299 7837
rect 11339 7840 11989 7868
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 7248 7772 8984 7800
rect 9048 7772 10701 7800
rect 7248 7760 7254 7772
rect 2740 7704 6031 7732
rect 2740 7692 2746 7704
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 6604 7704 7481 7732
rect 6604 7692 6610 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 8956 7732 8984 7772
rect 10689 7769 10701 7772
rect 10735 7769 10747 7803
rect 10689 7763 10747 7769
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8956 7704 9505 7732
rect 7469 7695 7527 7701
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 10502 7692 10508 7744
rect 10560 7732 10566 7744
rect 11339 7732 11367 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7868 12219 7871
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12207 7840 13185 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13173 7831 13231 7837
rect 13280 7840 14105 7868
rect 11422 7760 11428 7812
rect 11480 7800 11486 7812
rect 11698 7800 11704 7812
rect 11480 7772 11704 7800
rect 11480 7760 11486 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 13280 7800 13308 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14093 7831 14151 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19116 7840 19257 7868
rect 19116 7828 19122 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 20162 7868 20168 7880
rect 20123 7840 20168 7868
rect 19245 7831 19303 7837
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 11848 7772 13308 7800
rect 13541 7803 13599 7809
rect 11848 7760 11854 7772
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14918 7800 14924 7812
rect 13587 7772 14924 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 19886 7800 19892 7812
rect 18748 7772 19892 7800
rect 18748 7760 18754 7772
rect 19886 7760 19892 7772
rect 19944 7800 19950 7812
rect 20272 7800 20300 7831
rect 19944 7772 20300 7800
rect 19944 7760 19950 7772
rect 10560 7704 11367 7732
rect 11716 7732 11744 7760
rect 12342 7732 12348 7744
rect 11716 7704 12348 7732
rect 10560 7692 10566 7704
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 15010 7732 15016 7744
rect 14691 7704 15016 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 17034 7732 17040 7744
rect 16995 7704 17040 7732
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 19702 7732 19708 7744
rect 19663 7704 19708 7732
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5350 7528 5356 7540
rect 4939 7500 5356 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6270 7528 6276 7540
rect 5960 7500 6276 7528
rect 5960 7488 5966 7500
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 8386 7528 8392 7540
rect 6696 7500 8392 7528
rect 6696 7488 6702 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9272 7500 9965 7528
rect 9272 7488 9278 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1544 7432 3832 7460
rect 1544 7420 1550 7432
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3510 7392 3516 7404
rect 2823 7364 3516 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 3804 7324 3832 7432
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4120 7432 8340 7460
rect 4120 7420 4126 7432
rect 3970 7392 3976 7404
rect 3931 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5224 7364 5457 7392
rect 5224 7352 5230 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 7466 7392 7472 7404
rect 5445 7355 5503 7361
rect 7024 7364 7236 7392
rect 7427 7364 7472 7392
rect 7024 7324 7052 7364
rect 7208 7333 7236 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 3804 7296 7052 7324
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7650 7324 7656 7336
rect 7239 7296 7656 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 8202 7324 8208 7336
rect 8067 7296 8208 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8312 7324 8340 7432
rect 9968 7392 9996 7491
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 10192 7500 10241 7528
rect 10192 7488 10198 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 15102 7528 15108 7540
rect 10229 7491 10287 7497
rect 10336 7500 14780 7528
rect 15063 7500 15108 7528
rect 10045 7463 10103 7469
rect 10045 7429 10057 7463
rect 10091 7460 10103 7463
rect 10336 7460 10364 7500
rect 10091 7432 10364 7460
rect 10091 7429 10103 7432
rect 10045 7423 10103 7429
rect 11900 7404 11928 7500
rect 13078 7420 13084 7472
rect 13136 7460 13142 7472
rect 13136 7432 13216 7460
rect 13136 7420 13142 7432
rect 10781 7395 10839 7401
rect 10781 7392 10793 7395
rect 9968 7364 10793 7392
rect 10781 7361 10793 7364
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 8573 7327 8631 7333
rect 8312 7296 8432 7324
rect 3878 7256 3884 7268
rect 3839 7228 3884 7256
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 8404 7256 8432 7296
rect 8573 7293 8585 7327
rect 8619 7324 8631 7327
rect 8662 7324 8668 7336
rect 8619 7296 8668 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8840 7327 8898 7333
rect 8840 7293 8852 7327
rect 8886 7324 8898 7327
rect 10410 7324 10416 7336
rect 8886 7296 10416 7324
rect 8886 7293 8898 7296
rect 8840 7287 8898 7293
rect 10410 7284 10416 7296
rect 10468 7324 10474 7336
rect 11808 7324 11836 7355
rect 11882 7352 11888 7404
rect 11940 7352 11946 7404
rect 13188 7401 13216 7432
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13173 7355 13231 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13504 7364 13737 7392
rect 13504 7352 13510 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 10468 7296 11836 7324
rect 13081 7327 13139 7333
rect 10468 7284 10474 7296
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13127 7296 13645 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 14752 7324 14780 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 17218 7528 17224 7540
rect 16255 7500 17224 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 17586 7460 17592 7472
rect 16408 7432 17592 7460
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 16408 7392 16436 7432
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 20714 7460 20720 7472
rect 20180 7432 20720 7460
rect 16758 7392 16764 7404
rect 14976 7364 16436 7392
rect 16719 7364 16764 7392
rect 14976 7352 14982 7364
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 18690 7352 18696 7404
rect 18748 7392 18754 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 18748 7364 19257 7392
rect 18748 7352 18754 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 16577 7327 16635 7333
rect 16577 7324 16589 7327
rect 14752 7296 16589 7324
rect 13633 7287 13691 7293
rect 16577 7293 16589 7296
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 19058 7324 19064 7336
rect 16724 7296 16769 7324
rect 19019 7296 19064 7324
rect 16724 7284 16730 7296
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 20073 7327 20131 7333
rect 19668 7296 19840 7324
rect 19668 7284 19674 7296
rect 10962 7256 10968 7268
rect 5399 7228 8340 7256
rect 8404 7228 10968 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 2004 7160 2513 7188
rect 2004 7148 2010 7160
rect 2501 7157 2513 7160
rect 2547 7157 2559 7191
rect 2501 7151 2559 7157
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 3050 7188 3056 7200
rect 2639 7160 3056 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3786 7188 3792 7200
rect 3747 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 5040 7160 5273 7188
rect 5040 7148 5046 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 5592 7160 6837 7188
rect 5592 7148 5598 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 7248 7160 7297 7188
rect 7248 7148 7254 7160
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 7285 7151 7343 7157
rect 7837 7191 7895 7197
rect 7837 7157 7849 7191
rect 7883 7188 7895 7191
rect 8202 7188 8208 7200
rect 7883 7160 8208 7188
rect 7883 7157 7895 7160
rect 7837 7151 7895 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 8312 7188 8340 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 11974 7256 11980 7268
rect 11747 7228 11980 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 11974 7216 11980 7228
rect 12032 7216 12038 7268
rect 13998 7265 14004 7268
rect 13992 7219 14004 7265
rect 14056 7256 14062 7268
rect 15470 7256 15476 7268
rect 14056 7228 14092 7256
rect 15120 7228 15476 7256
rect 13998 7216 14004 7219
rect 14056 7216 14062 7228
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 8312 7160 10057 7188
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10594 7188 10600 7200
rect 10555 7160 10600 7188
rect 10045 7151 10103 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 10735 7160 11253 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 11514 7148 11520 7200
rect 11572 7188 11578 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 11572 7160 11621 7188
rect 11572 7148 11578 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 11609 7151 11667 7157
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12676 7160 12725 7188
rect 12676 7148 12682 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 12713 7151 12771 7157
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 13078 7188 13084 7200
rect 12860 7160 13084 7188
rect 12860 7148 12866 7160
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 15120 7188 15148 7228
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 15378 7188 15384 7200
rect 13679 7160 15148 7188
rect 15339 7160 15384 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 18233 7191 18291 7197
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 18506 7188 18512 7200
rect 18279 7160 18512 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 18690 7188 18696 7200
rect 18651 7160 18696 7188
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 19153 7191 19211 7197
rect 19153 7157 19165 7191
rect 19199 7188 19211 7191
rect 19705 7191 19763 7197
rect 19705 7188 19717 7191
rect 19199 7160 19717 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 19705 7157 19717 7160
rect 19751 7157 19763 7191
rect 19812 7188 19840 7296
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 20180 7324 20208 7432
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7392 20407 7395
rect 20622 7392 20628 7404
rect 20395 7364 20628 7392
rect 20395 7361 20407 7364
rect 20349 7355 20407 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20714 7324 20720 7336
rect 20119 7296 20208 7324
rect 20675 7296 20720 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19812 7160 20177 7188
rect 19705 7151 19763 7157
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 20165 7151 20223 7157
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20901 7191 20959 7197
rect 20901 7188 20913 7191
rect 20312 7160 20913 7188
rect 20312 7148 20318 7160
rect 20901 7157 20913 7160
rect 20947 7157 20959 7191
rect 20901 7151 20959 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 4120 6956 6929 6984
rect 4120 6944 4126 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 9953 6987 10011 6993
rect 6917 6947 6975 6953
rect 7668 6956 9076 6984
rect 4976 6919 5034 6925
rect 4976 6885 4988 6919
rect 5022 6916 5034 6919
rect 7466 6916 7472 6928
rect 5022 6888 7472 6916
rect 5022 6885 5034 6888
rect 4976 6879 5034 6885
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 1912 6820 2145 6848
rect 1912 6808 1918 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 2133 6811 2191 6817
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 2866 6848 2872 6860
rect 2446 6820 2872 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 6822 6848 6828 6860
rect 6783 6820 6828 6848
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7668 6848 7696 6956
rect 9048 6916 9076 6956
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10594 6984 10600 6996
rect 9999 6956 10600 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13170 6984 13176 6996
rect 12492 6956 13176 6984
rect 12492 6944 12498 6956
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13541 6987 13599 6993
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 15378 6984 15384 6996
rect 13587 6956 15384 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15804 6956 16037 6984
rect 15804 6944 15810 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 16025 6947 16083 6953
rect 16117 6987 16175 6993
rect 16117 6953 16129 6987
rect 16163 6984 16175 6987
rect 16298 6984 16304 6996
rect 16163 6956 16304 6984
rect 16163 6953 16175 6956
rect 16117 6947 16175 6953
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 17310 6984 17316 6996
rect 16715 6956 17316 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 17681 6987 17739 6993
rect 17681 6953 17693 6987
rect 17727 6984 17739 6987
rect 17954 6984 17960 6996
rect 17727 6956 17960 6984
rect 17727 6953 17739 6956
rect 17681 6947 17739 6953
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 18598 6984 18604 6996
rect 18559 6956 18604 6984
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 18969 6987 19027 6993
rect 18969 6984 18981 6987
rect 18748 6956 18981 6984
rect 18748 6944 18754 6956
rect 18969 6953 18981 6956
rect 19015 6953 19027 6987
rect 18969 6947 19027 6953
rect 19058 6944 19064 6996
rect 19116 6984 19122 6996
rect 19981 6987 20039 6993
rect 19981 6984 19993 6987
rect 19116 6956 19993 6984
rect 19116 6944 19122 6956
rect 19981 6953 19993 6956
rect 20027 6953 20039 6987
rect 19981 6947 20039 6953
rect 7024 6820 7696 6848
rect 7760 6888 8984 6916
rect 9048 6888 9996 6916
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 4724 6644 4752 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 7024 6780 7052 6820
rect 5776 6752 7052 6780
rect 7101 6783 7159 6789
rect 5776 6740 5782 6752
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7190 6780 7196 6792
rect 7147 6752 7196 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7190 6740 7196 6752
rect 7248 6780 7254 6792
rect 7760 6780 7788 6888
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6817 7895 6851
rect 8846 6848 8852 6860
rect 8807 6820 8852 6848
rect 7837 6811 7895 6817
rect 7248 6752 7788 6780
rect 7248 6740 7254 6752
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6712 6515 6715
rect 7852 6712 7880 6811
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 8956 6848 8984 6888
rect 9968 6848 9996 6888
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 10100 6888 10333 6916
rect 10100 6876 10106 6888
rect 10321 6885 10333 6888
rect 10367 6885 10379 6919
rect 17037 6919 17095 6925
rect 17037 6916 17049 6919
rect 10321 6879 10379 6885
rect 10428 6888 17049 6916
rect 10428 6848 10456 6888
rect 17037 6885 17049 6888
rect 17083 6885 17095 6919
rect 17037 6879 17095 6885
rect 17497 6919 17555 6925
rect 17497 6885 17509 6919
rect 17543 6916 17555 6919
rect 20073 6919 20131 6925
rect 20073 6916 20085 6919
rect 17543 6888 20085 6916
rect 17543 6885 17555 6888
rect 17497 6879 17555 6885
rect 20073 6885 20085 6888
rect 20119 6885 20131 6919
rect 20073 6879 20131 6885
rect 8956 6820 9076 6848
rect 9968 6820 10456 6848
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8294 6780 8300 6792
rect 8159 6752 8300 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 6503 6684 7880 6712
rect 7944 6712 7972 6743
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9048 6789 9076 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10962 6848 10968 6860
rect 10744 6820 10968 6848
rect 10744 6808 10750 6820
rect 10962 6808 10968 6820
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11324 6851 11382 6857
rect 11324 6817 11336 6851
rect 11370 6848 11382 6851
rect 12986 6848 12992 6860
rect 11370 6820 12992 6848
rect 11370 6817 11382 6820
rect 11324 6811 11382 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 13188 6820 14565 6848
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6780 9091 6783
rect 9490 6780 9496 6792
rect 9079 6752 9496 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10008 6752 10425 6780
rect 10008 6740 10014 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 12710 6780 12716 6792
rect 10560 6752 10605 6780
rect 12671 6752 12716 6780
rect 10560 6740 10566 6752
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 7944 6684 8493 6712
rect 6503 6681 6515 6684
rect 6457 6675 6515 6681
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 10042 6712 10048 6724
rect 9732 6684 10048 6712
rect 9732 6672 9738 6684
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 13188 6721 13216 6820
rect 14553 6817 14565 6820
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15378 6848 15384 6860
rect 15252 6820 15384 6848
rect 15252 6808 15258 6820
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 17126 6848 17132 6860
rect 17087 6820 17132 6848
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 13630 6780 13636 6792
rect 13591 6752 13636 6780
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 13998 6780 14004 6792
rect 13771 6752 14004 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14366 6740 14372 6792
rect 14424 6780 14430 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14424 6752 14657 6780
rect 14424 6740 14430 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15102 6780 15108 6792
rect 14875 6752 15108 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16758 6780 16764 6792
rect 16347 6752 16764 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16758 6740 16764 6752
rect 16816 6780 16822 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 16816 6752 17325 6780
rect 16816 6740 16822 6752
rect 17313 6749 17325 6752
rect 17359 6780 17371 6783
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17359 6752 17601 6780
rect 17359 6749 17371 6752
rect 17313 6743 17371 6749
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6681 13231 6715
rect 13173 6675 13231 6681
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 15010 6712 15016 6724
rect 14332 6684 15016 6712
rect 14332 6672 14338 6684
rect 15010 6672 15016 6684
rect 15068 6712 15074 6724
rect 17880 6712 17908 6811
rect 17954 6808 17960 6860
rect 18012 6848 18018 6860
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 18012 6820 18061 6848
rect 18012 6808 18018 6820
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 19024 6820 19073 6848
rect 19024 6808 19030 6820
rect 19061 6817 19073 6820
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6780 19303 6783
rect 19426 6780 19432 6792
rect 19291 6752 19432 6780
rect 19291 6749 19303 6752
rect 19245 6743 19303 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 20165 6783 20223 6789
rect 20165 6780 20177 6783
rect 19944 6752 20177 6780
rect 19944 6740 19950 6752
rect 20165 6749 20177 6752
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 15068 6684 17908 6712
rect 18233 6715 18291 6721
rect 15068 6672 15074 6684
rect 18233 6681 18245 6715
rect 18279 6712 18291 6715
rect 18874 6712 18880 6724
rect 18279 6684 18880 6712
rect 18279 6681 18291 6684
rect 18233 6675 18291 6681
rect 18874 6672 18880 6684
rect 18932 6672 18938 6724
rect 20622 6712 20628 6724
rect 18984 6684 20628 6712
rect 5350 6644 5356 6656
rect 4724 6616 5356 6644
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5500 6616 6101 6644
rect 5500 6604 5506 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 8938 6644 8944 6656
rect 7515 6616 8944 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 12250 6644 12256 6656
rect 9364 6616 12256 6644
rect 9364 6604 9370 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12400 6616 12449 6644
rect 12400 6604 12406 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 15194 6644 15200 6656
rect 14231 6616 15200 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15657 6647 15715 6653
rect 15657 6613 15669 6647
rect 15703 6644 15715 6647
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 15703 6616 17509 6644
rect 15703 6613 15715 6616
rect 15657 6607 15715 6613
rect 17497 6613 17509 6616
rect 17543 6613 17555 6647
rect 17497 6607 17555 6613
rect 17589 6647 17647 6653
rect 17589 6613 17601 6647
rect 17635 6644 17647 6647
rect 18984 6644 19012 6684
rect 20622 6672 20628 6684
rect 20680 6672 20686 6724
rect 19610 6644 19616 6656
rect 17635 6616 19012 6644
rect 19571 6616 19616 6644
rect 17635 6613 17647 6616
rect 17589 6607 17647 6613
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3108 6412 3341 6440
rect 3108 6400 3114 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3329 6403 3387 6409
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6788 6412 6837 6440
rect 6788 6400 6794 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7466 6440 7472 6452
rect 7156 6412 7472 6440
rect 7156 6400 7162 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 11241 6443 11299 6449
rect 11241 6440 11253 6443
rect 10560 6412 11253 6440
rect 10560 6400 10566 6412
rect 11241 6409 11253 6412
rect 11287 6409 11299 6443
rect 11241 6403 11299 6409
rect 11900 6412 12204 6440
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 9582 6372 9588 6384
rect 3844 6344 4016 6372
rect 9543 6344 9588 6372
rect 3844 6332 3850 6344
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3050 6304 3056 6316
rect 2924 6276 3056 6304
rect 2924 6264 2930 6276
rect 3050 6264 3056 6276
rect 3108 6304 3114 6316
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 3108 6276 3893 6304
rect 3108 6264 3114 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1762 6236 1768 6248
rect 1719 6208 1768 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3476 6208 3709 6236
rect 3476 6196 3482 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 1940 6171 1998 6177
rect 1940 6137 1952 6171
rect 1986 6168 1998 6171
rect 2498 6168 2504 6180
rect 1986 6140 2504 6168
rect 1986 6137 1998 6140
rect 1940 6131 1998 6137
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 3988 6168 4016 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 11900 6372 11928 6412
rect 11020 6344 11928 6372
rect 11977 6375 12035 6381
rect 11020 6332 11026 6344
rect 11977 6341 11989 6375
rect 12023 6372 12035 6375
rect 12066 6372 12072 6384
rect 12023 6344 12072 6372
rect 12023 6341 12035 6344
rect 11977 6335 12035 6341
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 12176 6372 12204 6412
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12308 6412 13400 6440
rect 12308 6400 12314 6412
rect 13372 6372 13400 6412
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 15010 6440 15016 6452
rect 14056 6412 15016 6440
rect 14056 6400 14062 6412
rect 15010 6400 15016 6412
rect 15068 6440 15074 6452
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 15068 6412 15761 6440
rect 15068 6400 15074 6412
rect 15749 6409 15761 6412
rect 15795 6409 15807 6443
rect 15749 6403 15807 6409
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 19150 6440 19156 6452
rect 17635 6412 19156 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 20530 6440 20536 6452
rect 20211 6412 20536 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 13817 6375 13875 6381
rect 12176 6344 12480 6372
rect 13372 6344 13492 6372
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 5442 6304 5448 6316
rect 4212 6276 5448 6304
rect 4212 6264 4218 6276
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 6822 6304 6828 6316
rect 6319 6276 6828 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6972 6276 7481 6304
rect 6972 6264 6978 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 7742 6304 7748 6316
rect 7515 6276 7748 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 9600 6304 9628 6332
rect 12452 6316 12480 6344
rect 9600 6276 9996 6304
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5534 6236 5540 6248
rect 5399 6208 5540 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 8110 6236 8116 6248
rect 6135 6208 8116 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8754 6236 8760 6248
rect 8251 6208 8760 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8754 6196 8760 6208
rect 8812 6236 8818 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 8812 6208 9873 6236
rect 8812 6196 8818 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9968 6236 9996 6276
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 12434 6304 12440 6316
rect 11204 6276 12204 6304
rect 12347 6276 12440 6304
rect 11204 6264 11210 6276
rect 10117 6239 10175 6245
rect 10117 6236 10129 6239
rect 9968 6208 10129 6236
rect 9861 6199 9919 6205
rect 10117 6205 10129 6208
rect 10163 6205 10175 6239
rect 10117 6199 10175 6205
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11698 6236 11704 6248
rect 11112 6208 11704 6236
rect 11112 6196 11118 6208
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 7193 6171 7251 6177
rect 7193 6168 7205 6171
rect 3988 6140 7205 6168
rect 7193 6137 7205 6140
rect 7239 6137 7251 6171
rect 7193 6131 7251 6137
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8450 6171 8508 6177
rect 8450 6168 8462 6171
rect 8352 6140 8462 6168
rect 8352 6128 8358 6140
rect 8450 6137 8462 6140
rect 8496 6137 8508 6171
rect 8450 6131 8508 6137
rect 10226 6128 10232 6180
rect 10284 6168 10290 6180
rect 10410 6168 10416 6180
rect 10284 6140 10416 6168
rect 10284 6128 10290 6140
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 11808 6168 11836 6199
rect 12176 6168 12204 6276
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 13464 6304 13492 6344
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 13909 6375 13967 6381
rect 13909 6372 13921 6375
rect 13863 6344 13921 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 13909 6341 13921 6344
rect 13955 6341 13967 6375
rect 13909 6335 13967 6341
rect 16025 6375 16083 6381
rect 16025 6341 16037 6375
rect 16071 6372 16083 6375
rect 16071 6344 18460 6372
rect 16071 6341 16083 6344
rect 16025 6335 16083 6341
rect 16669 6307 16727 6313
rect 13464 6276 14504 6304
rect 12452 6236 12480 6264
rect 13262 6236 13268 6248
rect 12452 6208 13268 6236
rect 13262 6196 13268 6208
rect 13320 6236 13326 6248
rect 14274 6236 14280 6248
rect 13320 6208 14035 6236
rect 14235 6208 14280 6236
rect 13320 6196 13326 6208
rect 12342 6168 12348 6180
rect 11808 6140 12112 6168
rect 12176 6140 12348 6168
rect 3050 6100 3056 6112
rect 3011 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 3835 6072 4905 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 5902 6100 5908 6112
rect 5408 6072 5908 6100
rect 5408 6060 5414 6072
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 10594 6100 10600 6112
rect 7331 6072 10600 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 12084 6100 12112 6140
rect 12342 6128 12348 6140
rect 12400 6168 12406 6180
rect 12682 6171 12740 6177
rect 12682 6168 12694 6171
rect 12400 6140 12694 6168
rect 12400 6128 12406 6140
rect 12682 6137 12694 6140
rect 12728 6137 12740 6171
rect 12682 6131 12740 6137
rect 13354 6128 13360 6180
rect 13412 6168 13418 6180
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 13412 6140 13921 6168
rect 13412 6128 13418 6140
rect 13909 6137 13921 6140
rect 13955 6137 13967 6171
rect 13909 6131 13967 6137
rect 12802 6100 12808 6112
rect 12084 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 14007 6100 14035 6208
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14476 6236 14504 6276
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 17034 6304 17040 6316
rect 16715 6276 17040 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 16485 6239 16543 6245
rect 16485 6236 16497 6239
rect 14476 6208 16497 6236
rect 14369 6199 14427 6205
rect 16485 6205 16497 6208
rect 16531 6205 16543 6239
rect 17402 6236 17408 6248
rect 17363 6208 17408 6236
rect 16485 6199 16543 6205
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 14007 6072 14105 6100
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 14384 6100 14412 6199
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18432 6245 18460 6344
rect 18690 6304 18696 6316
rect 18651 6276 18696 6304
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19484 6276 19717 6304
rect 19484 6264 19490 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20717 6307 20775 6313
rect 20717 6304 20729 6307
rect 19852 6276 20729 6304
rect 19852 6264 19858 6276
rect 20717 6273 20729 6276
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 19610 6236 19616 6248
rect 19567 6208 19616 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 14636 6171 14694 6177
rect 14636 6137 14648 6171
rect 14682 6168 14694 6171
rect 15102 6168 15108 6180
rect 14682 6140 15108 6168
rect 14682 6137 14694 6140
rect 14636 6131 14694 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 16390 6168 16396 6180
rect 16351 6140 16396 6168
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 17218 6128 17224 6180
rect 17276 6168 17282 6180
rect 17954 6168 17960 6180
rect 17276 6140 17960 6168
rect 17276 6128 17282 6140
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 20625 6171 20683 6177
rect 20625 6168 20637 6171
rect 18064 6140 20637 6168
rect 15746 6100 15752 6112
rect 14384 6072 15752 6100
rect 14093 6063 14151 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 18064 6109 18092 6140
rect 20625 6137 20637 6140
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18874 6100 18880 6112
rect 18555 6072 18880 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 19153 6103 19211 6109
rect 19153 6069 19165 6103
rect 19199 6100 19211 6103
rect 19242 6100 19248 6112
rect 19199 6072 19248 6100
rect 19199 6069 19211 6072
rect 19153 6063 19211 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19613 6103 19671 6109
rect 19613 6069 19625 6103
rect 19659 6100 19671 6103
rect 19702 6100 19708 6112
rect 19659 6072 19708 6100
rect 19659 6069 19671 6072
rect 19613 6063 19671 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 20530 6100 20536 6112
rect 20491 6072 20536 6100
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2455 5868 2973 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3200 5868 3433 5896
rect 3200 5856 3206 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5316 5868 5917 5896
rect 5316 5856 5322 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 7098 5896 7104 5908
rect 5905 5859 5963 5865
rect 6840 5868 7104 5896
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 4310 5831 4368 5837
rect 4310 5828 4322 5831
rect 3568 5800 4322 5828
rect 3568 5788 3574 5800
rect 4310 5797 4322 5800
rect 4356 5797 4368 5831
rect 4310 5791 4368 5797
rect 2314 5760 2320 5772
rect 2275 5732 2320 5760
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2740 5732 3341 5760
rect 2740 5720 2746 5732
rect 3329 5729 3341 5732
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6730 5760 6736 5772
rect 6319 5732 6736 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2866 5692 2872 5704
rect 2639 5664 2872 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 3970 5692 3976 5704
rect 3559 5664 3976 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 3528 5624 3556 5655
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6454 5692 6460 5704
rect 6411 5664 6460 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 4080 5624 4108 5655
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6840 5692 6868 5868
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8938 5896 8944 5908
rect 8899 5868 8944 5896
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 11977 5899 12035 5905
rect 9048 5868 10272 5896
rect 9048 5828 9076 5868
rect 7944 5800 9076 5828
rect 7190 5769 7196 5772
rect 7184 5723 7196 5769
rect 7248 5760 7254 5772
rect 7248 5732 7284 5760
rect 7190 5720 7196 5723
rect 7248 5720 7254 5732
rect 6595 5664 6868 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 6972 5664 7017 5692
rect 6972 5652 6978 5664
rect 5902 5624 5908 5636
rect 2556 5596 3556 5624
rect 3988 5596 4108 5624
rect 5276 5596 5908 5624
rect 2556 5584 2562 5596
rect 3510 5516 3516 5568
rect 3568 5556 3574 5568
rect 3988 5556 4016 5596
rect 5276 5556 5304 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 5442 5556 5448 5568
rect 3568 5528 5304 5556
rect 5403 5528 5448 5556
rect 3568 5516 3574 5528
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 7944 5556 7972 5800
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 10244 5828 10272 5868
rect 11977 5865 11989 5899
rect 12023 5896 12035 5899
rect 12618 5896 12624 5908
rect 12023 5868 12624 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 17402 5896 17408 5908
rect 12820 5868 17408 5896
rect 12820 5828 12848 5868
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5865 17555 5899
rect 17497 5859 17555 5865
rect 17589 5899 17647 5905
rect 17589 5865 17601 5899
rect 17635 5896 17647 5899
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 17635 5868 19257 5896
rect 17635 5865 17647 5868
rect 17589 5859 17647 5865
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 19429 5899 19487 5905
rect 19429 5865 19441 5899
rect 19475 5896 19487 5899
rect 20530 5896 20536 5908
rect 19475 5868 20536 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 9548 5800 10180 5828
rect 10244 5800 12848 5828
rect 12888 5831 12946 5837
rect 9548 5788 9554 5800
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9858 5760 9864 5772
rect 9456 5732 9864 5760
rect 9456 5720 9462 5732
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10152 5760 10180 5800
rect 12888 5797 12900 5831
rect 12934 5828 12946 5831
rect 13354 5828 13360 5840
rect 12934 5800 13360 5828
rect 12934 5797 12946 5800
rect 12888 5791 12946 5797
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 16384 5831 16442 5837
rect 16384 5797 16396 5831
rect 16430 5828 16442 5831
rect 16850 5828 16856 5840
rect 16430 5800 16856 5828
rect 16430 5797 16442 5800
rect 16384 5791 16442 5797
rect 16850 5788 16856 5800
rect 16908 5828 16914 5840
rect 17034 5828 17040 5840
rect 16908 5800 17040 5828
rect 16908 5788 16914 5800
rect 17034 5788 17040 5800
rect 17092 5788 17098 5840
rect 17512 5828 17540 5859
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 18040 5831 18098 5837
rect 18040 5828 18052 5831
rect 17512 5800 18052 5828
rect 18040 5797 18052 5800
rect 18086 5828 18098 5831
rect 18690 5828 18696 5840
rect 18086 5800 18696 5828
rect 18086 5797 18098 5800
rect 18040 5791 18098 5797
rect 18690 5788 18696 5800
rect 18748 5828 18754 5840
rect 18748 5800 20024 5828
rect 18748 5788 18754 5800
rect 11057 5763 11115 5769
rect 10152 5732 10272 5760
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8628 5664 9045 5692
rect 8628 5652 8634 5664
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9582 5692 9588 5704
rect 9263 5664 9588 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10134 5692 10140 5704
rect 9824 5664 10140 5692
rect 9824 5652 9830 5664
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10244 5701 10272 5732
rect 11057 5729 11069 5763
rect 11103 5760 11115 5763
rect 11698 5760 11704 5772
rect 11103 5732 11704 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12434 5760 12440 5772
rect 12115 5732 12440 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12584 5732 12633 5760
rect 12584 5720 12590 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 14274 5760 14280 5772
rect 14235 5732 14280 5760
rect 12621 5723 12679 5729
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 15562 5760 15568 5772
rect 15523 5732 15568 5760
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15804 5732 16129 5760
rect 15804 5720 15810 5732
rect 16117 5729 16129 5732
rect 16163 5760 16175 5763
rect 16163 5732 17172 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 11790 5692 11796 5704
rect 10229 5655 10287 5661
rect 10336 5664 11796 5692
rect 9858 5624 9864 5636
rect 8588 5596 9864 5624
rect 8294 5556 8300 5568
rect 6512 5528 7972 5556
rect 8255 5528 8300 5556
rect 6512 5516 6518 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8588 5565 8616 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5525 8631 5559
rect 8573 5519 8631 5525
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9088 5528 9689 5556
rect 9088 5516 9094 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 9677 5519 9735 5525
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10226 5556 10232 5568
rect 9824 5528 10232 5556
rect 9824 5516 9830 5528
rect 10226 5516 10232 5528
rect 10284 5556 10290 5568
rect 10336 5556 10364 5664
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 17144 5692 17172 5732
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17368 5732 17601 5760
rect 17368 5720 17374 5732
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5760 17831 5763
rect 17862 5760 17868 5772
rect 17819 5732 17868 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 17788 5692 17816 5723
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 18564 5732 19809 5760
rect 18564 5720 18570 5732
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 19886 5692 19892 5704
rect 12299 5664 12664 5692
rect 17144 5664 17816 5692
rect 19847 5664 19892 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 11609 5627 11667 5633
rect 11609 5593 11621 5627
rect 11655 5624 11667 5627
rect 12526 5624 12532 5636
rect 11655 5596 12532 5624
rect 11655 5593 11667 5596
rect 11609 5587 11667 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 10284 5528 10364 5556
rect 11241 5559 11299 5565
rect 10284 5516 10290 5528
rect 11241 5525 11253 5559
rect 11287 5556 11299 5559
rect 12342 5556 12348 5568
rect 11287 5528 12348 5556
rect 11287 5525 11299 5528
rect 11241 5519 11299 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 12636 5556 12664 5664
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 19996 5701 20024 5800
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 19153 5627 19211 5633
rect 19153 5593 19165 5627
rect 19199 5624 19211 5627
rect 19245 5627 19303 5633
rect 19245 5624 19257 5627
rect 19199 5596 19257 5624
rect 19199 5593 19211 5596
rect 19153 5587 19211 5593
rect 19245 5593 19257 5596
rect 19291 5624 19303 5627
rect 19794 5624 19800 5636
rect 19291 5596 19800 5624
rect 19291 5593 19303 5596
rect 19245 5587 19303 5593
rect 19794 5584 19800 5596
rect 19852 5584 19858 5636
rect 13630 5556 13636 5568
rect 12636 5528 13636 5556
rect 13630 5516 13636 5528
rect 13688 5556 13694 5568
rect 14001 5559 14059 5565
rect 14001 5556 14013 5559
rect 13688 5528 14013 5556
rect 13688 5516 13694 5528
rect 14001 5525 14013 5528
rect 14047 5525 14059 5559
rect 14001 5519 14059 5525
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 15286 5556 15292 5568
rect 14507 5528 15292 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 16758 5556 16764 5568
rect 15795 5528 16764 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 17494 5516 17500 5568
rect 17552 5556 17558 5568
rect 19058 5556 19064 5568
rect 17552 5528 19064 5556
rect 17552 5516 17558 5528
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 2314 5352 2320 5364
rect 2087 5324 2320 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 7006 5352 7012 5364
rect 6236 5324 7012 5352
rect 6236 5312 6242 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 8570 5352 8576 5364
rect 8531 5324 8576 5352
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 11054 5352 11060 5364
rect 9968 5324 11060 5352
rect 4709 5287 4767 5293
rect 4709 5253 4721 5287
rect 4755 5284 4767 5287
rect 5902 5284 5908 5296
rect 4755 5256 5908 5284
rect 4755 5253 4767 5256
rect 4709 5247 4767 5253
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6549 5287 6607 5293
rect 6549 5253 6561 5287
rect 6595 5284 6607 5287
rect 6595 5256 7604 5284
rect 6595 5253 6607 5256
rect 6549 5247 6607 5253
rect 2498 5176 2504 5228
rect 2556 5216 2562 5228
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2556 5188 2605 5216
rect 2556 5176 2562 5188
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 5132 5188 5273 5216
rect 5132 5176 5138 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 6273 5219 6331 5225
rect 6273 5216 6285 5219
rect 5500 5188 6285 5216
rect 5500 5176 5506 5188
rect 6273 5185 6285 5188
rect 6319 5185 6331 5219
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 6273 5179 6331 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7576 5216 7604 5256
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8352 5256 9168 5284
rect 8352 5244 8358 5256
rect 9030 5216 9036 5228
rect 7576 5188 8892 5216
rect 8991 5188 9036 5216
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1728 5120 2421 5148
rect 1728 5108 1734 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4028 5120 8156 5148
rect 4028 5108 4034 5120
rect 5169 5083 5227 5089
rect 5169 5049 5181 5083
rect 5215 5080 5227 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 5215 5052 6561 5080
rect 5215 5049 5227 5052
rect 5169 5043 5227 5049
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 7156 5052 7297 5080
rect 7156 5040 7162 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 8128 5080 8156 5120
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8260 5120 8493 5148
rect 8260 5108 8266 5120
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8864 5148 8892 5188
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9140 5225 9168 5256
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9766 5148 9772 5160
rect 8864 5120 9772 5148
rect 8481 5111 8539 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 9968 5080 9996 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12492 5324 12909 5352
rect 12492 5312 12498 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14366 5352 14372 5364
rect 14323 5324 14372 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 17770 5352 17776 5364
rect 16540 5324 17776 5352
rect 16540 5312 16546 5324
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 21174 5352 21180 5364
rect 19208 5324 21180 5352
rect 19208 5312 19214 5324
rect 21174 5312 21180 5324
rect 21232 5312 21238 5364
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 12618 5284 12624 5296
rect 10091 5256 12624 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 18417 5287 18475 5293
rect 13412 5256 13492 5284
rect 13412 5244 13418 5256
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11146 5216 11152 5228
rect 10735 5188 11152 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 13464 5225 13492 5256
rect 18417 5253 18429 5287
rect 18463 5284 18475 5287
rect 18874 5284 18880 5296
rect 18463 5256 18880 5284
rect 18463 5253 18475 5256
rect 18417 5247 18475 5253
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11480 5188 11713 5216
rect 11480 5176 11486 5188
rect 11701 5185 11713 5188
rect 11747 5216 11759 5219
rect 13449 5219 13507 5225
rect 11747 5188 12296 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5148 10471 5151
rect 11790 5148 11796 5160
rect 10459 5120 11796 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12268 5148 12296 5188
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14148 5188 14749 5216
rect 14148 5176 14154 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15010 5216 15016 5228
rect 14967 5188 15016 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15470 5216 15476 5228
rect 15335 5188 15476 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 15746 5216 15752 5228
rect 15707 5188 15752 5216
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 16908 5188 18981 5216
rect 16908 5176 16914 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 19058 5176 19064 5228
rect 19116 5216 19122 5228
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 19116 5188 19625 5216
rect 19116 5176 19122 5188
rect 19613 5185 19625 5188
rect 19659 5185 19671 5219
rect 19613 5179 19671 5185
rect 16016 5151 16074 5157
rect 12268 5120 14780 5148
rect 8128 5052 9996 5080
rect 10505 5083 10563 5089
rect 7285 5043 7343 5049
rect 10505 5049 10517 5083
rect 10551 5080 10563 5083
rect 11146 5080 11152 5092
rect 10551 5052 11152 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11425 5083 11483 5089
rect 11425 5049 11437 5083
rect 11471 5080 11483 5083
rect 12437 5083 12495 5089
rect 12437 5080 12449 5083
rect 11471 5052 12449 5080
rect 11471 5049 11483 5052
rect 11425 5043 11483 5049
rect 12437 5049 12449 5052
rect 12483 5049 12495 5083
rect 12437 5043 12495 5049
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 2774 5012 2780 5024
rect 2547 4984 2780 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 2774 4972 2780 4984
rect 2832 5012 2838 5024
rect 3234 5012 3240 5024
rect 2832 4984 3240 5012
rect 2832 4972 2838 4984
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 5040 4984 5089 5012
rect 5040 4972 5046 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5077 4975 5135 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5592 4984 5733 5012
rect 5592 4972 5598 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 6086 5012 6092 5024
rect 6047 4984 6092 5012
rect 5721 4975 5779 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6270 5012 6276 5024
rect 6227 4984 6276 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6270 4972 6276 4984
rect 6328 5012 6334 5024
rect 6730 5012 6736 5024
rect 6328 4984 6736 5012
rect 6328 4972 6334 4984
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7006 5012 7012 5024
rect 6871 4984 7012 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7190 5012 7196 5024
rect 7151 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8202 5012 8208 5024
rect 7524 4984 8208 5012
rect 7524 4972 7530 4984
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8846 5012 8852 5024
rect 8343 4984 8852 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9674 5012 9680 5024
rect 8987 4984 9680 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 10744 4984 11069 5012
rect 10744 4972 10750 4984
rect 11057 4981 11069 4984
rect 11103 4981 11115 5015
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 11057 4975 11115 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 12066 5012 12072 5024
rect 11664 4984 12072 5012
rect 11664 4972 11670 4984
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12544 5012 12572 5120
rect 13357 5083 13415 5089
rect 13357 5049 13369 5083
rect 13403 5080 13415 5083
rect 13446 5080 13452 5092
rect 13403 5052 13452 5080
rect 13403 5049 13415 5052
rect 13357 5043 13415 5049
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 12400 4984 12572 5012
rect 12400 4972 12406 4984
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 12676 4984 13277 5012
rect 12676 4972 12682 4984
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 13265 4975 13323 4981
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 14056 4984 14657 5012
rect 14056 4972 14062 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 14752 5012 14780 5120
rect 16016 5117 16028 5151
rect 16062 5148 16074 5151
rect 17310 5148 17316 5160
rect 16062 5120 17316 5148
rect 16062 5117 16074 5120
rect 16016 5111 16074 5117
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 17405 5151 17463 5157
rect 17405 5117 17417 5151
rect 17451 5148 17463 5151
rect 19518 5148 19524 5160
rect 17451 5120 19524 5148
rect 17451 5117 17463 5120
rect 17405 5111 17463 5117
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 18785 5083 18843 5089
rect 18785 5049 18797 5083
rect 18831 5080 18843 5083
rect 19150 5080 19156 5092
rect 18831 5052 19156 5080
rect 18831 5049 18843 5052
rect 18785 5043 18843 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 19794 5040 19800 5092
rect 19852 5089 19858 5092
rect 19852 5083 19916 5089
rect 19852 5049 19870 5083
rect 19904 5049 19916 5083
rect 19852 5043 19916 5049
rect 19852 5040 19858 5043
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 14752 4984 17141 5012
rect 14645 4975 14703 4981
rect 17129 4981 17141 4984
rect 17175 4981 17187 5015
rect 17129 4975 17187 4981
rect 17589 5015 17647 5021
rect 17589 4981 17601 5015
rect 17635 5012 17647 5015
rect 18690 5012 18696 5024
rect 17635 4984 18696 5012
rect 17635 4981 17647 4984
rect 17589 4975 17647 4981
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 18874 5012 18880 5024
rect 18835 4984 18880 5012
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 20622 5012 20628 5024
rect 20496 4984 20628 5012
rect 20496 4972 20502 4984
rect 20622 4972 20628 4984
rect 20680 5012 20686 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20680 4984 21005 5012
rect 20680 4972 20686 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3602 4808 3608 4820
rect 3559 4780 3608 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 9674 4808 9680 4820
rect 4120 4780 8984 4808
rect 9635 4780 9680 4808
rect 4120 4768 4126 4780
rect 4608 4743 4666 4749
rect 4608 4709 4620 4743
rect 4654 4740 4666 4743
rect 5442 4740 5448 4752
rect 4654 4712 5448 4740
rect 4654 4709 4666 4712
rect 4608 4703 4666 4709
rect 5442 4700 5448 4712
rect 5500 4740 5506 4752
rect 5500 4712 6224 4740
rect 5500 4700 5506 4712
rect 1762 4632 1768 4684
rect 1820 4672 1826 4684
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 1820 4644 2145 4672
rect 1820 4632 1826 4644
rect 2133 4641 2145 4644
rect 2179 4641 2191 4675
rect 2133 4635 2191 4641
rect 2400 4675 2458 4681
rect 2400 4641 2412 4675
rect 2446 4672 2458 4675
rect 3142 4672 3148 4684
rect 2446 4644 3148 4672
rect 2446 4641 2458 4644
rect 2400 4635 2458 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3510 4564 3516 4616
rect 3568 4604 3574 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 3568 4576 4353 4604
rect 3568 4564 3574 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 6196 4604 6224 4712
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6457 4743 6515 4749
rect 6457 4740 6469 4743
rect 6328 4712 6469 4740
rect 6328 4700 6334 4712
rect 6457 4709 6469 4712
rect 6503 4740 6515 4743
rect 6638 4740 6644 4752
rect 6503 4712 6644 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7653 4743 7711 4749
rect 7653 4709 7665 4743
rect 7699 4740 7711 4743
rect 7699 4712 8156 4740
rect 7699 4709 7711 4712
rect 7653 4703 7711 4709
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6196 4576 6561 4604
rect 4341 4567 4399 4573
rect 6549 4573 6561 4576
rect 6595 4573 6607 4607
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 6549 4567 6607 4573
rect 7116 4576 7757 4604
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 5408 4508 6316 4536
rect 5408 4496 5414 4508
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5721 4471 5779 4477
rect 5721 4468 5733 4471
rect 5132 4440 5733 4468
rect 5132 4428 5138 4440
rect 5721 4437 5733 4440
rect 5767 4437 5779 4471
rect 5994 4468 6000 4480
rect 5955 4440 6000 4468
rect 5721 4431 5779 4437
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6288 4468 6316 4508
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 6822 4536 6828 4548
rect 6420 4508 6828 4536
rect 6420 4496 6426 4508
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7116 4468 7144 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7282 4536 7288 4548
rect 7243 4508 7288 4536
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 7760 4536 7788 4567
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7892 4576 7937 4604
rect 7892 4564 7898 4576
rect 7926 4536 7932 4548
rect 7760 4508 7932 4536
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8128 4536 8156 4712
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8956 4740 8984 4780
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 9824 4780 11161 4808
rect 9824 4768 9830 4780
rect 11149 4777 11161 4780
rect 11195 4808 11207 4811
rect 11974 4808 11980 4820
rect 11195 4780 11980 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 15010 4808 15016 4820
rect 12943 4780 15016 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 17862 4808 17868 4820
rect 16071 4780 17868 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 19794 4808 19800 4820
rect 18279 4780 18828 4808
rect 19755 4780 19800 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 11057 4743 11115 4749
rect 11057 4740 11069 4743
rect 8352 4712 8892 4740
rect 8956 4712 11069 4740
rect 8352 4700 8358 4712
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 8260 4644 8677 4672
rect 8260 4632 8266 4644
rect 8665 4641 8677 4644
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8864 4613 8892 4712
rect 11057 4709 11069 4712
rect 11103 4709 11115 4743
rect 11057 4703 11115 4709
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 12069 4743 12127 4749
rect 12069 4740 12081 4743
rect 11388 4712 12081 4740
rect 11388 4700 11394 4712
rect 12069 4709 12081 4712
rect 12115 4709 12127 4743
rect 12069 4703 12127 4709
rect 12161 4743 12219 4749
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 12618 4740 12624 4752
rect 12207 4712 12624 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9766 4672 9772 4684
rect 8996 4644 9772 4672
rect 8996 4632 9002 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 12176 4672 12204 4703
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 13538 4749 13544 4752
rect 13532 4740 13544 4749
rect 13499 4712 13544 4740
rect 13532 4703 13544 4712
rect 13538 4700 13544 4703
rect 13596 4700 13602 4752
rect 13722 4700 13728 4752
rect 13780 4700 13786 4752
rect 15930 4740 15936 4752
rect 15304 4712 15936 4740
rect 10468 4644 12204 4672
rect 12713 4675 12771 4681
rect 10468 4632 10474 4644
rect 12713 4641 12725 4675
rect 12759 4672 12771 4675
rect 13740 4672 13768 4700
rect 12759 4644 13768 4672
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 14550 4672 14556 4684
rect 14148 4644 14556 4672
rect 14148 4632 14154 4644
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 15304 4681 15332 4712
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 16807 4712 17908 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4672 15899 4675
rect 16482 4672 16488 4684
rect 15887 4644 16488 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 16850 4672 16856 4684
rect 16632 4644 16856 4672
rect 16632 4632 16638 4644
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17773 4675 17831 4681
rect 17773 4672 17785 4675
rect 17696 4644 17785 4672
rect 8757 4607 8815 4613
rect 8757 4604 8769 4607
rect 8352 4576 8769 4604
rect 8352 4564 8358 4576
rect 8757 4573 8769 4576
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9950 4604 9956 4616
rect 9732 4576 9956 4604
rect 9732 4564 9738 4576
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 11422 4604 11428 4616
rect 11379 4576 11428 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 8662 4536 8668 4548
rect 8128 4508 8668 4536
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10336 4536 10364 4567
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13078 4604 13084 4616
rect 12584 4576 13084 4604
rect 12584 4564 12590 4576
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13262 4604 13268 4616
rect 13223 4576 13268 4604
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17000 4576 17045 4604
rect 17000 4564 17006 4576
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 9548 4508 10364 4536
rect 16393 4539 16451 4545
rect 9548 4496 9554 4508
rect 16393 4505 16405 4539
rect 16439 4536 16451 4539
rect 17420 4536 17448 4564
rect 16439 4508 17448 4536
rect 16439 4505 16451 4508
rect 16393 4499 16451 4505
rect 6288 4440 7144 4468
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 8297 4471 8355 4477
rect 8297 4468 8309 4471
rect 7432 4440 8309 4468
rect 7432 4428 7438 4440
rect 8297 4437 8309 4440
rect 8343 4437 8355 4471
rect 8297 4431 8355 4437
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 9824 4440 10701 4468
rect 9824 4428 9830 4440
rect 10689 4437 10701 4440
rect 10735 4437 10747 4471
rect 10689 4431 10747 4437
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11701 4471 11759 4477
rect 11701 4468 11713 4471
rect 11020 4440 11713 4468
rect 11020 4428 11026 4440
rect 11701 4437 11713 4440
rect 11747 4437 11759 4471
rect 11701 4431 11759 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14608 4440 14657 4468
rect 14608 4428 14614 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 17310 4468 17316 4480
rect 15519 4440 17316 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 17405 4471 17463 4477
rect 17405 4437 17417 4471
rect 17451 4468 17463 4471
rect 17494 4468 17500 4480
rect 17451 4440 17500 4468
rect 17451 4437 17463 4440
rect 17405 4431 17463 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17696 4468 17724 4644
rect 17773 4641 17785 4644
rect 17819 4641 17831 4675
rect 17880 4672 17908 4712
rect 17954 4700 17960 4752
rect 18012 4740 18018 4752
rect 18662 4743 18720 4749
rect 18662 4740 18674 4743
rect 18012 4712 18674 4740
rect 18012 4700 18018 4712
rect 18662 4709 18674 4712
rect 18708 4709 18720 4743
rect 18800 4740 18828 4780
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 20438 4740 20444 4752
rect 18800 4712 20444 4740
rect 18662 4703 18720 4709
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 18966 4672 18972 4684
rect 17880 4644 18972 4672
rect 17773 4635 17831 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 20257 4675 20315 4681
rect 20257 4641 20269 4675
rect 20303 4672 20315 4675
rect 21634 4672 21640 4684
rect 20303 4644 21640 4672
rect 20303 4641 20315 4644
rect 20257 4635 20315 4641
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18095 4576 18245 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 18233 4567 18291 4573
rect 17770 4496 17776 4548
rect 17828 4536 17834 4548
rect 17880 4536 17908 4567
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 17828 4508 17908 4536
rect 17828 4496 17834 4508
rect 19150 4468 19156 4480
rect 17696 4440 19156 4468
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 20441 4471 20499 4477
rect 20441 4437 20453 4471
rect 20487 4468 20499 4471
rect 22094 4468 22100 4480
rect 20487 4440 22100 4468
rect 20487 4437 20499 4440
rect 20441 4431 20499 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3142 4264 3148 4276
rect 3103 4236 3148 4264
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 4571 4236 5457 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7282 4264 7288 4276
rect 6972 4236 7288 4264
rect 6972 4224 6978 4236
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8941 4267 8999 4273
rect 7576 4236 8616 4264
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 3160 4128 3188 4224
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 6270 4196 6276 4208
rect 4120 4168 6276 4196
rect 4120 4156 4126 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3160 4100 3985 4128
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 3973 4091 4031 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 5684 4100 6101 4128
rect 5684 4088 5690 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 7576 4128 7604 4236
rect 6788 4100 7604 4128
rect 8588 4128 8616 4236
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 9490 4264 9496 4276
rect 8987 4236 9496 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 10060 4236 11376 4264
rect 10060 4208 10088 4236
rect 10042 4196 10048 4208
rect 9600 4168 10048 4196
rect 9600 4128 9628 4168
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 9766 4128 9772 4140
rect 8588 4100 9628 4128
rect 9727 4100 9772 4128
rect 6788 4088 6794 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9950 4128 9956 4140
rect 9911 4100 9956 4128
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 11348 4128 11376 4236
rect 16482 4224 16488 4276
rect 16540 4264 16546 4276
rect 18506 4264 18512 4276
rect 16540 4236 18512 4264
rect 16540 4224 16546 4236
rect 18506 4224 18512 4236
rect 18564 4264 18570 4276
rect 19058 4264 19064 4276
rect 18564 4236 19064 4264
rect 18564 4224 18570 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 18046 4196 18052 4208
rect 15712 4168 18052 4196
rect 15712 4156 15718 4168
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 11882 4128 11888 4140
rect 11348 4100 11888 4128
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13170 4088 13176 4140
rect 13228 4088 13234 4140
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13320 4100 13829 4128
rect 13320 4088 13326 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16942 4128 16948 4140
rect 16531 4100 16948 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16942 4088 16948 4100
rect 17000 4128 17006 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17000 4100 17509 4128
rect 17000 4088 17006 4100
rect 17497 4097 17509 4100
rect 17543 4128 17555 4131
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 17543 4100 18797 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 18785 4097 18797 4100
rect 18831 4128 18843 4131
rect 19058 4128 19064 4140
rect 18831 4100 19064 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19794 4128 19800 4140
rect 19755 4100 19800 4128
rect 19794 4088 19800 4100
rect 19852 4088 19858 4140
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20496 4100 20821 4128
rect 20496 4088 20502 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 5445 4063 5503 4069
rect 3927 4032 4752 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 2032 3995 2090 4001
rect 2032 3961 2044 3995
rect 2078 3992 2090 3995
rect 3326 3992 3332 4004
rect 2078 3964 3332 3992
rect 2078 3961 2090 3964
rect 2032 3955 2090 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3694 3992 3700 4004
rect 3436 3964 3700 3992
rect 3436 3933 3464 3964
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 4724 3992 4752 4032
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5491 4032 6009 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5997 4029 6009 4032
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 5902 3992 5908 4004
rect 4724 3964 5580 3992
rect 5863 3964 5908 3992
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3893 3479 3927
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3421 3887 3479 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4890 3924 4896 3936
rect 4851 3896 4896 3924
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5442 3924 5448 3936
rect 5031 3896 5448 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5552 3933 5580 3964
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7024 3992 7052 4023
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7340 4032 7573 4060
rect 7340 4020 7346 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 10042 4060 10048 4072
rect 7561 4023 7619 4029
rect 7760 4032 10048 4060
rect 7760 3992 7788 4032
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10410 4060 10416 4072
rect 10367 4032 10416 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 12618 4060 12624 4072
rect 10520 4032 12624 4060
rect 7024 3964 7788 3992
rect 7828 3995 7886 4001
rect 7828 3961 7840 3995
rect 7874 3992 7886 3995
rect 8754 3992 8760 4004
rect 7874 3964 8760 3992
rect 7874 3961 7886 3964
rect 7828 3955 7886 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 10520 3992 10548 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12768 4032 12817 4060
rect 12768 4020 12774 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 13188 4060 13216 4088
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 12805 4023 12863 4029
rect 12912 4032 13216 4060
rect 13740 4032 16221 4060
rect 9140 3964 10548 3992
rect 10588 3995 10646 4001
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 9140 3924 9168 3964
rect 10588 3961 10600 3995
rect 10634 3992 10646 3995
rect 11606 3992 11612 4004
rect 10634 3964 11612 3992
rect 10634 3961 10646 3964
rect 10588 3955 10646 3961
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 12912 4001 12940 4032
rect 12897 3995 12955 4001
rect 12897 3961 12909 3995
rect 12943 3961 12955 3995
rect 12897 3955 12955 3961
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 13740 3992 13768 4032
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 17218 4060 17224 4072
rect 17179 4032 17224 4060
rect 16209 4023 16267 4029
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 18472 4032 19564 4060
rect 18472 4020 18478 4032
rect 14090 4001 14096 4004
rect 14084 3992 14096 4001
rect 13228 3964 13768 3992
rect 14051 3964 14096 3992
rect 13228 3952 13234 3964
rect 14084 3955 14096 3964
rect 14090 3952 14096 3955
rect 14148 3952 14154 4004
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 14240 3964 16313 3992
rect 14240 3952 14246 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 17313 3995 17371 4001
rect 17313 3992 17325 3995
rect 16448 3964 17325 3992
rect 16448 3952 16454 3964
rect 17313 3961 17325 3964
rect 17359 3961 17371 3995
rect 19426 3992 19432 4004
rect 17313 3955 17371 3961
rect 19168 3964 19432 3992
rect 9306 3924 9312 3936
rect 7239 3896 9168 3924
rect 9267 3896 9312 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 10686 3924 10692 3936
rect 9723 3896 10692 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 10928 3896 11713 3924
rect 10928 3884 10934 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 11848 3896 12449 3924
rect 11848 3884 11854 3896
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 15160 3896 15209 3924
rect 15160 3884 15166 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 15841 3927 15899 3933
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 16666 3924 16672 3936
rect 15887 3896 16672 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 17460 3896 18153 3924
rect 17460 3884 17466 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18506 3924 18512 3936
rect 18467 3896 18512 3924
rect 18141 3887 18199 3893
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 18598 3884 18604 3936
rect 18656 3924 18662 3936
rect 19168 3933 19196 3964
rect 19426 3952 19432 3964
rect 19484 3952 19490 4004
rect 19536 3992 19564 4032
rect 19536 3964 20392 3992
rect 19153 3927 19211 3933
rect 18656 3896 18701 3924
rect 18656 3884 18662 3896
rect 19153 3893 19165 3927
rect 19199 3893 19211 3927
rect 19153 3887 19211 3893
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19521 3927 19579 3933
rect 19521 3924 19533 3927
rect 19300 3896 19533 3924
rect 19300 3884 19306 3896
rect 19521 3893 19533 3896
rect 19567 3893 19579 3927
rect 19521 3887 19579 3893
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 19668 3896 19713 3924
rect 19668 3884 19674 3896
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 20220 3896 20269 3924
rect 20220 3884 20226 3896
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20364 3924 20392 3964
rect 20530 3952 20536 4004
rect 20588 3992 20594 4004
rect 20717 3995 20775 4001
rect 20717 3992 20729 3995
rect 20588 3964 20729 3992
rect 20588 3952 20594 3964
rect 20717 3961 20729 3964
rect 20763 3961 20775 3995
rect 20717 3955 20775 3961
rect 20622 3924 20628 3936
rect 20364 3896 20628 3924
rect 20257 3887 20315 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3844 3692 4077 3720
rect 3844 3680 3850 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 5994 3720 6000 3732
rect 4948 3692 6000 3720
rect 4948 3680 4954 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7466 3720 7472 3732
rect 7147 3692 7472 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 8754 3720 8760 3732
rect 8715 3692 8760 3720
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 10686 3720 10692 3732
rect 9364 3692 10692 3720
rect 9364 3680 9370 3692
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 10919 3692 11529 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 11882 3720 11888 3732
rect 11843 3692 11888 3720
rect 11517 3683 11575 3689
rect 11882 3680 11888 3692
rect 11940 3720 11946 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 11940 3692 12357 3720
rect 11940 3680 11946 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3689 12587 3723
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12529 3683 12587 3689
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 6730 3652 6736 3664
rect 2004 3624 6736 3652
rect 2004 3612 2010 3624
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 10962 3652 10968 3664
rect 6972 3624 9720 3652
rect 10923 3624 10968 3652
rect 6972 3612 6978 3624
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4212 3556 4445 3584
rect 4212 3544 4218 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 5166 3584 5172 3596
rect 4571 3556 5172 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5988 3587 6046 3593
rect 5988 3553 6000 3587
rect 6034 3584 6046 3587
rect 6362 3584 6368 3596
rect 6034 3556 6368 3584
rect 6034 3553 6046 3556
rect 5988 3547 6046 3553
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7633 3587 7691 3593
rect 7633 3584 7645 3587
rect 7524 3556 7645 3584
rect 7524 3544 7530 3556
rect 7633 3553 7645 3556
rect 7679 3553 7691 3587
rect 7633 3547 7691 3553
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3584 9091 3587
rect 9122 3584 9128 3596
rect 9079 3556 9128 3584
rect 9079 3553 9091 3556
rect 9033 3547 9091 3553
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9692 3593 9720 3624
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 12544 3652 12572 3683
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13817 3723 13875 3729
rect 13817 3689 13829 3723
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 14599 3692 15301 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 15289 3683 15347 3689
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 16574 3720 16580 3732
rect 15795 3692 16580 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 11204 3624 12572 3652
rect 13832 3652 13860 3683
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17773 3723 17831 3729
rect 17773 3689 17785 3723
rect 17819 3720 17831 3723
rect 17954 3720 17960 3732
rect 17819 3692 17960 3720
rect 17819 3689 17831 3692
rect 17773 3683 17831 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 18874 3680 18880 3732
rect 18932 3720 18938 3732
rect 18969 3723 19027 3729
rect 18969 3720 18981 3723
rect 18932 3692 18981 3720
rect 18932 3680 18938 3692
rect 18969 3689 18981 3692
rect 19015 3689 19027 3723
rect 18969 3683 19027 3689
rect 19797 3723 19855 3729
rect 19797 3689 19809 3723
rect 19843 3720 19855 3723
rect 20070 3720 20076 3732
rect 19843 3692 20076 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 17126 3652 17132 3664
rect 13832 3624 17132 3652
rect 11204 3612 11210 3624
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 18984 3652 19012 3683
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20165 3655 20223 3661
rect 20165 3652 20177 3655
rect 18984 3624 20177 3652
rect 20165 3621 20177 3624
rect 20211 3621 20223 3655
rect 20165 3615 20223 3621
rect 20257 3655 20315 3661
rect 20257 3621 20269 3655
rect 20303 3652 20315 3655
rect 20806 3652 20812 3664
rect 20303 3624 20812 3652
rect 20303 3621 20315 3624
rect 20257 3615 20315 3621
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 10192 3556 11989 3584
rect 10192 3544 10198 3556
rect 11977 3553 11989 3556
rect 12023 3584 12035 3587
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12023 3556 12909 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 12897 3553 12909 3556
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3584 13691 3587
rect 15470 3584 15476 3596
rect 13679 3556 15476 3584
rect 13679 3553 13691 3556
rect 13633 3547 13691 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16298 3584 16304 3596
rect 15804 3556 16304 3584
rect 15804 3544 15810 3556
rect 16298 3544 16304 3556
rect 16356 3584 16362 3596
rect 16393 3587 16451 3593
rect 16393 3584 16405 3587
rect 16356 3556 16405 3584
rect 16356 3544 16362 3556
rect 16393 3553 16405 3556
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 16660 3587 16718 3593
rect 16660 3553 16672 3587
rect 16706 3584 16718 3587
rect 16942 3584 16948 3596
rect 16706 3556 16948 3584
rect 16706 3553 16718 3556
rect 16660 3547 16718 3553
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18782 3584 18788 3596
rect 18095 3556 18788 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 18966 3544 18972 3596
rect 19024 3584 19030 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 19024 3556 20913 3584
rect 19024 3544 19030 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 20901 3547 20959 3553
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3384 3488 4629 3516
rect 3384 3476 3390 3488
rect 4617 3485 4629 3488
rect 4663 3516 4675 3519
rect 4890 3516 4896 3528
rect 4663 3488 4896 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5626 3516 5632 3528
rect 5307 3488 5632 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 4908 3448 4936 3476
rect 5534 3448 5540 3460
rect 4908 3420 5540 3448
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 3510 3380 3516 3392
rect 1820 3352 3516 3380
rect 1820 3340 1826 3352
rect 3510 3340 3516 3352
rect 3568 3380 3574 3392
rect 5736 3380 5764 3479
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 7340 3488 7389 3516
rect 7340 3476 7346 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 7377 3479 7435 3485
rect 8404 3488 9873 3516
rect 3568 3352 5764 3380
rect 3568 3340 3574 3352
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 8404 3380 8432 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10870 3516 10876 3528
rect 10008 3488 10876 3516
rect 10008 3476 10014 3488
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10928 3488 11069 3516
rect 10928 3476 10934 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11664 3488 12081 3516
rect 11664 3476 11670 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14056 3488 14657 3516
rect 14056 3476 14062 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3516 14887 3519
rect 15102 3516 15108 3528
rect 14875 3488 15108 3516
rect 14875 3485 14887 3488
rect 14829 3479 14887 3485
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 9217 3451 9275 3457
rect 9217 3417 9229 3451
rect 9263 3448 9275 3451
rect 14366 3448 14372 3460
rect 9263 3420 14372 3448
rect 9263 3417 9275 3420
rect 9217 3411 9275 3417
rect 14366 3408 14372 3420
rect 14424 3408 14430 3460
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 15856 3448 15884 3479
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 18414 3516 18420 3528
rect 17736 3488 18420 3516
rect 17736 3476 17742 3488
rect 18414 3476 18420 3488
rect 18472 3516 18478 3528
rect 19061 3519 19119 3525
rect 19061 3516 19073 3519
rect 18472 3488 19073 3516
rect 18472 3476 18478 3488
rect 19061 3485 19073 3488
rect 19107 3485 19119 3519
rect 19061 3479 19119 3485
rect 19153 3519 19211 3525
rect 19153 3485 19165 3519
rect 19199 3516 19211 3519
rect 19334 3516 19340 3528
rect 19199 3488 19340 3516
rect 19199 3485 19211 3488
rect 19153 3479 19211 3485
rect 14792 3420 15884 3448
rect 14792 3408 14798 3420
rect 18782 3408 18788 3460
rect 18840 3448 18846 3460
rect 19168 3448 19196 3479
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 18840 3420 19196 3448
rect 18840 3408 18846 3420
rect 6512 3352 8432 3380
rect 6512 3340 6518 3352
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 10410 3380 10416 3392
rect 8996 3352 10416 3380
rect 8996 3340 9002 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10505 3383 10563 3389
rect 10505 3349 10517 3383
rect 10551 3380 10563 3383
rect 11146 3380 11152 3392
rect 10551 3352 11152 3380
rect 10551 3349 10563 3352
rect 10505 3343 10563 3349
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 13354 3380 13360 3392
rect 12391 3352 13360 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14185 3383 14243 3389
rect 14185 3349 14197 3383
rect 14231 3380 14243 3383
rect 16114 3380 16120 3392
rect 14231 3352 16120 3380
rect 14231 3349 14243 3352
rect 14185 3343 14243 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 19426 3380 19432 3392
rect 18279 3352 19432 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 4890 3176 4896 3188
rect 4851 3148 4896 3176
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 6411 3148 6653 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6641 3145 6653 3148
rect 6687 3145 6699 3179
rect 6914 3176 6920 3188
rect 6875 3148 6920 3176
rect 6641 3139 6699 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8202 3176 8208 3188
rect 7975 3148 8208 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 8956 3148 10333 3176
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 7282 3108 7288 3120
rect 4856 3080 7288 3108
rect 4856 3068 4862 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 7374 3068 7380 3120
rect 7432 3068 7438 3120
rect 8754 3108 8760 3120
rect 7576 3080 8760 3108
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 5074 3040 5080 3052
rect 4987 3012 5080 3040
rect 5000 2972 5028 3012
rect 5074 3000 5080 3012
rect 5132 3040 5138 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5132 3012 5733 3040
rect 5132 3000 5138 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 4632 2944 5028 2972
rect 4632 2916 4660 2944
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5442 2972 5448 2984
rect 5316 2944 5448 2972
rect 5316 2932 5322 2944
rect 5442 2932 5448 2944
rect 5500 2972 5506 2984
rect 5629 2975 5687 2981
rect 5629 2972 5641 2975
rect 5500 2944 5641 2972
rect 5500 2932 5506 2944
rect 5629 2941 5641 2944
rect 5675 2941 5687 2975
rect 5629 2935 5687 2941
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6454 2972 6460 2984
rect 6227 2944 6460 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7392 2981 7420 3068
rect 7576 3049 7604 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8846 3040 8852 3052
rect 8619 3012 8852 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8846 3000 8852 3012
rect 8904 3040 8910 3052
rect 8956 3040 8984 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 10321 3139 10379 3145
rect 10428 3148 13001 3176
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 10428 3108 10456 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 12989 3139 13047 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 16298 3136 16304 3188
rect 16356 3176 16362 3188
rect 16945 3179 17003 3185
rect 16356 3148 16436 3176
rect 16356 3136 16362 3148
rect 10100 3080 10456 3108
rect 10100 3068 10106 3080
rect 12434 3068 12440 3120
rect 12492 3108 12498 3120
rect 16408 3108 16436 3148
rect 16945 3145 16957 3179
rect 16991 3176 17003 3179
rect 19610 3176 19616 3188
rect 16991 3148 19616 3176
rect 16991 3145 17003 3148
rect 16945 3139 17003 3145
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 12492 3080 16344 3108
rect 16408 3080 18092 3108
rect 12492 3068 12498 3080
rect 8904 3012 8984 3040
rect 8904 3000 8910 3012
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10468 3012 10609 3040
rect 10468 3000 10474 3012
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 11790 3040 11796 3052
rect 10597 3003 10655 3009
rect 11624 3012 11796 3040
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7064 2944 7297 2972
rect 7064 2932 7070 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7800 2944 8309 2972
rect 7800 2932 7806 2944
rect 8297 2941 8309 2944
rect 8343 2972 8355 2975
rect 8386 2972 8392 2984
rect 8343 2944 8392 2972
rect 8343 2941 8355 2944
rect 8297 2935 8355 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8536 2944 8883 2972
rect 8536 2932 8542 2944
rect 3780 2907 3838 2913
rect 3780 2873 3792 2907
rect 3826 2904 3838 2907
rect 4614 2904 4620 2916
rect 3826 2876 4620 2904
rect 3826 2873 3838 2876
rect 3780 2867 3838 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 5718 2904 5724 2916
rect 5132 2876 5724 2904
rect 5132 2864 5138 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 8754 2904 8760 2916
rect 6687 2876 8760 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8855 2904 8883 2944
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 10134 2972 10140 2984
rect 8996 2944 9041 2972
rect 9131 2944 10140 2972
rect 8996 2932 9002 2944
rect 9131 2904 9159 2944
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10870 2981 10876 2984
rect 10864 2972 10876 2981
rect 10831 2944 10876 2972
rect 10864 2935 10876 2944
rect 10870 2932 10876 2935
rect 10928 2932 10934 2984
rect 11624 2972 11652 3012
rect 11790 3000 11796 3012
rect 11848 3040 11854 3052
rect 14645 3043 14703 3049
rect 11848 3012 14596 3040
rect 11848 3000 11854 3012
rect 10980 2944 11652 2972
rect 10980 2916 11008 2944
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12308 2944 12449 2972
rect 12308 2932 12314 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 12437 2935 12495 2941
rect 12544 2944 13185 2972
rect 8855 2876 9159 2904
rect 9208 2907 9266 2913
rect 9208 2873 9220 2907
rect 9254 2904 9266 2907
rect 9254 2876 10916 2904
rect 9254 2873 9266 2876
rect 9208 2867 9266 2873
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 4430 2836 4436 2848
rect 3099 2808 4436 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 5534 2836 5540 2848
rect 5495 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 8386 2836 8392 2848
rect 8347 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2836 8450 2848
rect 9674 2836 9680 2848
rect 8444 2808 9680 2836
rect 8444 2796 8450 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 10888 2836 10916 2876
rect 10962 2864 10968 2916
rect 11020 2864 11026 2916
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 12544 2904 12572 2944
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 14458 2972 14464 2984
rect 14419 2944 14464 2972
rect 13173 2935 13231 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14568 2972 14596 3012
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 16316 3049 16344 3080
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15528 3012 15577 3040
rect 15528 3000 15534 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 16301 3003 16359 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 17954 3040 17960 3052
rect 17635 3012 17960 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18064 3049 18092 3080
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 19429 3111 19487 3117
rect 19429 3108 19441 3111
rect 19116 3080 19441 3108
rect 19116 3068 19122 3080
rect 19429 3077 19441 3080
rect 19475 3077 19487 3111
rect 19429 3071 19487 3077
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 20438 3040 20444 3052
rect 20399 3012 20444 3040
rect 18049 3003 18107 3009
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 15378 2972 15384 2984
rect 14568 2944 14688 2972
rect 15339 2944 15384 2972
rect 11112 2876 12572 2904
rect 12713 2907 12771 2913
rect 11112 2864 11118 2876
rect 12713 2873 12725 2907
rect 12759 2904 12771 2907
rect 12802 2904 12808 2916
rect 12759 2876 12808 2904
rect 12759 2873 12771 2876
rect 12713 2867 12771 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 12989 2907 13047 2913
rect 12989 2873 13001 2907
rect 13035 2904 13047 2907
rect 13449 2907 13507 2913
rect 13449 2904 13461 2907
rect 13035 2876 13461 2904
rect 13035 2873 13047 2876
rect 12989 2867 13047 2873
rect 13449 2873 13461 2876
rect 13495 2873 13507 2907
rect 13449 2867 13507 2873
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 14660 2904 14688 2944
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 16264 2944 16528 2972
rect 16264 2932 16270 2944
rect 16390 2904 16396 2916
rect 13780 2876 14596 2904
rect 14660 2876 16396 2904
rect 13780 2864 13786 2876
rect 11422 2836 11428 2848
rect 10888 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2836 11486 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11480 2808 11989 2836
rect 11480 2796 11486 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 11977 2799 12035 2805
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 13170 2836 13176 2848
rect 12124 2808 13176 2836
rect 12124 2796 12130 2808
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 13412 2808 14381 2836
rect 13412 2796 13418 2808
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 14568 2836 14596 2876
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 16500 2904 16528 2944
rect 16666 2932 16672 2984
rect 16724 2972 16730 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 16724 2944 17325 2972
rect 16724 2932 16730 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 18316 2975 18374 2981
rect 18316 2941 18328 2975
rect 18362 2972 18374 2975
rect 18782 2972 18788 2984
rect 18362 2944 18788 2972
rect 18362 2941 18374 2944
rect 18316 2935 18374 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 20257 2975 20315 2981
rect 20257 2941 20269 2975
rect 20303 2972 20315 2975
rect 22554 2972 22560 2984
rect 20303 2944 22560 2972
rect 20303 2941 20315 2944
rect 20257 2935 20315 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 20806 2904 20812 2916
rect 16500 2876 20812 2904
rect 20806 2864 20812 2876
rect 20864 2864 20870 2916
rect 16298 2836 16304 2848
rect 14568 2808 16304 2836
rect 14369 2799 14427 2805
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4154 2632 4160 2644
rect 4111 2604 4160 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7190 2632 7196 2644
rect 6963 2604 7196 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 8294 2632 8300 2644
rect 8251 2604 8300 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9030 2632 9036 2644
rect 8711 2604 9036 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 10873 2635 10931 2641
rect 10873 2601 10885 2635
rect 10919 2632 10931 2635
rect 11054 2632 11060 2644
rect 10919 2604 11060 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11330 2632 11336 2644
rect 11291 2604 11336 2632
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12161 2635 12219 2641
rect 12161 2601 12173 2635
rect 12207 2632 12219 2635
rect 13722 2632 13728 2644
rect 12207 2604 13728 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 15654 2592 15660 2644
rect 15712 2632 15718 2644
rect 16209 2635 16267 2641
rect 16209 2632 16221 2635
rect 15712 2604 16221 2632
rect 15712 2592 15718 2604
rect 16209 2601 16221 2604
rect 16255 2601 16267 2635
rect 16209 2595 16267 2601
rect 16850 2592 16856 2644
rect 16908 2632 16914 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 16908 2604 17693 2632
rect 16908 2592 16914 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 18564 2604 18613 2632
rect 18564 2592 18570 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 18966 2632 18972 2644
rect 18927 2604 18972 2632
rect 18601 2595 18659 2601
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 2958 2564 2964 2576
rect 2832 2536 2964 2564
rect 2832 2524 2838 2536
rect 2958 2524 2964 2536
rect 3016 2564 3022 2576
rect 4525 2567 4583 2573
rect 4525 2564 4537 2567
rect 3016 2536 4537 2564
rect 3016 2524 3022 2536
rect 4525 2533 4537 2536
rect 4571 2533 4583 2567
rect 4525 2527 4583 2533
rect 6086 2524 6092 2576
rect 6144 2564 6150 2576
rect 6181 2567 6239 2573
rect 6181 2564 6193 2567
rect 6144 2536 6193 2564
rect 6144 2524 6150 2536
rect 6181 2533 6193 2536
rect 6227 2533 6239 2567
rect 6181 2527 6239 2533
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 6696 2536 7389 2564
rect 6696 2524 6702 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 11204 2536 11253 2564
rect 11204 2524 11210 2536
rect 11241 2533 11253 2536
rect 11287 2533 11299 2567
rect 11241 2527 11299 2533
rect 12526 2524 12532 2576
rect 12584 2564 12590 2576
rect 13357 2567 13415 2573
rect 12584 2536 13216 2564
rect 12584 2524 12590 2536
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 5684 2468 7297 2496
rect 5684 2456 5690 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 7285 2459 7343 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 9858 2496 9864 2508
rect 9815 2468 9864 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 11698 2496 11704 2508
rect 10091 2468 11704 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 12434 2496 12440 2508
rect 12023 2468 12440 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 13078 2496 13084 2508
rect 13039 2468 13084 2496
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 13188 2496 13216 2536
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 14274 2564 14280 2576
rect 13403 2536 14280 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 15620 2536 15761 2564
rect 15620 2524 15626 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 17586 2564 17592 2576
rect 17547 2536 17592 2564
rect 15749 2527 15807 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 19058 2564 19064 2576
rect 18104 2536 19064 2564
rect 18104 2524 18110 2536
rect 19058 2524 19064 2536
rect 19116 2524 19122 2576
rect 19518 2524 19524 2576
rect 19576 2564 19582 2576
rect 19889 2567 19947 2573
rect 19889 2564 19901 2567
rect 19576 2536 19901 2564
rect 19576 2524 19582 2536
rect 19889 2533 19901 2536
rect 19935 2533 19947 2567
rect 19889 2527 19947 2533
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13188 2468 13829 2496
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 13817 2459 13875 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14139 2468 14841 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15252 2468 15485 2496
rect 15252 2456 15258 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 17494 2496 17500 2508
rect 16715 2468 17500 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 19613 2499 19671 2505
rect 19613 2465 19625 2499
rect 19659 2496 19671 2499
rect 20346 2496 20352 2508
rect 19659 2468 20352 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 20530 2496 20536 2508
rect 20491 2468 20536 2496
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 6420 2400 6469 2428
rect 6420 2388 6426 2400
rect 6457 2397 6469 2400
rect 6503 2428 6515 2431
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 6503 2400 7573 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 7561 2397 7573 2400
rect 7607 2428 7619 2431
rect 8846 2428 8852 2440
rect 7607 2400 8852 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10870 2428 10876 2440
rect 10376 2400 10876 2428
rect 10376 2388 10382 2400
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11422 2428 11428 2440
rect 11383 2400 11428 2428
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 17954 2428 17960 2440
rect 17911 2400 17960 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 19153 2431 19211 2437
rect 19153 2428 19165 2431
rect 18840 2400 19165 2428
rect 18840 2388 18846 2400
rect 19153 2397 19165 2400
rect 19199 2397 19211 2431
rect 19153 2391 19211 2397
rect 5813 2363 5871 2369
rect 5813 2329 5825 2363
rect 5859 2360 5871 2363
rect 7098 2360 7104 2372
rect 5859 2332 7104 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 7098 2320 7104 2332
rect 7156 2320 7162 2372
rect 16853 2363 16911 2369
rect 16853 2329 16865 2363
rect 16899 2360 16911 2363
rect 18966 2360 18972 2372
rect 16899 2332 18972 2360
rect 16899 2329 16911 2332
rect 16853 2323 16911 2329
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 2406 2252 2412 2304
rect 2464 2292 2470 2304
rect 7742 2292 7748 2304
rect 2464 2264 7748 2292
rect 2464 2252 2470 2264
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 15838 2292 15844 2304
rect 15059 2264 15844 2292
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2292 17279 2295
rect 19150 2292 19156 2304
rect 17267 2264 19156 2292
rect 17267 2261 17279 2264
rect 17221 2255 17279 2261
rect 19150 2252 19156 2264
rect 19208 2252 19214 2304
rect 20714 2292 20720 2304
rect 20675 2264 20720 2292
rect 20714 2252 20720 2264
rect 20772 2252 20778 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 18598 2088 18604 2100
rect 17092 2060 18604 2088
rect 17092 2048 17098 2060
rect 18598 2048 18604 2060
rect 18656 2048 18662 2100
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 11974 2020 11980 2032
rect 11388 1992 11980 2020
rect 11388 1980 11394 1992
rect 11974 1980 11980 1992
rect 12032 1980 12038 2032
rect 1486 1844 1492 1896
rect 1544 1884 1550 1896
rect 8386 1884 8392 1896
rect 1544 1856 8392 1884
rect 1544 1844 1550 1856
rect 8386 1844 8392 1856
rect 8444 1844 8450 1896
rect 566 1776 572 1828
rect 624 1816 630 1828
rect 8570 1816 8576 1828
rect 624 1788 8576 1816
rect 624 1776 630 1788
rect 8570 1776 8576 1788
rect 8628 1776 8634 1828
rect 198 1640 204 1692
rect 256 1680 262 1692
rect 5810 1680 5816 1692
rect 256 1652 5816 1680
rect 256 1640 262 1652
rect 5810 1640 5816 1652
rect 5868 1640 5874 1692
rect 1026 1504 1032 1556
rect 1084 1544 1090 1556
rect 8478 1544 8484 1556
rect 1084 1516 8484 1544
rect 1084 1504 1090 1516
rect 8478 1504 8484 1516
rect 8536 1504 8542 1556
rect 3878 1096 3884 1148
rect 3936 1136 3942 1148
rect 5442 1136 5448 1148
rect 3936 1108 5448 1136
rect 3936 1096 3942 1108
rect 5442 1096 5448 1108
rect 5500 1096 5506 1148
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3884 19456 3936 19508
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 4988 19252 5040 19304
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 18420 19252 18472 19304
rect 19708 19252 19760 19304
rect 6092 19184 6144 19236
rect 2780 19116 2832 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 5632 18844 5684 18896
rect 18420 18887 18472 18896
rect 18420 18853 18429 18887
rect 18429 18853 18463 18887
rect 18463 18853 18472 18887
rect 18420 18844 18472 18853
rect 1492 18776 1544 18828
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 19616 18776 19668 18828
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 5724 18164 5776 18216
rect 8208 18164 8260 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1768 17756 1820 17808
rect 20536 17756 20588 17808
rect 6736 17688 6788 17740
rect 20260 17688 20312 17740
rect 7380 17620 7432 17672
rect 1676 17552 1728 17604
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 7104 17076 7156 17128
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1860 16736 1912 16788
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 4896 16600 4948 16652
rect 20628 16600 20680 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 17868 16192 17920 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20812 16192 20864 16244
rect 7472 16056 7524 16108
rect 3148 16031 3200 16040
rect 3148 15997 3157 16031
rect 3157 15997 3191 16031
rect 3191 15997 3200 16031
rect 3148 15988 3200 15997
rect 12808 15988 12860 16040
rect 19340 15988 19392 16040
rect 20168 15988 20220 16040
rect 4712 15920 4764 15972
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2412 15648 2464 15700
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 3148 15580 3200 15632
rect 12808 15623 12860 15632
rect 12808 15589 12817 15623
rect 12817 15589 12851 15623
rect 12851 15589 12860 15623
rect 12808 15580 12860 15589
rect 4252 15512 4304 15564
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 5080 15444 5132 15496
rect 19984 15512 20036 15564
rect 20812 15444 20864 15496
rect 5172 15376 5224 15428
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2780 15104 2832 15156
rect 20076 15104 20128 15156
rect 20352 15104 20404 15156
rect 1952 15079 2004 15088
rect 1952 15045 1961 15079
rect 1961 15045 1995 15079
rect 1995 15045 2004 15079
rect 1952 15036 2004 15045
rect 19616 15079 19668 15088
rect 19616 15045 19625 15079
rect 19625 15045 19659 15079
rect 19659 15045 19668 15079
rect 19616 15036 19668 15045
rect 2412 14968 2464 15020
rect 16396 14968 16448 15020
rect 17500 14968 17552 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 5908 14900 5960 14952
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 3792 14832 3844 14884
rect 12716 14832 12768 14884
rect 4160 14764 4212 14816
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16580 14807 16632 14816
rect 16580 14773 16589 14807
rect 16589 14773 16623 14807
rect 16623 14773 16632 14807
rect 16580 14764 16632 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 3424 14560 3476 14612
rect 11704 14560 11756 14612
rect 17132 14560 17184 14612
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 1768 14492 1820 14544
rect 7748 14492 7800 14544
rect 1860 14424 1912 14476
rect 2872 14424 2924 14476
rect 5356 14424 5408 14476
rect 9864 14424 9916 14476
rect 3332 14399 3384 14408
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 4160 14356 4212 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 10508 14399 10560 14408
rect 7564 14288 7616 14340
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 11152 14356 11204 14408
rect 12440 14424 12492 14476
rect 8208 14288 8260 14340
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 7196 14220 7248 14229
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 15292 14424 15344 14476
rect 16396 14424 16448 14476
rect 18604 14467 18656 14476
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 18696 14424 18748 14476
rect 19432 14492 19484 14544
rect 14740 14356 14792 14408
rect 15016 14356 15068 14408
rect 15568 14356 15620 14408
rect 13544 14220 13596 14272
rect 15200 14220 15252 14272
rect 16120 14220 16172 14272
rect 20536 14356 20588 14408
rect 17040 14288 17092 14340
rect 20628 14288 20680 14340
rect 17132 14263 17184 14272
rect 17132 14229 17141 14263
rect 17141 14229 17175 14263
rect 17175 14229 17184 14263
rect 17132 14220 17184 14229
rect 18880 14220 18932 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2412 14016 2464 14068
rect 2136 13880 2188 13932
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 11152 14016 11204 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 5264 13948 5316 14000
rect 7288 13948 7340 14000
rect 9772 13991 9824 14000
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 3240 13812 3292 13864
rect 4160 13812 4212 13864
rect 4804 13812 4856 13864
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 7564 13880 7616 13932
rect 8668 13855 8720 13864
rect 8668 13821 8702 13855
rect 8702 13821 8720 13855
rect 8668 13812 8720 13821
rect 3148 13744 3200 13796
rect 5080 13744 5132 13796
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8484 13744 8536 13796
rect 10140 13812 10192 13864
rect 10968 13744 11020 13796
rect 12440 13812 12492 13864
rect 13084 13812 13136 13864
rect 14464 13812 14516 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 11244 13744 11296 13796
rect 19248 14016 19300 14068
rect 17132 13880 17184 13932
rect 16212 13812 16264 13864
rect 19340 13948 19392 14000
rect 19708 13948 19760 14000
rect 18604 13880 18656 13932
rect 20812 13923 20864 13932
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 18788 13855 18840 13864
rect 18788 13821 18797 13855
rect 18797 13821 18831 13855
rect 18831 13821 18840 13855
rect 18788 13812 18840 13821
rect 19524 13812 19576 13864
rect 16856 13744 16908 13796
rect 17224 13744 17276 13796
rect 18604 13744 18656 13796
rect 19708 13744 19760 13796
rect 15752 13676 15804 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 16396 13676 16448 13685
rect 17408 13676 17460 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2872 13472 2924 13524
rect 3332 13472 3384 13524
rect 3516 13472 3568 13524
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 6000 13472 6052 13524
rect 6828 13472 6880 13524
rect 7196 13404 7248 13456
rect 11704 13472 11756 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 16580 13472 16632 13524
rect 19800 13472 19852 13524
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 3884 13336 3936 13388
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 7288 13379 7340 13388
rect 7288 13345 7297 13379
rect 7297 13345 7331 13379
rect 7331 13345 7340 13379
rect 7288 13336 7340 13345
rect 2504 13268 2556 13320
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 3792 13268 3844 13320
rect 4712 13268 4764 13320
rect 3976 13200 4028 13252
rect 5448 13268 5500 13320
rect 9956 13404 10008 13456
rect 10416 13447 10468 13456
rect 10416 13413 10425 13447
rect 10425 13413 10459 13447
rect 10459 13413 10468 13447
rect 10416 13404 10468 13413
rect 7564 13379 7616 13388
rect 7564 13345 7598 13379
rect 7598 13345 7616 13379
rect 7564 13336 7616 13345
rect 7840 13336 7892 13388
rect 10140 13268 10192 13320
rect 11060 13404 11112 13456
rect 11152 13404 11204 13456
rect 15568 13404 15620 13456
rect 17132 13404 17184 13456
rect 13084 13379 13136 13388
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 7196 13200 7248 13252
rect 10692 13268 10744 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 12808 13268 12860 13320
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 16304 13336 16356 13388
rect 18512 13404 18564 13456
rect 14740 13311 14792 13320
rect 10324 13132 10376 13184
rect 10784 13200 10836 13252
rect 12992 13200 13044 13252
rect 12348 13175 12400 13184
rect 12348 13141 12357 13175
rect 12357 13141 12391 13175
rect 12391 13141 12400 13175
rect 12348 13132 12400 13141
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 14464 13200 14516 13252
rect 19984 13336 20036 13388
rect 18512 13268 18564 13320
rect 19800 13268 19852 13320
rect 16672 13132 16724 13184
rect 19892 13132 19944 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 3424 12928 3476 12980
rect 3884 12928 3936 12980
rect 10508 12928 10560 12980
rect 10600 12928 10652 12980
rect 14280 12928 14332 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 18788 12928 18840 12980
rect 4068 12860 4120 12912
rect 4160 12860 4212 12912
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 3700 12724 3752 12776
rect 7012 12724 7064 12776
rect 8668 12860 8720 12912
rect 10784 12860 10836 12912
rect 12164 12860 12216 12912
rect 9680 12792 9732 12844
rect 10048 12792 10100 12844
rect 10140 12792 10192 12844
rect 10508 12792 10560 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 11980 12792 12032 12844
rect 15936 12860 15988 12912
rect 20260 12860 20312 12912
rect 12716 12792 12768 12844
rect 14464 12835 14516 12844
rect 3056 12656 3108 12708
rect 4712 12656 4764 12708
rect 2964 12588 3016 12640
rect 3792 12588 3844 12640
rect 4620 12588 4672 12640
rect 5448 12656 5500 12708
rect 12348 12724 12400 12776
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 16028 12792 16080 12844
rect 16396 12792 16448 12844
rect 16856 12792 16908 12844
rect 17408 12835 17460 12844
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 19984 12792 20036 12844
rect 14740 12724 14792 12776
rect 15568 12724 15620 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 9588 12656 9640 12708
rect 10508 12699 10560 12708
rect 9956 12588 10008 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 10508 12665 10517 12699
rect 10517 12665 10551 12699
rect 10551 12665 10560 12699
rect 10508 12656 10560 12665
rect 11704 12699 11756 12708
rect 11704 12665 11713 12699
rect 11713 12665 11747 12699
rect 11747 12665 11756 12699
rect 11704 12656 11756 12665
rect 12808 12699 12860 12708
rect 12808 12665 12817 12699
rect 12817 12665 12851 12699
rect 12851 12665 12860 12699
rect 12808 12656 12860 12665
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 11612 12588 11664 12640
rect 12072 12588 12124 12640
rect 17500 12656 17552 12708
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 15844 12588 15896 12597
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 16488 12588 16540 12640
rect 17592 12588 17644 12640
rect 18788 12631 18840 12640
rect 18788 12597 18797 12631
rect 18797 12597 18831 12631
rect 18831 12597 18840 12631
rect 18788 12588 18840 12597
rect 20536 12656 20588 12708
rect 20720 12699 20772 12708
rect 20720 12665 20729 12699
rect 20729 12665 20763 12699
rect 20763 12665 20772 12699
rect 20720 12656 20772 12665
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 19800 12588 19852 12597
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2320 12384 2372 12436
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 7564 12384 7616 12436
rect 7748 12384 7800 12436
rect 9312 12384 9364 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 10324 12427 10376 12436
rect 10324 12393 10333 12427
rect 10333 12393 10367 12427
rect 10367 12393 10376 12427
rect 10324 12384 10376 12393
rect 1400 12316 1452 12368
rect 3976 12316 4028 12368
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 3240 12248 3292 12300
rect 3516 12248 3568 12300
rect 4896 12248 4948 12300
rect 5448 12248 5500 12300
rect 6920 12248 6972 12300
rect 8024 12248 8076 12300
rect 10140 12316 10192 12368
rect 12808 12384 12860 12436
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 15844 12384 15896 12436
rect 18512 12384 18564 12436
rect 18972 12384 19024 12436
rect 19340 12384 19392 12436
rect 20536 12384 20588 12436
rect 10600 12316 10652 12368
rect 17500 12316 17552 12368
rect 3148 12180 3200 12232
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 6000 12180 6052 12232
rect 10968 12248 11020 12300
rect 11888 12248 11940 12300
rect 15660 12248 15712 12300
rect 18880 12316 18932 12368
rect 19892 12316 19944 12368
rect 19064 12248 19116 12300
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 8668 12180 8720 12232
rect 3240 12112 3292 12164
rect 1860 12044 1912 12096
rect 7288 12112 7340 12164
rect 7380 12112 7432 12164
rect 7932 12112 7984 12164
rect 8024 12112 8076 12164
rect 9772 12180 9824 12232
rect 12072 12180 12124 12232
rect 12992 12180 13044 12232
rect 8852 12112 8904 12164
rect 10692 12112 10744 12164
rect 12256 12155 12308 12164
rect 12256 12121 12265 12155
rect 12265 12121 12299 12155
rect 12299 12121 12308 12155
rect 12256 12112 12308 12121
rect 7104 12044 7156 12096
rect 7748 12044 7800 12096
rect 11796 12044 11848 12096
rect 12808 12044 12860 12096
rect 16580 12180 16632 12232
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 17960 12180 18012 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 17316 12112 17368 12164
rect 17408 12112 17460 12164
rect 16304 12044 16356 12096
rect 17960 12044 18012 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 5356 11840 5408 11892
rect 6184 11772 6236 11824
rect 7656 11840 7708 11892
rect 10600 11840 10652 11892
rect 10692 11840 10744 11892
rect 11888 11840 11940 11892
rect 8484 11815 8536 11824
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 2412 11636 2464 11688
rect 5264 11704 5316 11756
rect 5816 11704 5868 11756
rect 6552 11704 6604 11756
rect 8024 11747 8076 11756
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 8484 11781 8493 11815
rect 8493 11781 8527 11815
rect 8527 11781 8536 11815
rect 8484 11772 8536 11781
rect 11704 11772 11756 11824
rect 14096 11840 14148 11892
rect 15660 11883 15712 11892
rect 8208 11636 8260 11688
rect 2964 11568 3016 11620
rect 4160 11568 4212 11620
rect 4896 11568 4948 11620
rect 5172 11568 5224 11620
rect 5448 11611 5500 11620
rect 5448 11577 5457 11611
rect 5457 11577 5491 11611
rect 5491 11577 5500 11611
rect 5448 11568 5500 11577
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 2872 11543 2924 11552
rect 2320 11500 2372 11509
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 5816 11500 5868 11552
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 7380 11568 7432 11620
rect 7932 11611 7984 11620
rect 7932 11577 7941 11611
rect 7941 11577 7975 11611
rect 7975 11577 7984 11611
rect 7932 11568 7984 11577
rect 9588 11568 9640 11620
rect 8300 11500 8352 11552
rect 8484 11500 8536 11552
rect 11888 11704 11940 11756
rect 12348 11772 12400 11824
rect 12992 11747 13044 11756
rect 12164 11636 12216 11688
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 15844 11840 15896 11892
rect 19984 11840 20036 11892
rect 20996 11840 21048 11892
rect 18696 11772 18748 11824
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 17316 11704 17368 11756
rect 15292 11636 15344 11688
rect 17960 11636 18012 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 19340 11679 19392 11688
rect 19340 11645 19374 11679
rect 19374 11645 19392 11679
rect 19340 11636 19392 11645
rect 20720 11679 20772 11688
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 14556 11611 14608 11620
rect 14556 11577 14590 11611
rect 14590 11577 14608 11611
rect 14556 11568 14608 11577
rect 10232 11500 10284 11552
rect 10968 11500 11020 11552
rect 12348 11500 12400 11552
rect 13084 11500 13136 11552
rect 17592 11500 17644 11552
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 19340 11500 19392 11552
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 1768 11160 1820 11212
rect 2412 11160 2464 11212
rect 4068 11160 4120 11212
rect 6000 11296 6052 11348
rect 6828 11296 6880 11348
rect 7748 11296 7800 11348
rect 3608 11092 3660 11144
rect 8300 11228 8352 11280
rect 10784 11228 10836 11280
rect 12256 11228 12308 11280
rect 12440 11228 12492 11280
rect 12992 11296 13044 11348
rect 13544 11228 13596 11280
rect 14096 11296 14148 11348
rect 18788 11296 18840 11348
rect 20352 11296 20404 11348
rect 15476 11228 15528 11280
rect 15844 11228 15896 11280
rect 5448 11160 5500 11212
rect 3516 11024 3568 11076
rect 5540 11024 5592 11076
rect 7472 11160 7524 11212
rect 7656 11067 7708 11076
rect 7656 11033 7665 11067
rect 7665 11033 7699 11067
rect 7699 11033 7708 11067
rect 7656 11024 7708 11033
rect 9772 11160 9824 11212
rect 10968 11160 11020 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 15568 11160 15620 11212
rect 10232 11092 10284 11101
rect 14556 11092 14608 11144
rect 16856 11228 16908 11280
rect 16948 11160 17000 11212
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 17776 11160 17828 11212
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 17868 11135 17920 11144
rect 16856 11092 16908 11101
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18880 11092 18932 11144
rect 19064 11092 19116 11144
rect 20352 11135 20404 11144
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 3148 10956 3200 11008
rect 4160 10956 4212 11008
rect 4988 10956 5040 11008
rect 7840 10956 7892 11008
rect 9680 10999 9732 11008
rect 9680 10965 9689 10999
rect 9689 10965 9723 10999
rect 9723 10965 9732 10999
rect 9680 10956 9732 10965
rect 16580 11024 16632 11076
rect 18512 11024 18564 11076
rect 12900 10956 12952 11008
rect 17040 10956 17092 11008
rect 20076 10956 20128 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1676 10752 1728 10804
rect 3148 10752 3200 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 3516 10616 3568 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 3976 10616 4028 10668
rect 6184 10659 6236 10668
rect 3884 10548 3936 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 8484 10752 8536 10804
rect 9772 10752 9824 10804
rect 10140 10752 10192 10804
rect 7840 10684 7892 10736
rect 12164 10752 12216 10804
rect 12348 10684 12400 10736
rect 13820 10684 13872 10736
rect 15292 10727 15344 10736
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 11612 10616 11664 10668
rect 12256 10616 12308 10668
rect 13544 10616 13596 10668
rect 14372 10616 14424 10668
rect 15292 10693 15301 10727
rect 15301 10693 15335 10727
rect 15335 10693 15344 10727
rect 15292 10684 15344 10693
rect 16396 10727 16448 10736
rect 16396 10693 16405 10727
rect 16405 10693 16439 10727
rect 16439 10693 16448 10727
rect 16396 10684 16448 10693
rect 15016 10616 15068 10668
rect 4160 10480 4212 10532
rect 5172 10480 5224 10532
rect 5264 10480 5316 10532
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 12992 10548 13044 10600
rect 16212 10616 16264 10668
rect 16672 10616 16724 10668
rect 19064 10752 19116 10804
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 19432 10548 19484 10600
rect 20444 10548 20496 10600
rect 7748 10480 7800 10532
rect 10968 10480 11020 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 5724 10455 5776 10464
rect 3516 10412 3568 10421
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6920 10412 6972 10464
rect 9312 10412 9364 10464
rect 10324 10412 10376 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 11704 10455 11756 10464
rect 10508 10412 10560 10421
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 11796 10412 11848 10464
rect 12624 10480 12676 10532
rect 12900 10412 12952 10464
rect 12992 10412 13044 10464
rect 14464 10412 14516 10464
rect 17132 10480 17184 10532
rect 15292 10412 15344 10464
rect 16028 10412 16080 10464
rect 17960 10412 18012 10464
rect 20352 10412 20404 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2044 10208 2096 10260
rect 2504 10208 2556 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 5356 10208 5408 10260
rect 2596 10140 2648 10192
rect 3608 10140 3660 10192
rect 5724 10140 5776 10192
rect 1768 10115 1820 10124
rect 1768 10081 1777 10115
rect 1777 10081 1811 10115
rect 1811 10081 1820 10115
rect 1768 10072 1820 10081
rect 2044 10115 2096 10124
rect 2044 10081 2078 10115
rect 2078 10081 2096 10115
rect 2044 10072 2096 10081
rect 5632 10115 5684 10124
rect 5632 10081 5641 10115
rect 5641 10081 5675 10115
rect 5675 10081 5684 10115
rect 5632 10072 5684 10081
rect 7012 10208 7064 10260
rect 7472 10208 7524 10260
rect 7748 10208 7800 10260
rect 8208 10208 8260 10260
rect 9588 10208 9640 10260
rect 11980 10251 12032 10260
rect 7104 10140 7156 10192
rect 7380 10140 7432 10192
rect 5540 10004 5592 10056
rect 6000 10072 6052 10124
rect 6184 10072 6236 10124
rect 7564 10072 7616 10124
rect 8208 10072 8260 10124
rect 9680 10140 9732 10192
rect 10232 10072 10284 10124
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 13820 10208 13872 10260
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 15936 10208 15988 10260
rect 16672 10208 16724 10260
rect 20168 10208 20220 10260
rect 17684 10140 17736 10192
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 13912 10072 13964 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 19432 10140 19484 10192
rect 9128 10047 9180 10056
rect 5448 9936 5500 9988
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 8484 9936 8536 9988
rect 11060 10004 11112 10056
rect 11796 10004 11848 10056
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 12440 10004 12492 10056
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 14556 10047 14608 10056
rect 13176 10004 13228 10013
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 4068 9868 4120 9920
rect 10876 9868 10928 9920
rect 11796 9868 11848 9920
rect 16120 9868 16172 9920
rect 19800 10072 19852 10124
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 20628 9936 20680 9988
rect 18788 9868 18840 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2412 9664 2464 9716
rect 3976 9664 4028 9716
rect 10048 9664 10100 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 10784 9664 10836 9716
rect 3332 9596 3384 9648
rect 4804 9639 4856 9648
rect 4804 9605 4813 9639
rect 4813 9605 4847 9639
rect 4847 9605 4856 9639
rect 4804 9596 4856 9605
rect 6736 9596 6788 9648
rect 7564 9596 7616 9648
rect 1860 9528 1912 9580
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 2688 9528 2740 9580
rect 5080 9528 5132 9580
rect 6920 9528 6972 9580
rect 7748 9528 7800 9580
rect 8484 9528 8536 9580
rect 2872 9460 2924 9512
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 3608 9460 3660 9512
rect 7196 9460 7248 9512
rect 7656 9460 7708 9512
rect 4068 9392 4120 9444
rect 10692 9460 10744 9512
rect 11336 9596 11388 9648
rect 15660 9596 15712 9648
rect 16764 9664 16816 9716
rect 17960 9664 18012 9716
rect 17776 9596 17828 9648
rect 14556 9528 14608 9580
rect 11244 9460 11296 9512
rect 12532 9460 12584 9512
rect 16396 9528 16448 9580
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 18788 9528 18840 9580
rect 19432 9528 19484 9580
rect 15476 9460 15528 9512
rect 17776 9460 17828 9512
rect 18604 9460 18656 9512
rect 20352 9460 20404 9512
rect 9864 9392 9916 9444
rect 10876 9435 10928 9444
rect 10876 9401 10885 9435
rect 10885 9401 10919 9435
rect 10919 9401 10928 9435
rect 10876 9392 10928 9401
rect 13084 9392 13136 9444
rect 2964 9324 3016 9376
rect 3056 9324 3108 9376
rect 6920 9324 6972 9376
rect 8300 9324 8352 9376
rect 8484 9324 8536 9376
rect 14004 9392 14056 9444
rect 13912 9324 13964 9376
rect 17408 9435 17460 9444
rect 17408 9401 17417 9435
rect 17417 9401 17451 9435
rect 17451 9401 17460 9435
rect 17408 9392 17460 9401
rect 20444 9392 20496 9444
rect 16304 9324 16356 9376
rect 18420 9367 18472 9376
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 18604 9324 18656 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2320 9120 2372 9172
rect 5632 9120 5684 9172
rect 7564 9163 7616 9172
rect 7564 9129 7573 9163
rect 7573 9129 7607 9163
rect 7607 9129 7616 9163
rect 7564 9120 7616 9129
rect 4068 9052 4120 9104
rect 9772 9052 9824 9104
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10876 9120 10928 9172
rect 11336 9120 11388 9172
rect 12532 9120 12584 9172
rect 10140 9052 10192 9061
rect 12348 9052 12400 9104
rect 3148 8984 3200 9036
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6736 8984 6788 9036
rect 7196 8984 7248 9036
rect 7656 8984 7708 9036
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 2872 8916 2924 8968
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 8392 8984 8444 9036
rect 9036 8984 9088 9036
rect 9956 8984 10008 9036
rect 10784 8984 10836 9036
rect 8484 8959 8536 8968
rect 5080 8848 5132 8900
rect 6368 8780 6420 8832
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 8668 8916 8720 8968
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 13084 9120 13136 9172
rect 15752 9120 15804 9172
rect 15936 9120 15988 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 12716 9052 12768 9104
rect 12900 9052 12952 9104
rect 13084 8984 13136 9036
rect 15292 9052 15344 9104
rect 16304 9052 16356 9104
rect 18420 9120 18472 9172
rect 19800 9163 19852 9172
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 14648 8959 14700 8968
rect 8116 8848 8168 8900
rect 7288 8780 7340 8832
rect 8300 8780 8352 8832
rect 9496 8780 9548 8832
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 9864 8848 9916 8900
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 17684 8984 17736 9036
rect 19432 8984 19484 9036
rect 19892 8984 19944 9036
rect 15292 8959 15344 8968
rect 14556 8848 14608 8900
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 17960 8916 18012 8968
rect 14832 8848 14884 8900
rect 13820 8780 13872 8832
rect 14372 8780 14424 8832
rect 19616 8848 19668 8900
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2596 8576 2648 8628
rect 3516 8576 3568 8628
rect 4896 8576 4948 8628
rect 7840 8576 7892 8628
rect 8208 8576 8260 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 10692 8576 10744 8628
rect 4436 8508 4488 8560
rect 4988 8508 5040 8560
rect 3608 8440 3660 8492
rect 4528 8440 4580 8492
rect 6920 8508 6972 8560
rect 9588 8508 9640 8560
rect 10324 8508 10376 8560
rect 12256 8576 12308 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 14648 8576 14700 8628
rect 18972 8576 19024 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 12532 8508 12584 8560
rect 14832 8551 14884 8560
rect 14832 8517 14841 8551
rect 14841 8517 14875 8551
rect 14875 8517 14884 8551
rect 14832 8508 14884 8517
rect 19616 8508 19668 8560
rect 19984 8508 20036 8560
rect 7380 8440 7432 8492
rect 7564 8440 7616 8492
rect 9496 8440 9548 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3884 8372 3936 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 6736 8372 6788 8424
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 8576 8372 8628 8424
rect 2596 8304 2648 8356
rect 6460 8304 6512 8356
rect 10232 8372 10284 8424
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 12256 8440 12308 8492
rect 12716 8440 12768 8492
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 16396 8483 16448 8492
rect 16396 8449 16405 8483
rect 16405 8449 16439 8483
rect 16439 8449 16448 8483
rect 16396 8440 16448 8449
rect 9220 8304 9272 8356
rect 9404 8304 9456 8356
rect 11336 8304 11388 8356
rect 11888 8304 11940 8356
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 4896 8236 4948 8288
rect 6276 8279 6328 8288
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 7472 8236 7524 8288
rect 14004 8304 14056 8356
rect 14280 8304 14332 8356
rect 16212 8372 16264 8424
rect 17684 8372 17736 8424
rect 17960 8372 18012 8424
rect 19800 8440 19852 8492
rect 18696 8372 18748 8424
rect 19248 8372 19300 8424
rect 20812 8372 20864 8424
rect 18512 8304 18564 8356
rect 18604 8304 18656 8356
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13268 8236 13320 8288
rect 13636 8236 13688 8288
rect 16120 8236 16172 8288
rect 17224 8279 17276 8288
rect 17224 8245 17233 8279
rect 17233 8245 17267 8279
rect 17267 8245 17276 8279
rect 17224 8236 17276 8245
rect 17316 8279 17368 8288
rect 17316 8245 17325 8279
rect 17325 8245 17359 8279
rect 17359 8245 17368 8279
rect 17316 8236 17368 8245
rect 19984 8236 20036 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2228 8032 2280 8084
rect 3792 8032 3844 8084
rect 4160 8032 4212 8084
rect 4988 8032 5040 8084
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 4804 7964 4856 8016
rect 5172 7964 5224 8016
rect 2688 7896 2740 7948
rect 4528 7896 4580 7948
rect 5632 7939 5684 7948
rect 2228 7828 2280 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 3608 7871 3660 7880
rect 2596 7828 2648 7837
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 4160 7828 4212 7880
rect 4620 7828 4672 7880
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6276 7964 6328 8016
rect 7380 8032 7432 8084
rect 10232 8075 10284 8084
rect 10232 8041 10241 8075
rect 10241 8041 10275 8075
rect 10275 8041 10284 8075
rect 10232 8032 10284 8041
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 11428 8032 11480 8084
rect 12072 8032 12124 8084
rect 12900 8032 12952 8084
rect 13912 8032 13964 8084
rect 14004 8075 14056 8084
rect 14004 8041 14013 8075
rect 14013 8041 14047 8075
rect 14047 8041 14056 8075
rect 14004 8032 14056 8041
rect 9956 7964 10008 8016
rect 10968 7964 11020 8016
rect 12348 7964 12400 8016
rect 16488 8032 16540 8084
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 2872 7760 2924 7812
rect 8484 7896 8536 7948
rect 10048 7896 10100 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 11336 7896 11388 7948
rect 2688 7692 2740 7744
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 6828 7760 6880 7812
rect 7656 7828 7708 7880
rect 9220 7871 9272 7880
rect 7196 7760 7248 7812
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 10232 7828 10284 7880
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 15752 7964 15804 8016
rect 15936 8007 15988 8016
rect 15936 7973 15970 8007
rect 15970 7973 15988 8007
rect 15936 7964 15988 7973
rect 16764 7964 16816 8016
rect 15016 7896 15068 7948
rect 15292 7896 15344 7948
rect 17960 7896 18012 7948
rect 20076 7939 20128 7948
rect 20076 7905 20085 7939
rect 20085 7905 20119 7939
rect 20119 7905 20128 7939
rect 20076 7896 20128 7905
rect 10416 7828 10468 7837
rect 6552 7692 6604 7744
rect 10508 7692 10560 7744
rect 11428 7760 11480 7812
rect 11704 7760 11756 7812
rect 11796 7760 11848 7812
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 19064 7828 19116 7880
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 14924 7760 14976 7812
rect 18696 7760 18748 7812
rect 19892 7760 19944 7812
rect 12348 7692 12400 7744
rect 15016 7692 15068 7744
rect 17040 7735 17092 7744
rect 17040 7701 17049 7735
rect 17049 7701 17083 7735
rect 17083 7701 17092 7735
rect 17040 7692 17092 7701
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 5356 7488 5408 7540
rect 5908 7488 5960 7540
rect 6276 7488 6328 7540
rect 6644 7488 6696 7540
rect 8392 7488 8444 7540
rect 9220 7488 9272 7540
rect 1492 7420 1544 7472
rect 3516 7352 3568 7404
rect 4068 7420 4120 7472
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 5172 7352 5224 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 7656 7284 7708 7336
rect 8208 7284 8260 7336
rect 10140 7488 10192 7540
rect 15108 7531 15160 7540
rect 13084 7420 13136 7472
rect 3884 7259 3936 7268
rect 3884 7225 3893 7259
rect 3893 7225 3927 7259
rect 3927 7225 3936 7259
rect 3884 7216 3936 7225
rect 8668 7284 8720 7336
rect 10416 7284 10468 7336
rect 11888 7352 11940 7404
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 13452 7352 13504 7404
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 17224 7488 17276 7540
rect 14924 7352 14976 7404
rect 17592 7420 17644 7472
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 18696 7352 18748 7404
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 19064 7327 19116 7336
rect 16672 7284 16724 7293
rect 19064 7293 19073 7327
rect 19073 7293 19107 7327
rect 19107 7293 19116 7327
rect 19064 7284 19116 7293
rect 19616 7284 19668 7336
rect 1952 7148 2004 7200
rect 3056 7148 3108 7200
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 4988 7148 5040 7200
rect 5540 7148 5592 7200
rect 7196 7148 7248 7200
rect 8208 7148 8260 7200
rect 10968 7216 11020 7268
rect 11980 7216 12032 7268
rect 14004 7259 14056 7268
rect 14004 7225 14038 7259
rect 14038 7225 14056 7259
rect 14004 7216 14056 7225
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 11520 7148 11572 7200
rect 12624 7148 12676 7200
rect 12808 7148 12860 7200
rect 13084 7148 13136 7200
rect 15476 7216 15528 7268
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 18512 7148 18564 7200
rect 18696 7191 18748 7200
rect 18696 7157 18705 7191
rect 18705 7157 18739 7191
rect 18739 7157 18748 7191
rect 18696 7148 18748 7157
rect 20720 7420 20772 7472
rect 20628 7352 20680 7404
rect 20720 7327 20772 7336
rect 20720 7293 20729 7327
rect 20729 7293 20763 7327
rect 20763 7293 20772 7327
rect 20720 7284 20772 7293
rect 20260 7148 20312 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 4068 6944 4120 6996
rect 7472 6876 7524 6928
rect 1860 6808 1912 6860
rect 2872 6808 2924 6860
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 10600 6944 10652 6996
rect 12440 6944 12492 6996
rect 13176 6944 13228 6996
rect 15384 6944 15436 6996
rect 15752 6944 15804 6996
rect 16304 6944 16356 6996
rect 17316 6944 17368 6996
rect 17960 6944 18012 6996
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 18696 6944 18748 6996
rect 19064 6944 19116 6996
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 5724 6740 5776 6792
rect 7196 6740 7248 6792
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 10048 6876 10100 6928
rect 8300 6740 8352 6792
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 10692 6808 10744 6860
rect 10968 6808 11020 6860
rect 12992 6808 13044 6860
rect 9496 6740 9548 6792
rect 9956 6740 10008 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 12716 6783 12768 6792
rect 10508 6740 10560 6749
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 9680 6672 9732 6724
rect 10048 6672 10100 6724
rect 15200 6808 15252 6860
rect 15384 6808 15436 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 14004 6740 14056 6792
rect 14372 6740 14424 6792
rect 15108 6740 15160 6792
rect 16764 6740 16816 6792
rect 14280 6672 14332 6724
rect 15016 6672 15068 6724
rect 17960 6808 18012 6860
rect 18972 6808 19024 6860
rect 19432 6740 19484 6792
rect 19892 6740 19944 6792
rect 18880 6672 18932 6724
rect 5356 6604 5408 6656
rect 5448 6604 5500 6656
rect 8944 6604 8996 6656
rect 9312 6604 9364 6656
rect 12256 6604 12308 6656
rect 12348 6604 12400 6656
rect 15200 6604 15252 6656
rect 20628 6672 20680 6724
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 19616 6604 19668 6613
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 3056 6400 3108 6452
rect 6736 6400 6788 6452
rect 7104 6400 7156 6452
rect 7472 6400 7524 6452
rect 10508 6400 10560 6452
rect 3792 6332 3844 6384
rect 9588 6375 9640 6384
rect 2872 6264 2924 6316
rect 3056 6264 3108 6316
rect 1768 6196 1820 6248
rect 3424 6196 3476 6248
rect 2504 6128 2556 6180
rect 9588 6341 9597 6375
rect 9597 6341 9631 6375
rect 9631 6341 9640 6375
rect 9588 6332 9640 6341
rect 10968 6332 11020 6384
rect 12072 6332 12124 6384
rect 12256 6400 12308 6452
rect 14004 6400 14056 6452
rect 15016 6400 15068 6452
rect 19156 6400 19208 6452
rect 20536 6400 20588 6452
rect 4160 6264 4212 6316
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 6828 6264 6880 6316
rect 6920 6264 6972 6316
rect 7748 6264 7800 6316
rect 5540 6196 5592 6248
rect 8116 6196 8168 6248
rect 8760 6196 8812 6248
rect 11152 6264 11204 6316
rect 12440 6307 12492 6316
rect 11060 6196 11112 6248
rect 11704 6196 11756 6248
rect 8300 6128 8352 6180
rect 10232 6128 10284 6180
rect 10416 6128 10468 6180
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 13268 6196 13320 6248
rect 14280 6239 14332 6248
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 5356 6060 5408 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 10600 6060 10652 6112
rect 12348 6128 12400 6180
rect 13360 6128 13412 6180
rect 12808 6060 12860 6112
rect 14280 6205 14289 6239
rect 14289 6205 14323 6239
rect 14323 6205 14332 6239
rect 14280 6196 14332 6205
rect 17040 6264 17092 6316
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 19432 6264 19484 6316
rect 19800 6264 19852 6316
rect 19616 6196 19668 6248
rect 15108 6128 15160 6180
rect 16396 6171 16448 6180
rect 16396 6137 16405 6171
rect 16405 6137 16439 6171
rect 16439 6137 16448 6171
rect 16396 6128 16448 6137
rect 17224 6128 17276 6180
rect 17960 6128 18012 6180
rect 15752 6060 15804 6112
rect 18880 6060 18932 6112
rect 19248 6060 19300 6112
rect 19708 6060 19760 6112
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 3148 5856 3200 5908
rect 5264 5856 5316 5908
rect 3516 5788 3568 5840
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2688 5720 2740 5772
rect 6736 5720 6788 5772
rect 2872 5652 2924 5704
rect 2504 5584 2556 5636
rect 3976 5652 4028 5704
rect 6460 5652 6512 5704
rect 7104 5856 7156 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 7196 5763 7248 5772
rect 7196 5729 7230 5763
rect 7230 5729 7248 5763
rect 7196 5720 7248 5729
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 3516 5516 3568 5568
rect 5908 5584 5960 5636
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 6460 5516 6512 5568
rect 9496 5788 9548 5840
rect 12624 5856 12676 5908
rect 17408 5856 17460 5908
rect 9404 5720 9456 5772
rect 9864 5720 9916 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 13360 5788 13412 5840
rect 16856 5788 16908 5840
rect 17040 5788 17092 5840
rect 20536 5856 20588 5908
rect 18696 5788 18748 5840
rect 8576 5652 8628 5704
rect 9588 5652 9640 5704
rect 9772 5652 9824 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11704 5720 11756 5772
rect 12440 5720 12492 5772
rect 12532 5720 12584 5772
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 15752 5720 15804 5772
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 9864 5584 9916 5636
rect 9036 5516 9088 5568
rect 9772 5516 9824 5568
rect 10232 5516 10284 5568
rect 11796 5652 11848 5704
rect 17316 5720 17368 5772
rect 17868 5720 17920 5772
rect 18512 5720 18564 5772
rect 19892 5695 19944 5704
rect 12532 5584 12584 5636
rect 12348 5516 12400 5568
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 19800 5584 19852 5636
rect 13636 5516 13688 5568
rect 15292 5516 15344 5568
rect 16764 5516 16816 5568
rect 17500 5516 17552 5568
rect 19064 5516 19116 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2320 5312 2372 5364
rect 6184 5312 6236 5364
rect 7012 5312 7064 5364
rect 8576 5355 8628 5364
rect 8576 5321 8585 5355
rect 8585 5321 8619 5355
rect 8619 5321 8628 5355
rect 8576 5312 8628 5321
rect 5908 5244 5960 5296
rect 2504 5176 2556 5228
rect 5080 5176 5132 5228
rect 5448 5176 5500 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8300 5244 8352 5296
rect 9036 5219 9088 5228
rect 1676 5108 1728 5160
rect 3976 5108 4028 5160
rect 7104 5040 7156 5092
rect 8208 5108 8260 5160
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9772 5108 9824 5160
rect 11060 5312 11112 5364
rect 12440 5312 12492 5364
rect 14372 5312 14424 5364
rect 16488 5312 16540 5364
rect 17776 5312 17828 5364
rect 19156 5312 19208 5364
rect 21180 5312 21232 5364
rect 12624 5244 12676 5296
rect 13360 5244 13412 5296
rect 11152 5176 11204 5228
rect 11428 5176 11480 5228
rect 18880 5244 18932 5296
rect 11796 5108 11848 5160
rect 14096 5176 14148 5228
rect 15016 5176 15068 5228
rect 15476 5176 15528 5228
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 16856 5176 16908 5228
rect 19064 5176 19116 5228
rect 11152 5040 11204 5092
rect 2780 4972 2832 5024
rect 3240 4972 3292 5024
rect 4988 4972 5040 5024
rect 5540 4972 5592 5024
rect 6092 5015 6144 5024
rect 6092 4981 6101 5015
rect 6101 4981 6135 5015
rect 6135 4981 6144 5015
rect 6092 4972 6144 4981
rect 6276 4972 6328 5024
rect 6736 4972 6788 5024
rect 7012 4972 7064 5024
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7472 4972 7524 5024
rect 8208 4972 8260 5024
rect 8852 4972 8904 5024
rect 9680 4972 9732 5024
rect 10692 4972 10744 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11612 4972 11664 5024
rect 12072 4972 12124 5024
rect 12348 4972 12400 5024
rect 13452 5040 13504 5092
rect 12624 4972 12676 5024
rect 14004 4972 14056 5024
rect 17316 5108 17368 5160
rect 19524 5108 19576 5160
rect 19156 5040 19208 5092
rect 19800 5040 19852 5092
rect 18696 4972 18748 5024
rect 18880 5015 18932 5024
rect 18880 4981 18889 5015
rect 18889 4981 18923 5015
rect 18923 4981 18932 5015
rect 18880 4972 18932 4981
rect 20444 4972 20496 5024
rect 20628 4972 20680 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 3608 4768 3660 4820
rect 4068 4768 4120 4820
rect 9680 4811 9732 4820
rect 5448 4700 5500 4752
rect 1768 4632 1820 4684
rect 3148 4632 3200 4684
rect 3516 4564 3568 4616
rect 6276 4700 6328 4752
rect 6644 4700 6696 4752
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 5356 4496 5408 4548
rect 5080 4428 5132 4480
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 6368 4496 6420 4548
rect 6828 4496 6880 4548
rect 7288 4539 7340 4548
rect 7288 4505 7297 4539
rect 7297 4505 7331 4539
rect 7331 4505 7340 4539
rect 7288 4496 7340 4505
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 7932 4496 7984 4548
rect 8300 4700 8352 4752
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 9772 4768 9824 4820
rect 11980 4768 12032 4820
rect 15016 4768 15068 4820
rect 17868 4768 17920 4820
rect 19800 4811 19852 4820
rect 8208 4632 8260 4684
rect 8300 4564 8352 4616
rect 11336 4700 11388 4752
rect 8944 4632 8996 4684
rect 9772 4632 9824 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 10416 4632 10468 4684
rect 12624 4700 12676 4752
rect 13544 4743 13596 4752
rect 13544 4709 13578 4743
rect 13578 4709 13596 4743
rect 13544 4700 13596 4709
rect 13728 4700 13780 4752
rect 14096 4632 14148 4684
rect 14556 4632 14608 4684
rect 15936 4700 15988 4752
rect 16488 4632 16540 4684
rect 16580 4632 16632 4684
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 9680 4564 9732 4616
rect 9956 4564 10008 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 8668 4496 8720 4548
rect 9496 4496 9548 4548
rect 11428 4564 11480 4616
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 12532 4564 12584 4616
rect 13084 4564 13136 4616
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 16948 4607 17000 4616
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 17408 4564 17460 4616
rect 7380 4428 7432 4480
rect 9772 4428 9824 4480
rect 10968 4428 11020 4480
rect 14556 4428 14608 4480
rect 17316 4428 17368 4480
rect 17500 4428 17552 4480
rect 17960 4700 18012 4752
rect 19800 4777 19809 4811
rect 19809 4777 19843 4811
rect 19843 4777 19852 4811
rect 19800 4768 19852 4777
rect 20444 4700 20496 4752
rect 18972 4632 19024 4684
rect 21640 4632 21692 4684
rect 18420 4607 18472 4616
rect 17776 4496 17828 4548
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 19156 4428 19208 4480
rect 22100 4428 22152 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3148 4267 3200 4276
rect 3148 4233 3157 4267
rect 3157 4233 3191 4267
rect 3191 4233 3200 4267
rect 3148 4224 3200 4233
rect 6920 4224 6972 4276
rect 7288 4224 7340 4276
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 4068 4156 4120 4208
rect 6276 4156 6328 4208
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 5632 4088 5684 4140
rect 6736 4088 6788 4140
rect 9496 4224 9548 4276
rect 10048 4156 10100 4208
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 16488 4224 16540 4276
rect 18512 4224 18564 4276
rect 19064 4224 19116 4276
rect 15660 4156 15712 4208
rect 18052 4156 18104 4208
rect 11888 4088 11940 4140
rect 12900 4088 12952 4140
rect 13176 4088 13228 4140
rect 13268 4088 13320 4140
rect 16948 4088 17000 4140
rect 19064 4088 19116 4140
rect 19800 4131 19852 4140
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 20444 4088 20496 4140
rect 3332 3952 3384 4004
rect 3700 3952 3752 4004
rect 5908 3995 5960 4004
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5448 3884 5500 3936
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 7288 4020 7340 4072
rect 10048 4020 10100 4072
rect 10416 4020 10468 4072
rect 8760 3952 8812 4004
rect 12624 4020 12676 4072
rect 12716 4020 12768 4072
rect 11612 3952 11664 4004
rect 13176 3952 13228 4004
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 18420 4020 18472 4072
rect 14096 3995 14148 4004
rect 14096 3961 14130 3995
rect 14130 3961 14148 3995
rect 14096 3952 14148 3961
rect 14188 3952 14240 4004
rect 16396 3952 16448 4004
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 10692 3884 10744 3936
rect 10876 3884 10928 3936
rect 11796 3884 11848 3936
rect 15108 3884 15160 3936
rect 16672 3884 16724 3936
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 17408 3884 17460 3936
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 18512 3884 18564 3893
rect 18604 3927 18656 3936
rect 18604 3893 18613 3927
rect 18613 3893 18647 3927
rect 18647 3893 18656 3927
rect 19432 3952 19484 4004
rect 18604 3884 18656 3893
rect 19248 3884 19300 3936
rect 19616 3927 19668 3936
rect 19616 3893 19625 3927
rect 19625 3893 19659 3927
rect 19659 3893 19668 3927
rect 19616 3884 19668 3893
rect 20168 3884 20220 3936
rect 20536 3952 20588 4004
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 20628 3884 20680 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3792 3680 3844 3732
rect 4896 3680 4948 3732
rect 6000 3680 6052 3732
rect 7472 3680 7524 3732
rect 8760 3723 8812 3732
rect 8760 3689 8769 3723
rect 8769 3689 8803 3723
rect 8803 3689 8812 3723
rect 8760 3680 8812 3689
rect 9312 3680 9364 3732
rect 10692 3680 10744 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12992 3723 13044 3732
rect 1952 3612 2004 3664
rect 6736 3612 6788 3664
rect 6920 3612 6972 3664
rect 10968 3655 11020 3664
rect 4160 3544 4212 3596
rect 5172 3544 5224 3596
rect 6368 3544 6420 3596
rect 7472 3544 7524 3596
rect 9128 3544 9180 3596
rect 10968 3621 10977 3655
rect 10977 3621 11011 3655
rect 11011 3621 11020 3655
rect 10968 3612 11020 3621
rect 11152 3612 11204 3664
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 16580 3680 16632 3732
rect 17960 3680 18012 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 18880 3680 18932 3732
rect 17132 3612 17184 3664
rect 20076 3680 20128 3732
rect 20812 3612 20864 3664
rect 10140 3544 10192 3596
rect 15476 3544 15528 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 15752 3544 15804 3596
rect 16304 3544 16356 3596
rect 16948 3544 17000 3596
rect 18788 3544 18840 3596
rect 18972 3544 19024 3596
rect 3332 3476 3384 3528
rect 4896 3476 4948 3528
rect 5632 3476 5684 3528
rect 5540 3408 5592 3460
rect 1768 3340 1820 3392
rect 3516 3340 3568 3392
rect 7288 3476 7340 3528
rect 6460 3340 6512 3392
rect 9956 3476 10008 3528
rect 10876 3476 10928 3528
rect 11612 3476 11664 3528
rect 12992 3476 13044 3528
rect 14004 3476 14056 3528
rect 15108 3476 15160 3528
rect 14372 3408 14424 3460
rect 14740 3408 14792 3460
rect 17684 3476 17736 3528
rect 18420 3476 18472 3528
rect 18788 3408 18840 3460
rect 19340 3476 19392 3528
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 8944 3340 8996 3392
rect 10416 3340 10468 3392
rect 11152 3340 11204 3392
rect 13360 3340 13412 3392
rect 16120 3340 16172 3392
rect 19432 3340 19484 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 4896 3179 4948 3188
rect 4896 3145 4905 3179
rect 4905 3145 4939 3179
rect 4939 3145 4948 3179
rect 4896 3136 4948 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8208 3136 8260 3188
rect 4804 3068 4856 3120
rect 7288 3068 7340 3120
rect 7380 3068 7432 3120
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 5080 3000 5132 3052
rect 5264 2932 5316 2984
rect 5448 2932 5500 2984
rect 6460 2932 6512 2984
rect 7012 2932 7064 2984
rect 8760 3068 8812 3120
rect 8852 3000 8904 3052
rect 10048 3068 10100 3120
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 16304 3136 16356 3188
rect 12440 3068 12492 3120
rect 19616 3136 19668 3188
rect 10416 3000 10468 3052
rect 7748 2932 7800 2984
rect 8392 2932 8444 2984
rect 8484 2932 8536 2984
rect 4620 2864 4672 2916
rect 5080 2864 5132 2916
rect 5724 2864 5776 2916
rect 8760 2864 8812 2916
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 10140 2932 10192 2984
rect 10876 2975 10928 2984
rect 10876 2941 10910 2975
rect 10910 2941 10928 2975
rect 10876 2932 10928 2941
rect 11796 3000 11848 3052
rect 12256 2932 12308 2984
rect 4436 2796 4488 2848
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 9680 2796 9732 2848
rect 10968 2864 11020 2916
rect 11060 2864 11112 2916
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 14740 3000 14792 3052
rect 15476 3000 15528 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 17960 3000 18012 3052
rect 19064 3068 19116 3120
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 15384 2975 15436 2984
rect 12808 2864 12860 2916
rect 13728 2864 13780 2916
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 16212 2932 16264 2984
rect 11428 2796 11480 2848
rect 12072 2796 12124 2848
rect 13176 2796 13228 2848
rect 13360 2796 13412 2848
rect 16396 2864 16448 2916
rect 16672 2932 16724 2984
rect 18788 2932 18840 2984
rect 22560 2932 22612 2984
rect 20812 2864 20864 2916
rect 16304 2796 16356 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4160 2592 4212 2644
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 7196 2592 7248 2644
rect 8300 2592 8352 2644
rect 9036 2592 9088 2644
rect 11060 2592 11112 2644
rect 11336 2635 11388 2644
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 13728 2592 13780 2644
rect 15660 2592 15712 2644
rect 16856 2592 16908 2644
rect 18512 2592 18564 2644
rect 18972 2635 19024 2644
rect 18972 2601 18981 2635
rect 18981 2601 19015 2635
rect 19015 2601 19024 2635
rect 18972 2592 19024 2601
rect 2780 2524 2832 2576
rect 2964 2524 3016 2576
rect 6092 2524 6144 2576
rect 6644 2524 6696 2576
rect 11152 2524 11204 2576
rect 12532 2524 12584 2576
rect 5632 2456 5684 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 9864 2456 9916 2508
rect 11704 2456 11756 2508
rect 12440 2456 12492 2508
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 14280 2524 14332 2576
rect 15568 2524 15620 2576
rect 17592 2567 17644 2576
rect 17592 2533 17601 2567
rect 17601 2533 17635 2567
rect 17635 2533 17644 2567
rect 17592 2524 17644 2533
rect 18052 2524 18104 2576
rect 19064 2567 19116 2576
rect 19064 2533 19073 2567
rect 19073 2533 19107 2567
rect 19107 2533 19116 2567
rect 19064 2524 19116 2533
rect 19524 2524 19576 2576
rect 15200 2456 15252 2508
rect 17500 2456 17552 2508
rect 20352 2456 20404 2508
rect 20536 2499 20588 2508
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 6368 2388 6420 2440
rect 8852 2431 8904 2440
rect 8852 2397 8861 2431
rect 8861 2397 8895 2431
rect 8895 2397 8904 2431
rect 8852 2388 8904 2397
rect 10324 2388 10376 2440
rect 10876 2388 10928 2440
rect 11428 2431 11480 2440
rect 11428 2397 11437 2431
rect 11437 2397 11471 2431
rect 11471 2397 11480 2431
rect 11428 2388 11480 2397
rect 17960 2388 18012 2440
rect 18788 2388 18840 2440
rect 7104 2320 7156 2372
rect 18972 2320 19024 2372
rect 2412 2252 2464 2304
rect 7748 2252 7800 2304
rect 15844 2252 15896 2304
rect 19156 2252 19208 2304
rect 20720 2295 20772 2304
rect 20720 2261 20729 2295
rect 20729 2261 20763 2295
rect 20763 2261 20772 2295
rect 20720 2252 20772 2261
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 17040 2048 17092 2100
rect 18604 2048 18656 2100
rect 11336 1980 11388 2032
rect 11980 1980 12032 2032
rect 1492 1844 1544 1896
rect 8392 1844 8444 1896
rect 572 1776 624 1828
rect 8576 1776 8628 1828
rect 204 1640 256 1692
rect 5816 1640 5868 1692
rect 1032 1504 1084 1556
rect 8484 1504 8536 1556
rect 3884 1096 3936 1148
rect 5448 1096 5500 1148
<< metal2 >>
rect 2962 22536 3018 22545
rect 2962 22471 3018 22480
rect 2502 22128 2558 22137
rect 2502 22063 2558 22072
rect 2410 21176 2466 21185
rect 2410 21111 2466 21120
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1964 18970 1992 19207
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18864 2006 18873
rect 1492 18828 1544 18834
rect 1950 18799 2006 18808
rect 1492 18770 1544 18776
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1412 12374 1440 13330
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 1504 7478 1532 18770
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1674 18320 1730 18329
rect 1674 18255 1730 18264
rect 1688 17610 1716 18255
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 17814 1808 18158
rect 1950 17912 2006 17921
rect 1950 17847 2006 17856
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1858 17368 1914 17377
rect 1964 17338 1992 17847
rect 1858 17303 1914 17312
rect 1952 17332 2004 17338
rect 1872 16794 1900 17303
rect 1952 17274 2004 17280
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 2424 15706 2452 21111
rect 2516 16250 2544 22063
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2792 19174 2820 20159
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2792 15162 2820 15535
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 1952 15088 2004 15094
rect 1950 15056 1952 15065
rect 2004 15056 2006 15065
rect 1950 14991 2006 15000
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1674 14648 1730 14657
rect 1674 14583 1676 14592
rect 1728 14583 1730 14592
rect 1676 14554 1728 14560
rect 1780 14550 1808 14894
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1582 14104 1638 14113
rect 1582 14039 1638 14048
rect 1596 13530 1624 14039
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 10810 1716 12242
rect 1872 12102 1900 14418
rect 2424 14074 2452 14962
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2424 13938 2452 14010
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 10130 1808 11154
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1872 9586 1900 11494
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2056 10130 2084 10202
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1872 6866 1900 8366
rect 2148 7546 2176 13874
rect 2884 13530 2912 14418
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2332 12442 2360 13330
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12986 2544 13262
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2976 12850 3004 22471
rect 5722 22320 5778 22800
rect 17130 22320 17186 22800
rect 17958 22536 18014 22545
rect 17958 22471 18014 22480
rect 3422 21584 3478 21593
rect 3422 21519 3478 21528
rect 3330 16960 3386 16969
rect 3330 16895 3386 16904
rect 3344 16250 3372 16895
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3160 15638 3188 15982
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3436 14618 3464 21519
rect 3882 20632 3938 20641
rect 3882 20567 3938 20576
rect 3896 19514 3924 20567
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3160 12889 3188 13738
rect 3146 12880 3202 12889
rect 2964 12844 3016 12850
rect 3146 12815 3148 12824
rect 2964 12786 3016 12792
rect 3200 12815 3202 12824
rect 3148 12786 3200 12792
rect 2976 12646 3004 12786
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2240 8090 2268 11494
rect 2332 9178 2360 11494
rect 2424 11218 2452 11630
rect 2792 11354 2820 12242
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2412 11212 2464 11218
rect 2464 11172 2544 11200
rect 2412 11154 2464 11160
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 9722 2452 10406
rect 2516 10266 2544 11172
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9586 2544 10202
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2608 8634 2636 10134
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2700 8974 2728 9522
rect 2884 9518 2912 11494
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2976 9382 3004 11562
rect 3068 9466 3096 12650
rect 3160 12238 3188 12786
rect 3252 12306 3280 13806
rect 3344 13530 3372 14350
rect 3804 13734 3832 14826
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14414 4200 14758
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3792 13728 3844 13734
rect 3514 13696 3570 13705
rect 3792 13670 3844 13676
rect 3514 13631 3570 13640
rect 3528 13530 3556 13631
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3804 13326 3832 13670
rect 4080 13512 4108 13874
rect 4172 13870 4200 14350
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4080 13484 4200 13512
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3424 13320 3476 13326
rect 3792 13320 3844 13326
rect 3424 13262 3476 13268
rect 3606 13288 3662 13297
rect 3436 12986 3464 13262
rect 3792 13262 3844 13268
rect 3606 13223 3662 13232
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3620 12442 3648 13223
rect 3896 12986 3924 13330
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3700 12776 3752 12782
rect 3988 12753 4016 13194
rect 4080 12918 4108 13330
rect 4172 12918 4200 13484
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 3700 12718 3752 12724
rect 3974 12744 4030 12753
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3606 12336 3662 12345
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3516 12300 3568 12306
rect 3606 12271 3662 12280
rect 3516 12242 3568 12248
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10810 3188 10950
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3252 9518 3280 12106
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 9654 3372 11494
rect 3436 10554 3464 11698
rect 3528 11082 3556 12242
rect 3620 11150 3648 12271
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3528 10674 3556 11018
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 10554 3648 10610
rect 3436 10526 3648 10554
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3240 9512 3292 9518
rect 3068 9438 3188 9466
rect 3240 9454 3292 9460
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9194 3096 9318
rect 2976 9166 3096 9194
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2596 8356 2648 8362
rect 2700 8344 2728 8910
rect 2648 8316 2728 8344
rect 2596 8298 2648 8304
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2608 7886 2636 8298
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1860 6860 1912 6866
rect 1780 6820 1860 6848
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 5166 1716 6734
rect 1780 6254 1808 6820
rect 1860 6802 1912 6808
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1780 4690 1808 6190
rect 1964 5914 1992 7142
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1780 4146 1808 4626
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1780 3398 1808 4082
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1492 1896 1544 1902
rect 1492 1838 1544 1844
rect 572 1828 624 1834
rect 572 1770 624 1776
rect 204 1692 256 1698
rect 204 1634 256 1640
rect 216 480 244 1634
rect 584 480 612 1770
rect 1032 1556 1084 1562
rect 1032 1498 1084 1504
rect 1044 480 1072 1498
rect 1504 480 1532 1838
rect 1964 480 1992 3606
rect 2240 2009 2268 7822
rect 2700 7750 2728 7890
rect 2884 7818 2912 8910
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2332 5370 2360 5714
rect 2516 5642 2544 6122
rect 2700 5778 2728 7686
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6322 2912 6802
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2516 5234 2544 5578
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2700 2553 2728 5714
rect 2884 5710 2912 6258
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 3505 2820 4966
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2792 2582 2820 2751
rect 2780 2576 2832 2582
rect 2686 2544 2742 2553
rect 2780 2518 2832 2524
rect 2686 2479 2742 2488
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 2424 480 2452 2246
rect 2884 480 2912 3567
rect 2976 2582 3004 9166
rect 3160 9042 3188 9438
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6458 3096 7142
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3068 6118 3096 6258
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3160 5914 3188 8978
rect 3148 5908 3200 5914
rect 3068 5868 3148 5896
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 3068 1601 3096 5868
rect 3148 5850 3200 5856
rect 3252 5030 3280 9454
rect 3528 8634 3556 10406
rect 3620 10198 3648 10526
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3620 9518 3648 10134
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 7886 3648 8434
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 6254 3464 7142
rect 3528 6662 3556 7346
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3528 5846 3556 6598
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4282 3188 4626
rect 3528 4622 3556 5510
rect 3620 4826 3648 7822
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3344 3534 3372 3946
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3528 3398 3556 4558
rect 3712 4010 3740 12718
rect 3974 12679 4030 12688
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 9330 3832 12582
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3988 11801 4016 12310
rect 4068 12232 4120 12238
rect 4172 12220 4200 12854
rect 4120 12192 4200 12220
rect 4068 12174 4120 12180
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 10606 3924 11494
rect 4080 11218 4108 12174
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 10674 4016 10775
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4080 10606 4108 11154
rect 4172 11014 4200 11562
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3988 9722 4016 10367
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9926 4108 9959
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4066 9480 4122 9489
rect 4066 9415 4068 9424
rect 4120 9415 4122 9424
rect 4068 9386 4120 9392
rect 3804 9302 3924 9330
rect 3896 8430 3924 9302
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4080 8537 4108 9046
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3804 7206 3832 8026
rect 3896 7274 3924 8366
rect 4172 8090 4200 10474
rect 4264 10266 4292 15506
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4724 13326 4752 15914
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4434 12880 4490 12889
rect 4724 12832 4752 13126
rect 4434 12815 4436 12824
rect 4488 12815 4490 12824
rect 4436 12786 4488 12792
rect 4632 12804 4752 12832
rect 4632 12646 4660 12804
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4448 8294 4476 8502
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4540 7954 4568 8434
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4160 7880 4212 7886
rect 4620 7880 4672 7886
rect 4160 7822 4212 7828
rect 4618 7848 4620 7857
rect 4672 7848 4674 7857
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4080 7478 4108 7511
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3804 6390 3832 7142
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3804 4162 3832 6326
rect 3988 6066 4016 7346
rect 4066 7168 4122 7177
rect 4172 7154 4200 7822
rect 4618 7783 4674 7792
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4172 7126 4292 7154
rect 4066 7103 4122 7112
rect 4080 7002 4108 7103
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4172 6066 4200 6258
rect 3988 6038 4200 6066
rect 3988 5710 4016 6038
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3988 4865 4016 5102
rect 3974 4856 4030 4865
rect 3974 4791 4030 4800
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4321 4108 4762
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4068 4208 4120 4214
rect 3804 4134 3924 4162
rect 4068 4150 4120 4156
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3738 3832 3878
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3896 3618 3924 4134
rect 3620 3590 3924 3618
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3058 3556 3334
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3422 2816 3478 2825
rect 3422 2751 3478 2760
rect 3054 1592 3110 1601
rect 3054 1527 3110 1536
rect 3436 1442 3464 2751
rect 3344 1414 3464 1442
rect 3344 480 3372 1414
rect 3620 649 3648 3590
rect 4080 3516 4108 4150
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3712 3488 4108 3516
rect 3606 640 3662 649
rect 3606 575 3662 584
rect 3712 480 3740 3488
rect 4172 2650 4200 3538
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4264 2530 4292 7126
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4448 2650 4476 2790
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4172 2502 4292 2530
rect 3884 1148 3936 1154
rect 3884 1090 3936 1096
rect 3896 1057 3924 1090
rect 3882 1048 3938 1057
rect 3882 983 3938 992
rect 4172 480 4200 2502
rect 4632 2446 4660 2858
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1442 4752 12650
rect 4816 9654 4844 13806
rect 4908 12306 4936 16594
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4802 8936 4858 8945
rect 4802 8871 4858 8880
rect 4816 8022 4844 8871
rect 4908 8634 4936 11562
rect 5000 11014 5028 19246
rect 5644 18902 5672 19246
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5736 18222 5764 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 13802 5120 15438
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 13530 5120 13738
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5184 11626 5212 15370
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5276 11762 5304 13942
rect 5368 11898 5396 14418
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12714 5488 13262
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 12442 5488 12650
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 8294 4936 8570
rect 5000 8566 5028 10950
rect 5276 10690 5304 11698
rect 5368 11694 5396 11834
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5460 11626 5488 12242
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5828 11558 5856 11698
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5184 10662 5304 10690
rect 5184 10538 5212 10662
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8906 5120 9522
rect 5184 8974 5212 10474
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4816 3126 4844 7958
rect 5000 7206 5028 8026
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 5030 5028 7142
rect 5092 5352 5120 8842
rect 5184 8022 5212 8910
rect 5276 8090 5304 10474
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7410 5212 7958
rect 5368 7546 5396 10202
rect 5460 9994 5488 10746
rect 5552 10062 5580 11018
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10198 5764 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5644 9178 5672 10066
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5540 8424 5592 8430
rect 5538 8392 5540 8401
rect 5592 8392 5594 8401
rect 5538 8327 5594 8336
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5644 7721 5672 7890
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5630 7712 5686 7721
rect 5630 7647 5686 7656
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5368 6118 5396 6598
rect 5460 6322 5488 6598
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5552 6254 5580 7142
rect 5736 6798 5764 7822
rect 5920 7546 5948 14894
rect 6012 13530 6040 18770
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6012 11558 6040 12174
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 11354 6040 11494
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6012 10130 6040 11290
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6104 10033 6132 19178
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6196 10674 6224 11766
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6090 10024 6146 10033
rect 6090 9959 6146 9968
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5092 5324 5304 5352
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3738 4936 3878
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4908 3194 4936 3470
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4632 1414 4752 1442
rect 4632 480 4660 1414
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2410 0 2466 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3698 0 3754 480
rect 4158 0 4214 480
rect 4618 0 4674 480
rect 5000 241 5028 4966
rect 5092 4486 5120 5170
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5092 4146 5120 4422
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3058 5120 4082
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3194 5212 3538
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5276 2990 5304 5324
rect 5460 5234 5488 5510
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4758 5488 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5092 480 5120 2858
rect 5368 1034 5396 4490
rect 5552 4026 5580 4966
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5460 3998 5580 4026
rect 5460 3942 5488 3998
rect 5448 3936 5500 3942
rect 5644 3890 5672 4082
rect 5448 3878 5500 3884
rect 5552 3862 5672 3890
rect 5552 3466 5580 3862
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 1154 5488 2926
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2009 5580 2790
rect 5644 2514 5672 3470
rect 5736 2922 5764 6734
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5814 5808 5870 5817
rect 5814 5743 5870 5752
rect 5828 4185 5856 5743
rect 5920 5642 5948 6054
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5998 5264 6054 5273
rect 5814 4176 5870 4185
rect 5814 4111 5870 4120
rect 5920 4010 5948 5238
rect 5998 5199 6054 5208
rect 6012 4570 6040 5199
rect 6104 5030 6132 9959
rect 6196 9042 6224 10066
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6288 8022 6316 8230
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6012 4542 6132 4570
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 6012 3738 6040 4422
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5814 3360 5870 3369
rect 5814 3295 5870 3304
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5828 1698 5856 3295
rect 6104 2582 6132 4542
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 5816 1692 5868 1698
rect 5816 1634 5868 1640
rect 5448 1148 5500 1154
rect 5448 1090 5500 1096
rect 5368 1006 5580 1034
rect 5552 480 5580 1006
rect 6196 898 6224 5306
rect 6288 5030 6316 7482
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6288 4214 6316 4694
rect 6380 4690 6408 8774
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6472 7818 6500 8298
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6564 7750 6592 11698
rect 6748 9654 6776 17682
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13530 6868 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 9466 6868 11290
rect 6932 10470 6960 12242
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 9586 6960 10406
rect 7024 10266 7052 12718
rect 7116 12102 7144 17070
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13462 7236 14214
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7300 13394 7328 13942
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7194 13288 7250 13297
rect 7194 13223 7196 13232
rect 7248 13223 7250 13232
rect 7196 13194 7248 13200
rect 7392 12170 7420 17614
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10192 7156 10198
rect 7024 10140 7104 10146
rect 7024 10134 7156 10140
rect 7024 10118 7144 10134
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6748 9438 6868 9466
rect 6748 9042 6776 9438
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8514 6776 8978
rect 6932 8566 6960 9318
rect 6920 8560 6972 8566
rect 6748 8486 6868 8514
rect 6920 8502 6972 8508
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6550 6624 6606 6633
rect 6550 6559 6606 6568
rect 6460 5704 6512 5710
rect 6564 5692 6592 6559
rect 6512 5664 6592 5692
rect 6460 5646 6512 5652
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4554 6408 4626
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6472 3913 6500 5510
rect 6458 3904 6514 3913
rect 6458 3839 6514 3848
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6274 3496 6330 3505
rect 6274 3431 6330 3440
rect 6288 2825 6316 3431
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 6288 2650 6316 2751
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6380 2446 6408 3538
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 2990 6500 3334
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6564 2836 6592 5664
rect 6656 4758 6684 7482
rect 6748 6458 6776 8366
rect 6840 7818 6868 8486
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 7018 6868 7754
rect 6840 6990 6960 7018
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6840 6322 6868 6802
rect 6932 6322 6960 6990
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6734 5808 6790 5817
rect 6734 5743 6736 5752
rect 6788 5743 6790 5752
rect 6736 5714 6788 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6644 4752 6696 4758
rect 6748 4729 6776 4966
rect 6644 4694 6696 4700
rect 6734 4720 6790 4729
rect 6734 4655 6790 4664
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6472 2808 6592 2836
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6012 870 6224 898
rect 6012 480 6040 870
rect 6472 480 6500 2808
rect 6656 2582 6684 3975
rect 6748 3670 6776 4082
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6840 480 6868 4490
rect 6932 4282 6960 5646
rect 7024 5370 7052 10118
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 9042 7236 9454
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7300 8922 7328 12106
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 10577 7420 11562
rect 7484 11218 7512 16050
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 13938 7604 14282
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7576 13394 7604 13874
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7576 12442 7604 13330
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7668 11898 7696 14350
rect 7760 12442 7788 14486
rect 8220 14346 8248 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 15638 12848 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 13297 7880 13330
rect 7838 13288 7894 13297
rect 7838 13223 7894 13232
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 12170 8064 12242
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 11354 7788 12038
rect 7944 11626 7972 12106
rect 8036 11762 8064 12106
rect 8496 11830 8524 13738
rect 8680 12918 8708 13806
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 12753 9720 12786
rect 9678 12744 9734 12753
rect 9588 12708 9640 12714
rect 9678 12679 9734 12688
rect 9588 12650 9640 12656
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 8668 12232 8720 12238
rect 8720 12180 8892 12186
rect 8668 12174 8892 12180
rect 8680 12170 8892 12174
rect 8680 12164 8904 12170
rect 8680 12158 8852 12164
rect 8852 12106 8904 12112
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7378 10568 7434 10577
rect 7378 10503 7434 10512
rect 7392 10198 7420 10503
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7208 8894 7328 8922
rect 7208 7818 7236 8894
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7206 7236 7754
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7116 5914 7144 6394
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7208 5778 7236 6734
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6932 3194 6960 3606
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 2990 7052 4966
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7116 2378 7144 5034
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 2650 7236 4966
rect 7300 4554 7328 8774
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 8090 7420 8434
rect 7484 8378 7512 10202
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9654 7604 10066
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7576 9178 7604 9590
rect 7668 9518 7696 11018
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10742 7880 10950
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7760 10266 7788 10474
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 11630
rect 8496 11558 8524 11766
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8312 11286 8340 11494
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8496 10810 8524 11494
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7760 9586 7788 10202
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8498 7604 9114
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7484 8350 7604 8378
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7484 7410 7512 8230
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7484 6934 7512 7346
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7484 6458 7512 6870
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 5030 7512 5170
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 4078 7328 4218
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7300 3534 7328 4014
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7300 3233 7328 3470
rect 7286 3224 7342 3233
rect 7286 3159 7342 3168
rect 7392 3126 7420 4422
rect 7484 3738 7512 4966
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 3602 7512 3674
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7300 480 7328 3062
rect 7576 1986 7604 8350
rect 7668 7886 7696 8978
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7852 8537 7880 8570
rect 7838 8528 7894 8537
rect 7838 8463 7894 8472
rect 8128 8430 8156 8842
rect 8220 8634 8248 10066
rect 8496 9994 8524 10746
rect 9324 10470 9352 12378
rect 9600 11744 9628 12650
rect 9784 12238 9812 13942
rect 9876 12442 9904 14418
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10140 13864 10192 13870
rect 10060 13824 10140 13852
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 12646 9996 13398
rect 10060 12850 10088 13824
rect 10140 13806 10192 13812
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12850 10180 13262
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 10152 12374 10180 12582
rect 10336 12442 10364 13126
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9508 11716 9628 11744
rect 9508 11257 9536 11716
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9494 11248 9550 11257
rect 9494 11183 9550 11192
rect 9600 10674 9628 11562
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8496 9586 8524 9930
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8312 8838 8340 9318
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7654 7440 7710 7449
rect 7654 7375 7710 7384
rect 7668 7342 7696 7375
rect 8220 7342 8248 8570
rect 8404 7546 8432 8978
rect 8496 8974 8524 9318
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8668 8968 8720 8974
rect 9048 8945 9076 8978
rect 8668 8910 8720 8916
rect 9034 8936 9090 8945
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8496 7721 8524 7890
rect 8482 7712 8538 7721
rect 8482 7647 8538 7656
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 4604 7788 6258
rect 8116 6248 8168 6254
rect 8220 6236 8248 7142
rect 8300 6792 8352 6798
rect 8496 6769 8524 7647
rect 8588 7324 8616 8366
rect 8680 7857 8708 8910
rect 9034 8871 9090 8880
rect 8666 7848 8722 7857
rect 8666 7783 8722 7792
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8668 7336 8720 7342
rect 8588 7296 8668 7324
rect 8720 7296 8800 7324
rect 8668 7278 8720 7284
rect 8300 6734 8352 6740
rect 8482 6760 8538 6769
rect 8168 6208 8248 6236
rect 8116 6190 8168 6196
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5166 8248 6208
rect 8312 6186 8340 6734
rect 8482 6695 8538 6704
rect 8772 6254 8800 7296
rect 8864 6866 8892 7783
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8760 6248 8812 6254
rect 8864 6225 8892 6802
rect 8944 6792 8996 6798
rect 8996 6752 9076 6780
rect 8944 6734 8996 6740
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8760 6190 8812 6196
rect 8850 6216 8906 6225
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5574 8340 6122
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5302 8340 5510
rect 8588 5370 8616 5646
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8208 5024 8260 5030
rect 8772 5012 8800 6190
rect 8850 6151 8906 6160
rect 8956 5914 8984 6598
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9048 5794 9076 6752
rect 8956 5766 9076 5794
rect 8852 5024 8904 5030
rect 8208 4966 8260 4972
rect 8390 4992 8446 5001
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8220 4842 8248 4966
rect 8772 4984 8852 5012
rect 8852 4966 8904 4972
rect 8390 4927 8446 4936
rect 8220 4814 8340 4842
rect 8312 4758 8340 4814
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7840 4616 7892 4622
rect 7760 4576 7840 4604
rect 7840 4558 7892 4564
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7944 4049 7972 4490
rect 7930 4040 7986 4049
rect 7930 3975 7986 3984
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3194 8248 4626
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 2310 7788 2926
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8312 2650 8340 4558
rect 8404 2990 8432 4927
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 3913 8708 4490
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8666 3904 8722 3913
rect 8666 3839 8722 3848
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8574 2952 8630 2961
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8206 2408 8262 2417
rect 8206 2343 8262 2352
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7576 1958 7788 1986
rect 7760 480 7788 1958
rect 8220 480 8248 2343
rect 8404 1902 8432 2790
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8496 1562 8524 2926
rect 8574 2887 8630 2896
rect 8588 2514 8616 2887
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8588 1834 8616 2450
rect 8576 1828 8628 1834
rect 8576 1770 8628 1776
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8680 480 8708 3839
rect 8772 3738 8800 3946
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8772 3126 8800 3674
rect 8864 3380 8892 4966
rect 8956 4690 8984 5766
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5234 9076 5510
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9034 5128 9090 5137
rect 9034 5063 9090 5072
rect 9048 4729 9076 5063
rect 9034 4720 9090 4729
rect 8944 4684 8996 4690
rect 9034 4655 9090 4664
rect 8944 4626 8996 4632
rect 8956 3641 8984 4626
rect 8942 3632 8998 3641
rect 8942 3567 8998 3576
rect 8944 3392 8996 3398
rect 8864 3352 8944 3380
rect 8944 3334 8996 3340
rect 8956 3233 8984 3334
rect 8942 3224 8998 3233
rect 8942 3159 8998 3168
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 2825 8800 2858
rect 8758 2816 8814 2825
rect 8758 2751 8814 2760
rect 8864 2446 8892 2994
rect 8956 2990 8984 3159
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9048 2650 9076 4655
rect 9140 3602 9168 9998
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 7886 9260 8298
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7546 9260 7822
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 6746 9352 10406
rect 9600 10266 9628 10610
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9692 10198 9720 10950
rect 9784 10810 9812 11154
rect 10244 11150 10272 11494
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10152 10810 10180 11086
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10324 10464 10376 10470
rect 10322 10432 10324 10441
rect 10376 10432 10378 10441
rect 10322 10367 10378 10376
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 10060 9722 10088 10231
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9722 10272 10066
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9770 9208 9826 9217
rect 9770 9143 9826 9152
rect 9784 9110 9812 9143
rect 9772 9104 9824 9110
rect 9586 9072 9642 9081
rect 9772 9046 9824 9052
rect 9586 9007 9642 9016
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8362 9444 8910
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8498 9536 8774
rect 9600 8566 9628 9007
rect 9678 8936 9734 8945
rect 9876 8906 9904 9386
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9678 8871 9680 8880
rect 9732 8871 9734 8880
rect 9864 8900 9916 8906
rect 9680 8842 9732 8848
rect 9864 8842 9916 8848
rect 9876 8634 9904 8842
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9770 8528 9826 8537
rect 9496 8492 9548 8498
rect 9770 8463 9826 8472
rect 9496 8434 9548 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9232 6718 9352 6746
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9232 3482 9260 6718
rect 9312 6656 9364 6662
rect 9310 6624 9312 6633
rect 9364 6624 9366 6633
rect 9310 6559 9366 6568
rect 9508 5846 9536 6734
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9496 5840 9548 5846
rect 9402 5808 9458 5817
rect 9496 5782 9548 5788
rect 9402 5743 9404 5752
rect 9456 5743 9458 5752
rect 9404 5714 9456 5720
rect 9416 4162 9444 5714
rect 9508 4554 9536 5782
rect 9600 5710 9628 6326
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9692 5522 9720 6666
rect 9784 5710 9812 8463
rect 9968 8022 9996 8978
rect 10046 8120 10102 8129
rect 10046 8055 10102 8064
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 10060 7954 10088 8055
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10152 7546 10180 9046
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10244 8090 10272 8366
rect 10336 8090 10364 8502
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 7970 10456 13398
rect 10520 12986 10548 14350
rect 11164 14074 11192 14350
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10980 13326 11008 13738
rect 11164 13462 11192 14010
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10968 13320 11020 13326
rect 11072 13308 11100 13398
rect 11256 13308 11284 13738
rect 11716 13530 11744 14554
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 13870 12480 14418
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11072 13280 11284 13308
rect 10968 13262 11020 13268
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10520 12714 10548 12786
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10612 12646 10640 12922
rect 10704 12850 10732 13262
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12918 10824 13194
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10612 11898 10640 12310
rect 10980 12306 11008 13262
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11898 10732 12106
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10980 11558 11008 12242
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9722 10548 10406
rect 10796 9722 10824 11222
rect 10980 11218 11008 11494
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10874 10160 10930 10169
rect 10874 10095 10930 10104
rect 10888 9926 10916 10095
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9081 10732 9454
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 9178 10916 9386
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10690 9072 10746 9081
rect 10690 9007 10746 9016
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10704 8430 10732 8570
rect 10692 8424 10744 8430
rect 10506 8392 10562 8401
rect 10692 8366 10744 8372
rect 10506 8327 10562 8336
rect 10336 7942 10456 7970
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9862 6080 9918 6089
rect 9862 6015 9918 6024
rect 9876 5778 9904 6015
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9600 5494 9720 5522
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9600 5001 9628 5494
rect 9784 5166 9812 5510
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 5024 9732 5030
rect 9586 4992 9642 5001
rect 9680 4966 9732 4972
rect 9586 4927 9642 4936
rect 9692 4826 9720 4966
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9784 4690 9812 4762
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9508 4282 9536 4490
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9416 4134 9628 4162
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3738 9352 3878
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9140 3454 9260 3482
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9140 480 9168 3454
rect 9600 480 9628 4134
rect 9692 2854 9720 4558
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4146 9812 4422
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9876 2514 9904 5578
rect 9968 4865 9996 6734
rect 10060 6730 10088 6870
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10244 6186 10272 7822
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10138 5808 10194 5817
rect 10048 5772 10100 5778
rect 10138 5743 10194 5752
rect 10048 5714 10100 5720
rect 10060 5681 10088 5714
rect 10152 5710 10180 5743
rect 10140 5704 10192 5710
rect 10046 5672 10102 5681
rect 10140 5646 10192 5652
rect 10046 5607 10102 5616
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9968 4622 9996 4791
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10060 4214 10088 4626
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3534 9996 4082
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10060 3126 10088 4014
rect 10152 3602 10180 4558
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10152 2990 10180 3538
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10244 2836 10272 5510
rect 9968 2808 10272 2836
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9968 480 9996 2808
rect 10336 2446 10364 7942
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7342 10456 7822
rect 10520 7750 10548 8327
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 6780 10456 7278
rect 10520 6882 10548 7686
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 7002 10640 7142
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10520 6854 10640 6882
rect 10704 6866 10732 8366
rect 10508 6792 10560 6798
rect 10428 6752 10508 6780
rect 10508 6734 10560 6740
rect 10520 6458 10548 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10612 6338 10640 6854
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10520 6310 10640 6338
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10428 4690 10456 6122
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3398 10456 4014
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10428 3058 10456 3334
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10520 2938 10548 6310
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10428 2910 10548 2938
rect 10612 2938 10640 6054
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 3942 10732 4966
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10704 3233 10732 3674
rect 10690 3224 10746 3233
rect 10690 3159 10746 3168
rect 10796 3097 10824 8978
rect 10888 5681 10916 9114
rect 10980 8022 11008 10474
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 8673 11100 9998
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 10980 7274 11008 7958
rect 11060 7948 11112 7954
rect 11164 7936 11192 13280
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11808 12940 12112 12968
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10674 11652 12582
rect 11716 11914 11744 12650
rect 11808 12102 11836 12940
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11900 12306 11928 12786
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11716 11886 11836 11914
rect 11900 11898 11928 12242
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11716 10554 11744 11766
rect 11624 10526 11744 10554
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11244 9512 11296 9518
rect 11242 9480 11244 9489
rect 11296 9480 11298 9489
rect 11242 9415 11298 9424
rect 11348 9178 11376 9590
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7954 11376 8298
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11112 7908 11192 7936
rect 11336 7948 11388 7954
rect 11060 7890 11112 7896
rect 11336 7890 11388 7896
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11072 6905 11100 7890
rect 11440 7818 11468 8026
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11520 7200 11572 7206
rect 11518 7168 11520 7177
rect 11572 7168 11574 7177
rect 11518 7103 11574 7112
rect 11058 6896 11114 6905
rect 10968 6860 11020 6866
rect 11058 6831 11114 6840
rect 10968 6802 11020 6808
rect 10980 6390 11008 6802
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10874 5672 10930 5681
rect 10874 5607 10930 5616
rect 11072 5522 11100 6190
rect 10980 5494 11100 5522
rect 10980 5148 11008 5494
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5273 11100 5306
rect 11058 5264 11114 5273
rect 11164 5234 11192 6258
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11518 5264 11574 5273
rect 11058 5199 11114 5208
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11428 5228 11480 5234
rect 11518 5199 11574 5208
rect 11428 5170 11480 5176
rect 10980 5120 11100 5148
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3534 10916 3878
rect 10980 3670 11008 4422
rect 11072 3777 11100 5120
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11058 3768 11114 3777
rect 11058 3703 11114 3712
rect 11164 3670 11192 5034
rect 11336 4752 11388 4758
rect 11334 4720 11336 4729
rect 11388 4720 11390 4729
rect 11334 4655 11390 4664
rect 11440 4622 11468 5170
rect 11532 5030 11560 5199
rect 11624 5030 11652 10526
rect 11808 10470 11836 11886
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11716 9908 11744 10406
rect 11808 10062 11836 10406
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11796 9920 11848 9926
rect 11716 9880 11796 9908
rect 11796 9862 11848 9868
rect 11808 7993 11836 9862
rect 11900 8362 11928 11698
rect 11992 10266 12020 12786
rect 12084 12646 12112 12940
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 12238 12112 12582
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12176 11778 12204 12854
rect 12360 12782 12388 13126
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12084 11750 12204 11778
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12084 10146 12112 11750
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11393 12204 11630
rect 12162 11384 12218 11393
rect 12162 11319 12218 11328
rect 12268 11286 12296 12106
rect 12360 11830 12388 12718
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11280 12308 11286
rect 12162 11248 12218 11257
rect 12256 11222 12308 11228
rect 12162 11183 12218 11192
rect 12176 10810 12204 11183
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10674 12296 11222
rect 12360 10742 12388 11494
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12452 10606 12480 11222
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11992 10118 12112 10146
rect 12452 10146 12480 10542
rect 12544 10248 12572 15506
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12728 12850 12756 14826
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 13394 13124 13806
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12458 12756 12786
rect 12820 12714 12848 13262
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12728 12442 12848 12458
rect 13004 12442 13032 13194
rect 12728 12436 12860 12442
rect 12728 12430 12808 12436
rect 12808 12378 12860 12384
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12820 12347 12848 12378
rect 12992 12232 13044 12238
rect 13044 12192 13124 12220
rect 12992 12174 13044 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11694 12848 12038
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12806 11384 12862 11393
rect 13004 11354 13032 11698
rect 13096 11558 13124 12192
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12806 11319 12862 11328
rect 12992 11348 13044 11354
rect 12622 10568 12678 10577
rect 12622 10503 12624 10512
rect 12676 10503 12678 10512
rect 12624 10474 12676 10480
rect 12624 10260 12676 10266
rect 12544 10220 12624 10248
rect 12624 10202 12676 10208
rect 12452 10118 12572 10146
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11794 7984 11850 7993
rect 11794 7919 11850 7928
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11716 6254 11744 7754
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11428 4616 11480 4622
rect 11480 4576 11652 4604
rect 11428 4558 11480 4564
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4010 11652 4576
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11624 3534 11652 3946
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 10782 3088 10838 3097
rect 10782 3023 10838 3032
rect 10888 2990 10916 3470
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11164 3176 11192 3334
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11072 3108 11100 3159
rect 11164 3148 11376 3176
rect 11072 3080 11192 3108
rect 10876 2984 10928 2990
rect 10612 2910 10824 2938
rect 10876 2926 10928 2932
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10428 480 10456 2910
rect 10796 2802 10824 2910
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10980 2802 11008 2858
rect 10796 2774 11008 2802
rect 11072 2650 11100 2858
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11164 2582 11192 3080
rect 11348 2650 11376 3148
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11440 2446 11468 2790
rect 11716 2514 11744 5714
rect 11808 5710 11836 7754
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11808 3942 11836 5102
rect 11900 4264 11928 7346
rect 11992 7274 12020 10118
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12084 8090 12112 9998
rect 12162 8936 12218 8945
rect 12162 8871 12218 8880
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11992 7177 12020 7210
rect 11978 7168 12034 7177
rect 11978 7103 12034 7112
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11992 4826 12020 6559
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 12084 5545 12112 6326
rect 12070 5536 12126 5545
rect 12070 5471 12126 5480
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11900 4236 12020 4264
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11900 3738 11928 4082
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 10888 480 10916 2382
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11348 480 11376 1974
rect 11808 480 11836 2994
rect 11992 2038 12020 4236
rect 12084 2938 12112 4966
rect 12176 4536 12204 8871
rect 12268 8634 12296 9998
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12268 8498 12296 8570
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12360 8106 12388 9046
rect 12452 8634 12480 9998
rect 12544 9518 12572 10118
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12544 8566 12572 9114
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12728 8498 12756 9046
rect 12820 8537 12848 11319
rect 12992 11290 13044 11296
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10470 12940 10950
rect 13004 10606 13032 11290
rect 13556 11286 13584 14214
rect 14292 12986 14320 14418
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14752 14074 14780 14350
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15028 13870 15056 14350
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14476 13530 14504 13806
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14476 13258 14504 13466
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14476 12850 14504 13194
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14752 12782 14780 13262
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13556 10674 13584 11222
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12898 9208 12954 9217
rect 12898 9143 12954 9152
rect 12912 9110 12940 9143
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12806 8528 12862 8537
rect 12716 8492 12768 8498
rect 12806 8463 12862 8472
rect 12716 8434 12768 8440
rect 12360 8078 12480 8106
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12360 7750 12388 7958
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12452 7002 12480 8078
rect 12820 7206 12848 8463
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 8090 12940 8230
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12268 6458 12296 6598
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12360 6186 12388 6598
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12452 5896 12480 6258
rect 12636 5914 12664 7142
rect 13004 6866 13032 10406
rect 13266 10296 13322 10305
rect 13266 10231 13322 10240
rect 13176 10056 13228 10062
rect 13096 10016 13176 10044
rect 13096 9450 13124 10016
rect 13176 9998 13228 10004
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 9178 13124 9386
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13082 9072 13138 9081
rect 13082 9007 13084 9016
rect 13136 9007 13138 9016
rect 13084 8978 13136 8984
rect 13096 7478 13124 8978
rect 13280 8294 13308 10231
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 13464 7410 13492 8434
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12624 5908 12676 5914
rect 12452 5868 12572 5896
rect 12544 5778 12572 5868
rect 12624 5850 12676 5856
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5409 12388 5510
rect 12346 5400 12402 5409
rect 12452 5370 12480 5714
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12346 5335 12402 5344
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12544 5250 12572 5578
rect 12452 5222 12572 5250
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4622 12388 4966
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12176 4508 12296 4536
rect 12268 2990 12296 4508
rect 12452 3652 12480 5222
rect 12636 5148 12664 5238
rect 12544 5120 12664 5148
rect 12544 4622 12572 5120
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4865 12664 4966
rect 12622 4856 12678 4865
rect 12622 4791 12678 4800
rect 12624 4752 12676 4758
rect 12622 4720 12624 4729
rect 12676 4720 12678 4729
rect 12622 4655 12678 4664
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12728 4078 12756 6734
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12636 3924 12664 4014
rect 12636 3896 12756 3924
rect 12452 3624 12572 3652
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12256 2984 12308 2990
rect 12084 2910 12204 2938
rect 12256 2926 12308 2932
rect 12072 2848 12124 2854
rect 12070 2816 12072 2825
rect 12176 2836 12204 2910
rect 12124 2816 12126 2825
rect 12176 2808 12296 2836
rect 12070 2751 12126 2760
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 12268 480 12296 2808
rect 12452 2514 12480 3062
rect 12544 2582 12572 3624
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12728 480 12756 3896
rect 12820 2922 12848 6054
rect 13004 5352 13032 6802
rect 12912 5324 13032 5352
rect 12912 4146 12940 5324
rect 13096 5284 13124 7142
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13188 6361 13216 6938
rect 13174 6352 13230 6361
rect 13174 6287 13230 6296
rect 13004 5256 13124 5284
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3516 12940 4082
rect 13004 3738 13032 5256
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12992 3528 13044 3534
rect 12912 3488 12992 3516
rect 12992 3470 13044 3476
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 13096 2514 13124 4558
rect 13188 4146 13216 6287
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 4622 13308 6190
rect 13372 6186 13400 7346
rect 13450 7304 13506 7313
rect 13450 7239 13506 7248
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13372 5846 13400 6122
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13372 5302 13400 5782
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13464 5098 13492 7239
rect 13648 6798 13676 8230
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13636 5568 13688 5574
rect 13556 5528 13636 5556
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13556 4758 13584 5528
rect 13636 5510 13688 5516
rect 13634 5400 13690 5409
rect 13634 5335 13690 5344
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13280 4146 13308 4558
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 13188 3913 13216 3946
rect 13174 3904 13230 3913
rect 13174 3839 13230 3848
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 2854 13400 3334
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13360 2848 13412 2854
rect 13648 2802 13676 5335
rect 13740 4758 13768 11562
rect 14108 11354 14136 11834
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14568 11150 14596 11562
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14094 10976 14150 10985
rect 14094 10911 14150 10920
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13832 10266 13860 10678
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13924 10130 13952 10367
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13832 8838 13860 10066
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13924 8090 13952 9318
rect 14016 8362 14044 9386
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14016 7993 14044 8026
rect 14002 7984 14058 7993
rect 14002 7919 14058 7928
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14016 6798 14044 7210
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6458 14044 6734
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13910 5536 13966 5545
rect 13910 5471 13966 5480
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13924 3074 13952 5471
rect 14108 5234 14136 10911
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 8838 14412 10610
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14568 10062 14596 11086
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 10056 14608 10062
rect 14462 10024 14518 10033
rect 14556 9998 14608 10004
rect 14462 9959 14518 9968
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 7886 14320 8298
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14292 6254 14320 6666
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14004 5024 14056 5030
rect 14002 4992 14004 5001
rect 14056 4992 14058 5001
rect 14002 4927 14058 4936
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14108 4010 14136 4626
rect 14186 4040 14242 4049
rect 14096 4004 14148 4010
rect 14186 3975 14188 3984
rect 14096 3946 14148 3952
rect 14240 3975 14242 3984
rect 14188 3946 14240 3952
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3194 14044 3470
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 13924 3046 14044 3074
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13360 2790 13412 2796
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13188 480 13216 2790
rect 13556 2774 13676 2802
rect 13556 480 13584 2774
rect 13740 2650 13768 2858
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 14016 480 14044 3046
rect 14292 2582 14320 5714
rect 14384 5370 14412 6734
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 14384 1714 14412 3402
rect 14476 2990 14504 9959
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 8906 14596 9522
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14660 8634 14688 8910
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14844 8566 14872 8842
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 7954 15056 10610
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14936 7410 14964 7754
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15028 6730 15056 7686
rect 15120 7546 15148 13330
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 6798 15148 7482
rect 15212 6866 15240 14214
rect 15304 13530 15332 14418
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15580 13462 15608 14350
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 10742 15332 11630
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 9110 15332 10406
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 7954 15332 8910
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15396 7290 15424 13330
rect 15764 13326 15792 13670
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15488 11286 15516 12543
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15488 9518 15516 11222
rect 15580 11218 15608 12718
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11898 15700 12242
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15764 11393 15792 13262
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12442 15884 12582
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15750 11384 15806 11393
rect 15750 11319 15806 11328
rect 15856 11286 15884 11834
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15856 10146 15884 11222
rect 15948 10266 15976 12854
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16040 10470 16068 12786
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15660 10124 15712 10130
rect 15856 10118 16068 10146
rect 15660 10066 15712 10072
rect 15672 9654 15700 10066
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15764 9178 15792 9998
rect 15948 9178 15976 9998
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15842 8392 15898 8401
rect 15842 8327 15898 8336
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15304 7262 15424 7290
rect 15476 7268 15528 7274
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15200 6656 15252 6662
rect 15304 6633 15332 7262
rect 15476 7210 15528 7216
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 7002 15424 7142
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15200 6598 15252 6604
rect 15290 6624 15346 6633
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5234 15056 6394
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14568 4486 14596 4626
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 3652 14596 4422
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14568 3624 14780 3652
rect 14752 3466 14780 3624
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 3058 14780 3402
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15028 2258 15056 4762
rect 15120 3942 15148 6122
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3534 15148 3878
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15212 2514 15240 6598
rect 15290 6559 15346 6568
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 2802 15332 5510
rect 15396 2990 15424 6802
rect 15488 5234 15516 7210
rect 15764 7002 15792 7958
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15764 6780 15792 6938
rect 15672 6752 15792 6780
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15488 3058 15516 3538
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15304 2774 15424 2802
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14936 2230 15056 2258
rect 14384 1686 14504 1714
rect 14476 480 14504 1686
rect 14936 480 14964 2230
rect 15396 480 15424 2774
rect 15580 2582 15608 5714
rect 15672 4214 15700 6752
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5234 15792 5714
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15764 3602 15792 5170
rect 15856 5148 15884 8327
rect 15948 8022 15976 9114
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 16040 7834 16068 10118
rect 16132 9926 16160 14214
rect 16224 13870 16252 14758
rect 16408 14482 16436 14962
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16408 13734 16436 14418
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16592 13530 16620 14758
rect 17144 14618 17172 22320
rect 17866 16960 17922 16969
rect 17866 16895 17922 16904
rect 17880 16250 17908 16895
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 10674 16252 12582
rect 16316 12102 16344 13330
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16394 12880 16450 12889
rect 16394 12815 16396 12824
rect 16448 12815 16450 12824
rect 16396 12786 16448 12792
rect 16394 12744 16450 12753
rect 16394 12679 16450 12688
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11762 16344 12038
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16408 10742 16436 12679
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16304 9376 16356 9382
rect 16224 9324 16304 9330
rect 16224 9318 16356 9324
rect 16224 9302 16344 9318
rect 16224 8430 16252 9302
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16120 8288 16172 8294
rect 16118 8256 16120 8265
rect 16172 8256 16174 8265
rect 16118 8191 16174 8200
rect 15948 7806 16068 7834
rect 15948 5273 15976 7806
rect 15934 5264 15990 5273
rect 15934 5199 15990 5208
rect 15856 5120 15976 5148
rect 15948 4758 15976 5120
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15672 2650 15700 3538
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16132 2990 16160 3334
rect 16224 2990 16252 8366
rect 16316 7002 16344 9046
rect 16408 8498 16436 9522
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16500 8090 16528 12582
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16592 11082 16620 12174
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16684 10674 16712 13126
rect 16868 12986 16896 13738
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 11286 16896 12786
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16868 11150 16896 11222
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10266 16712 10610
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16776 9722 16804 11086
rect 16854 10160 16910 10169
rect 16854 10095 16910 10104
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16868 9058 16896 10095
rect 16960 9178 16988 11154
rect 17052 11014 17080 14282
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 13938 17172 14214
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 13462 17172 13874
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16868 9030 16988 9058
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16764 8016 16816 8022
rect 16670 7984 16726 7993
rect 16764 7958 16816 7964
rect 16670 7919 16726 7928
rect 16684 7342 16712 7919
rect 16776 7410 16804 7958
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16316 5681 16344 6938
rect 16776 6798 16804 7346
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16394 6216 16450 6225
rect 16394 6151 16396 6160
rect 16448 6151 16450 6160
rect 16396 6122 16448 6128
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16302 5672 16358 5681
rect 16302 5607 16358 5616
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16500 4690 16528 5306
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 4162 16528 4218
rect 16316 4134 16528 4162
rect 16316 3602 16344 4134
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16316 3194 16344 3538
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16408 2922 16436 3946
rect 16592 3738 16620 4626
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16684 2990 16712 3878
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16304 2848 16356 2854
rect 16776 2802 16804 5510
rect 16868 5234 16896 5782
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16960 4706 16988 9030
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 6322 17080 7686
rect 17144 6866 17172 10474
rect 17236 8401 17264 13738
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 12850 17448 13670
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17512 12714 17540 14962
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 12368 17552 12374
rect 17604 12322 17632 12582
rect 17552 12316 17632 12322
rect 17500 12310 17632 12316
rect 17512 12294 17632 12310
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17328 11762 17356 12106
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17420 9450 17448 12106
rect 17604 11801 17632 12294
rect 17972 12238 18000 22471
rect 19798 22128 19854 22137
rect 19798 22063 19854 22072
rect 19154 20632 19210 20641
rect 19154 20567 19210 20576
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 19168 19514 19196 20567
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 18432 18902 18460 19246
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 19430 18320 19486 18329
rect 19430 18255 19486 18264
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19154 15600 19210 15609
rect 19154 15535 19210 15544
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18616 13938 18644 14418
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18524 13326 18552 13398
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12442 18552 13262
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17590 11792 17646 11801
rect 17590 11727 17646 11736
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17512 8974 17540 9522
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17222 8392 17278 8401
rect 17222 8327 17278 8336
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17236 7546 17264 8230
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17328 7002 17356 8230
rect 17604 8129 17632 11494
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17696 10198 17724 11154
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17788 9654 17816 11154
rect 17880 11150 17908 12174
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11694 18000 12038
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 18524 11082 18552 11494
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 9722 18000 10406
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 18616 9518 18644 13738
rect 18708 11830 18736 14418
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18800 12986 18828 13806
rect 18892 13705 18920 14214
rect 18878 13696 18934 13705
rect 18878 13631 18934 13640
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18800 11354 18828 12582
rect 18984 12442 19012 12786
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18694 11248 18750 11257
rect 18694 11183 18750 11192
rect 18708 10441 18736 11183
rect 18892 11150 18920 12310
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11694 19104 12242
rect 19064 11688 19116 11694
rect 19062 11656 19064 11665
rect 19116 11656 19118 11665
rect 19062 11591 19118 11600
rect 19168 11234 19196 15535
rect 19352 14770 19380 15982
rect 19444 15042 19472 18255
rect 19628 15201 19656 18770
rect 19614 15192 19670 15201
rect 19614 15127 19670 15136
rect 19616 15088 19668 15094
rect 19614 15056 19616 15065
rect 19668 15056 19670 15065
rect 19444 15014 19564 15042
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19260 14742 19380 14770
rect 19260 14074 19288 14742
rect 19338 14648 19394 14657
rect 19338 14583 19340 14592
rect 19392 14583 19394 14592
rect 19340 14554 19392 14560
rect 19444 14550 19472 14894
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19536 13954 19564 15014
rect 19614 14991 19670 15000
rect 19720 14006 19748 19246
rect 19708 14000 19760 14006
rect 19352 12594 19380 13942
rect 19536 13926 19656 13954
rect 19708 13942 19760 13948
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 18984 11206 19196 11234
rect 19260 12566 19380 12594
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18694 10432 18750 10441
rect 18694 10367 18750 10376
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18800 9586 18828 9862
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18786 9480 18842 9489
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17696 8430 17724 8978
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17590 8120 17646 8129
rect 17590 8055 17646 8064
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17052 5846 17080 6258
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 17038 5672 17094 5681
rect 17038 5607 17094 5616
rect 16868 4690 16988 4706
rect 16856 4684 16988 4690
rect 16908 4678 16988 4684
rect 16856 4626 16908 4632
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16960 4146 16988 4558
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16304 2790 16356 2796
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 480 15884 2246
rect 16316 480 16344 2790
rect 16684 2774 16804 2802
rect 16684 480 16712 2774
rect 16868 2650 16896 3878
rect 16960 3602 16988 4082
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17052 2106 17080 5607
rect 17144 3924 17172 6802
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17236 4185 17264 6122
rect 17420 5914 17448 6190
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5166 17356 5714
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17222 4176 17278 4185
rect 17222 4111 17278 4120
rect 17236 4078 17264 4111
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17144 3896 17264 3924
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 17144 480 17172 3606
rect 17236 3505 17264 3896
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 17328 2292 17356 4422
rect 17420 4026 17448 4558
rect 17512 4486 17540 5510
rect 17500 4480 17552 4486
rect 17604 4468 17632 7414
rect 17696 5148 17724 8366
rect 17788 5370 17816 9454
rect 18786 9415 18842 9424
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18432 9178 18460 9318
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 8430 18000 8910
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18616 8514 18644 9318
rect 18524 8486 18644 8514
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17972 7954 18000 8366
rect 18524 8362 18552 8486
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7018 18000 7890
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 17880 7002 18000 7018
rect 17880 6996 18012 7002
rect 17880 6990 17960 6996
rect 17880 5778 17908 6990
rect 17960 6938 18012 6944
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17972 6186 18000 6802
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18524 5778 18552 7142
rect 18616 7002 18644 8298
rect 18708 8090 18736 8366
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7818 18736 8026
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7410 18736 7754
rect 18800 7585 18828 9415
rect 18984 8786 19012 11206
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10810 19104 11086
rect 19154 10840 19210 10849
rect 19064 10804 19116 10810
rect 19154 10775 19210 10784
rect 19064 10746 19116 10752
rect 19168 10674 19196 10775
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19260 10169 19288 12566
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19352 11694 19380 12378
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19430 11656 19486 11665
rect 19430 11591 19486 11600
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19246 10160 19302 10169
rect 19246 10095 19302 10104
rect 19154 9480 19210 9489
rect 19154 9415 19210 9424
rect 18892 8758 19012 8786
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18786 7168 18842 7177
rect 18708 7002 18736 7142
rect 18786 7103 18842 7112
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18708 5846 18736 6258
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 17958 5672 18014 5681
rect 17958 5607 18014 5616
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17696 5120 17816 5148
rect 17972 5137 18000 5607
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17788 4554 17816 5120
rect 17958 5128 18014 5137
rect 17958 5063 18014 5072
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17604 4440 17724 4468
rect 17500 4422 17552 4428
rect 17420 3998 17632 4026
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17498 3904 17554 3913
rect 17420 3058 17448 3878
rect 17498 3839 17554 3848
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17512 2514 17540 3839
rect 17604 2582 17632 3998
rect 17696 3534 17724 4440
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17592 2576 17644 2582
rect 17788 2553 17816 4490
rect 17592 2518 17644 2524
rect 17774 2544 17830 2553
rect 17500 2508 17552 2514
rect 17774 2479 17830 2488
rect 17500 2450 17552 2456
rect 17328 2264 17632 2292
rect 17604 480 17632 2264
rect 17880 2258 17908 4762
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17972 3738 18000 4694
rect 18420 4616 18472 4622
rect 18472 4576 18552 4604
rect 18420 4558 18472 4564
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18524 4282 18552 4576
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17972 3058 18000 3674
rect 18064 3380 18092 4150
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18432 3534 18460 4014
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18055 3352 18092 3380
rect 18055 3176 18083 3352
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18055 3148 18092 3176
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17972 2446 18000 2994
rect 18064 2582 18092 3148
rect 18524 2650 18552 3878
rect 18616 3738 18644 3878
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18052 2576 18104 2582
rect 18708 2530 18736 4966
rect 18800 3602 18828 7103
rect 18892 6730 18920 8758
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18984 6866 19012 8570
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7342 19104 7822
rect 19168 7449 19196 9415
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19154 7440 19210 7449
rect 19154 7375 19210 7384
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5302 18920 6054
rect 19076 5574 19104 6938
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19168 5370 19196 6394
rect 19260 6118 19288 8366
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19352 5930 19380 11494
rect 19444 10606 19472 11591
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19444 10198 19472 10542
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19444 9586 19472 10134
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8634 19472 8978
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19444 6798 19472 8570
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6322 19472 6734
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19536 6202 19564 13806
rect 19628 8906 19656 13926
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19720 8634 19748 13738
rect 19812 13530 19840 22063
rect 20350 21584 20406 21593
rect 20350 21519 20406 21528
rect 20074 21176 20130 21185
rect 20074 21111 20130 21120
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 14113 19932 15302
rect 19890 14104 19946 14113
rect 19890 14039 19946 14048
rect 19996 13546 20024 15506
rect 20088 15162 20116 21111
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20166 16552 20222 16561
rect 20166 16487 20222 16496
rect 20180 16250 20208 16487
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19800 13524 19852 13530
rect 19996 13518 20116 13546
rect 19800 13466 19852 13472
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19812 12646 19840 13262
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12850 19932 13126
rect 19996 12850 20024 13330
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19800 12640 19852 12646
rect 19798 12608 19800 12617
rect 19852 12608 19854 12617
rect 19798 12543 19854 12552
rect 19904 12374 19932 12786
rect 19892 12368 19944 12374
rect 19892 12310 19944 12316
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19996 11898 20024 12242
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11098 20116 13518
rect 20180 12889 20208 15982
rect 20272 12918 20300 17682
rect 20364 15162 20392 21519
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19514 20760 19751
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20810 19272 20866 19281
rect 20810 19207 20866 19216
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20732 18426 20760 18799
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 17814 20576 18158
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20442 17368 20498 17377
rect 20732 17338 20760 17847
rect 20442 17303 20498 17312
rect 20720 17332 20772 17338
rect 20456 16794 20484 17303
rect 20720 17274 20772 17280
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20442 16008 20498 16017
rect 20442 15943 20498 15952
rect 20456 15706 20484 15943
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20442 15192 20498 15201
rect 20352 15156 20404 15162
rect 20442 15127 20498 15136
rect 20352 15098 20404 15104
rect 20260 12912 20312 12918
rect 20166 12880 20222 12889
rect 20260 12854 20312 12860
rect 20166 12815 20222 12824
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19996 11070 20116 11098
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 9178 19840 10066
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19628 7857 19656 8502
rect 19812 8498 19840 9114
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19904 8378 19932 8978
rect 19996 8566 20024 11070
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 19812 8350 19932 8378
rect 19614 7848 19670 7857
rect 19614 7783 19670 7792
rect 19628 7342 19656 7783
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19628 6254 19656 6598
rect 19260 5902 19380 5930
rect 19444 6174 19564 6202
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 3738 18920 4966
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18800 2990 18828 3402
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18052 2518 18104 2524
rect 18524 2502 18736 2530
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17880 2230 18000 2258
rect 17972 1986 18000 2230
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1958 18092 1986
rect 18064 480 18092 1958
rect 18524 480 18552 2502
rect 18800 2446 18828 2926
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18616 1601 18644 2042
rect 18602 1592 18658 1601
rect 18602 1527 18658 1536
rect 18892 1057 18920 3674
rect 18984 3602 19012 4626
rect 19076 4282 19104 5170
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19168 4486 19196 5034
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18970 3360 19026 3369
rect 18970 3295 19026 3304
rect 18984 2961 19012 3295
rect 19076 3126 19104 4082
rect 19168 3369 19196 4422
rect 19260 4026 19288 5902
rect 19260 3998 19380 4026
rect 19444 4010 19472 6174
rect 19720 6118 19748 7686
rect 19812 6610 19840 8350
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 20088 8242 20116 10950
rect 20180 10266 20208 11154
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20272 10130 20300 12174
rect 20364 11354 20392 12582
rect 20456 11642 20484 15127
rect 20548 14414 20576 17070
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20640 14346 20668 16594
rect 20824 16250 20852 19207
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20824 13938 20852 15438
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20626 13288 20682 13297
rect 20626 13223 20682 13232
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20548 12442 20576 12650
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20456 11614 20576 11642
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20364 10470 20392 11086
rect 20456 10606 20484 11494
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20364 9518 20392 10406
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19904 6798 19932 7754
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19812 6582 19932 6610
rect 19904 6361 19932 6582
rect 19890 6352 19946 6361
rect 19800 6316 19852 6322
rect 19890 6287 19946 6296
rect 19800 6258 19852 6264
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19812 5642 19840 6258
rect 19904 5710 19932 6287
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19800 5636 19852 5642
rect 19800 5578 19852 5584
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19154 3360 19210 3369
rect 19154 3295 19210 3304
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18970 2952 19026 2961
rect 19260 2938 19288 3878
rect 19352 3534 19380 3998
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 18970 2887 19026 2896
rect 19076 2910 19288 2938
rect 18984 2650 19012 2887
rect 19076 2666 19104 2910
rect 18972 2644 19024 2650
rect 19076 2638 19196 2666
rect 18972 2586 19024 2592
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 18878 1048 18934 1057
rect 18878 983 18934 992
rect 18984 480 19012 2314
rect 19076 2009 19104 2518
rect 19168 2310 19196 2638
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19062 2000 19118 2009
rect 19062 1935 19118 1944
rect 19444 480 19472 3334
rect 19536 2582 19564 5102
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 19812 4826 19840 5034
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19812 4146 19840 4762
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19628 3194 19656 3878
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19996 2836 20024 8230
rect 20088 8214 20392 8242
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 20088 3738 20116 7890
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 3942 20208 7822
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19904 2808 20024 2836
rect 19904 2666 19932 2808
rect 19812 2638 19932 2666
rect 19524 2576 19576 2582
rect 19524 2518 19576 2524
rect 19812 480 19840 2638
rect 20272 480 20300 7142
rect 20364 2514 20392 8214
rect 20456 5794 20484 9386
rect 20548 6458 20576 11614
rect 20640 9994 20668 13223
rect 20812 12776 20864 12782
rect 20718 12744 20774 12753
rect 20812 12718 20864 12724
rect 20718 12679 20720 12688
rect 20772 12679 20774 12688
rect 20720 12650 20772 12656
rect 20824 12345 20852 12718
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 21008 11898 21036 20159
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20732 8265 20760 11630
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20732 7478 20760 8191
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20640 6730 20668 7346
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5914 20576 6054
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20456 5766 20576 5794
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4758 20484 4966
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20456 4146 20484 4694
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20456 3534 20484 4082
rect 20548 4010 20576 5766
rect 20640 5030 20668 6666
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20732 4321 20760 7278
rect 20824 5273 20852 8366
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 20810 5264 20866 5273
rect 20810 5199 20866 5208
rect 20718 4312 20774 4321
rect 20718 4247 20774 4256
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20628 3936 20680 3942
rect 20534 3904 20590 3913
rect 20628 3878 20680 3884
rect 20534 3839 20590 3848
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20442 3088 20498 3097
rect 20442 3023 20444 3032
rect 20496 3023 20498 3032
rect 20444 2994 20496 3000
rect 20548 2514 20576 3839
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 4986 232 5042 241
rect 4986 167 5042 176
rect 5078 0 5134 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 6826 0 6882 480
rect 7286 0 7342 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9586 0 9642 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13542 0 13598 480
rect 14002 0 14058 480
rect 14462 0 14518 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15842 0 15898 480
rect 16302 0 16358 480
rect 16670 0 16726 480
rect 17130 0 17186 480
rect 17590 0 17646 480
rect 18050 0 18106 480
rect 18510 0 18566 480
rect 18970 0 19026 480
rect 19430 0 19486 480
rect 19798 0 19854 480
rect 20258 0 20314 480
rect 20640 241 20668 3878
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20824 2922 20852 3606
rect 20812 2916 20864 2922
rect 20812 2858 20864 2864
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20732 480 20760 2246
rect 20824 649 20852 2858
rect 20810 640 20866 649
rect 20810 575 20866 584
rect 21192 480 21220 5306
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21652 480 21680 4626
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 480 22140 4422
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22572 480 22600 2926
rect 20626 232 20682 241
rect 20626 167 20682 176
rect 20718 0 20774 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22098 0 22154 480
rect 22558 0 22614 480
<< via2 >>
rect 2962 22480 3018 22536
rect 2502 22072 2558 22128
rect 2410 21120 2466 21176
rect 1950 19760 2006 19816
rect 1950 19216 2006 19272
rect 1950 18808 2006 18864
rect 1674 18264 1730 18320
rect 1950 17856 2006 17912
rect 1858 17312 1914 17368
rect 1950 16496 2006 16552
rect 1950 15952 2006 16008
rect 2778 20168 2834 20224
rect 2778 15544 2834 15600
rect 1950 15036 1952 15056
rect 1952 15036 2004 15056
rect 2004 15036 2006 15056
rect 1950 15000 2006 15036
rect 1674 14612 1730 14648
rect 1674 14592 1676 14612
rect 1676 14592 1728 14612
rect 1728 14592 1730 14612
rect 1582 14048 1638 14104
rect 17958 22480 18014 22536
rect 3422 21528 3478 21584
rect 3330 16904 3386 16960
rect 3882 20576 3938 20632
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 3146 12844 3202 12880
rect 3146 12824 3148 12844
rect 3148 12824 3200 12844
rect 3200 12824 3202 12844
rect 3514 13640 3570 13696
rect 3606 13232 3662 13288
rect 3606 12280 3662 12336
rect 2870 3576 2926 3632
rect 2778 3440 2834 3496
rect 2778 2760 2834 2816
rect 2686 2488 2742 2544
rect 2226 1944 2282 2000
rect 3974 12688 4030 12744
rect 3974 11736 4030 11792
rect 3974 10784 4030 10840
rect 3974 10376 4030 10432
rect 4066 9968 4122 10024
rect 4066 9444 4122 9480
rect 4066 9424 4068 9444
rect 4068 9424 4120 9444
rect 4120 9424 4122 9444
rect 4066 8472 4122 8528
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4434 12844 4490 12880
rect 4434 12824 4436 12844
rect 4436 12824 4488 12844
rect 4488 12824 4490 12844
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4618 7828 4620 7848
rect 4620 7828 4672 7848
rect 4672 7828 4674 7848
rect 4066 7520 4122 7576
rect 4066 7112 4122 7168
rect 4618 7792 4674 7828
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 3974 4800 4030 4856
rect 4066 4256 4122 4312
rect 3422 2760 3478 2816
rect 3054 1536 3110 1592
rect 3606 584 3662 640
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 3882 992 3938 1048
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4802 8880 4858 8936
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 5538 8372 5540 8392
rect 5540 8372 5592 8392
rect 5592 8372 5594 8392
rect 5538 8336 5594 8372
rect 5630 7656 5686 7712
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 6090 9968 6146 10024
rect 5814 5752 5870 5808
rect 5814 4120 5870 4176
rect 5998 5208 6054 5264
rect 5814 3304 5870 3360
rect 5538 1944 5594 2000
rect 7194 13252 7250 13288
rect 7194 13232 7196 13252
rect 7196 13232 7248 13252
rect 7248 13232 7250 13252
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 6550 6568 6606 6624
rect 6458 3848 6514 3904
rect 6274 3440 6330 3496
rect 6274 2760 6330 2816
rect 6734 5772 6790 5808
rect 6734 5752 6736 5772
rect 6736 5752 6788 5772
rect 6788 5752 6790 5772
rect 6734 4664 6790 4720
rect 6642 3984 6698 4040
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7838 13232 7894 13288
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 9678 12688 9734 12744
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7378 10512 7434 10568
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7286 3168 7342 3224
rect 7838 8472 7894 8528
rect 9494 11192 9550 11248
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7654 7384 7710 7440
rect 8482 7656 8538 7712
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 9034 8880 9090 8936
rect 8666 7792 8722 7848
rect 8850 7792 8906 7848
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8482 6704 8538 6760
rect 8850 6160 8906 6216
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 8390 4936 8446 4992
rect 7930 3984 7986 4040
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8666 3848 8722 3904
rect 8206 2352 8262 2408
rect 8574 2896 8630 2952
rect 9034 5072 9090 5128
rect 9034 4664 9090 4720
rect 8942 3576 8998 3632
rect 8942 3168 8998 3224
rect 8758 2760 8814 2816
rect 10322 10412 10324 10432
rect 10324 10412 10376 10432
rect 10376 10412 10378 10432
rect 10322 10376 10378 10412
rect 10046 10240 10102 10296
rect 9770 9152 9826 9208
rect 9586 9016 9642 9072
rect 9678 8900 9734 8936
rect 9678 8880 9680 8900
rect 9680 8880 9732 8900
rect 9732 8880 9734 8900
rect 9770 8472 9826 8528
rect 9310 6604 9312 6624
rect 9312 6604 9364 6624
rect 9364 6604 9366 6624
rect 9310 6568 9366 6604
rect 9402 5772 9458 5808
rect 9402 5752 9404 5772
rect 9404 5752 9456 5772
rect 9456 5752 9458 5772
rect 10046 8064 10102 8120
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 10874 10104 10930 10160
rect 10690 9016 10746 9072
rect 10506 8336 10562 8392
rect 9862 6024 9918 6080
rect 9586 4936 9642 4992
rect 10138 5752 10194 5808
rect 10046 5616 10102 5672
rect 9954 4800 10010 4856
rect 10690 3168 10746 3224
rect 11058 8608 11114 8664
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11242 9460 11244 9480
rect 11244 9460 11296 9480
rect 11296 9460 11298 9480
rect 11242 9424 11298 9460
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11518 7148 11520 7168
rect 11520 7148 11572 7168
rect 11572 7148 11574 7168
rect 11518 7112 11574 7148
rect 11058 6840 11114 6896
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 10874 5616 10930 5672
rect 11058 5208 11114 5264
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11518 5208 11574 5264
rect 11058 3712 11114 3768
rect 11334 4700 11336 4720
rect 11336 4700 11388 4720
rect 11388 4700 11390 4720
rect 11334 4664 11390 4700
rect 12162 11328 12218 11384
rect 12162 11192 12218 11248
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 12806 11328 12862 11384
rect 12622 10532 12678 10568
rect 12622 10512 12624 10532
rect 12624 10512 12676 10532
rect 12676 10512 12678 10532
rect 11794 7928 11850 7984
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 10782 3032 10838 3088
rect 11058 3168 11114 3224
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 12162 8880 12218 8936
rect 11978 7112 12034 7168
rect 11978 6568 12034 6624
rect 12070 5480 12126 5536
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 12898 9152 12954 9208
rect 12806 8472 12862 8528
rect 13266 10240 13322 10296
rect 13082 9036 13138 9072
rect 13082 9016 13084 9036
rect 13084 9016 13136 9036
rect 13136 9016 13138 9036
rect 12346 5344 12402 5400
rect 12622 4800 12678 4856
rect 12622 4700 12624 4720
rect 12624 4700 12676 4720
rect 12676 4700 12678 4720
rect 12622 4664 12678 4700
rect 12070 2796 12072 2816
rect 12072 2796 12124 2816
rect 12124 2796 12126 2816
rect 12070 2760 12126 2796
rect 13174 6296 13230 6352
rect 13450 7248 13506 7304
rect 13634 5344 13690 5400
rect 13174 3848 13230 3904
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14094 10920 14150 10976
rect 13910 10376 13966 10432
rect 14002 7928 14058 7984
rect 13910 5480 13966 5536
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14462 9968 14518 10024
rect 14002 4972 14004 4992
rect 14004 4972 14056 4992
rect 14056 4972 14058 4992
rect 14002 4936 14058 4972
rect 14186 4004 14242 4040
rect 14186 3984 14188 4004
rect 14188 3984 14240 4004
rect 14240 3984 14242 4004
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 15474 12552 15530 12608
rect 15750 11328 15806 11384
rect 15842 8336 15898 8392
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15290 6568 15346 6624
rect 17866 16904 17922 16960
rect 16394 12844 16450 12880
rect 16394 12824 16396 12844
rect 16396 12824 16448 12844
rect 16448 12824 16450 12844
rect 16394 12688 16450 12744
rect 16118 8236 16120 8256
rect 16120 8236 16172 8256
rect 16172 8236 16174 8256
rect 16118 8200 16174 8236
rect 15934 5208 15990 5264
rect 16854 10104 16910 10160
rect 16670 7928 16726 7984
rect 16394 6180 16450 6216
rect 16394 6160 16396 6180
rect 16396 6160 16448 6180
rect 16448 6160 16450 6180
rect 16302 5616 16358 5672
rect 19798 22072 19854 22128
rect 19154 20576 19210 20632
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 19430 18264 19486 18320
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 19154 15544 19210 15600
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17590 11736 17646 11792
rect 17222 8336 17278 8392
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18878 13640 18934 13696
rect 18694 11192 18750 11248
rect 19062 11636 19064 11656
rect 19064 11636 19116 11656
rect 19116 11636 19118 11656
rect 19062 11600 19118 11636
rect 19614 15136 19670 15192
rect 19338 14612 19394 14648
rect 19338 14592 19340 14612
rect 19340 14592 19392 14612
rect 19392 14592 19394 14612
rect 19614 15036 19616 15056
rect 19616 15036 19668 15056
rect 19668 15036 19670 15056
rect 19614 15000 19670 15036
rect 18694 10376 18750 10432
rect 17590 8064 17646 8120
rect 17038 5616 17094 5672
rect 17222 4120 17278 4176
rect 17222 3440 17278 3496
rect 18786 9424 18842 9480
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 19154 10784 19210 10840
rect 19430 11600 19486 11656
rect 19246 10104 19302 10160
rect 19154 9424 19210 9480
rect 18786 7520 18842 7576
rect 18786 7112 18842 7168
rect 17958 5616 18014 5672
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 5072 18014 5128
rect 17498 3848 17554 3904
rect 17774 2488 17830 2544
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 19154 7384 19210 7440
rect 20350 21528 20406 21584
rect 20074 21120 20130 21176
rect 19890 14048 19946 14104
rect 20166 16496 20222 16552
rect 19798 12588 19800 12608
rect 19800 12588 19852 12608
rect 19852 12588 19854 12608
rect 19798 12552 19854 12588
rect 20994 20168 21050 20224
rect 20718 19760 20774 19816
rect 20810 19216 20866 19272
rect 20718 18808 20774 18864
rect 20718 17856 20774 17912
rect 20442 17312 20498 17368
rect 20442 15952 20498 16008
rect 20442 15136 20498 15192
rect 20166 12824 20222 12880
rect 19614 7792 19670 7848
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18602 1536 18658 1592
rect 18970 3304 19026 3360
rect 20626 13232 20682 13288
rect 19890 6296 19946 6352
rect 19154 3304 19210 3360
rect 18970 2896 19026 2952
rect 18878 992 18934 1048
rect 19062 1944 19118 2000
rect 20718 12708 20774 12744
rect 20718 12688 20720 12708
rect 20720 12688 20772 12708
rect 20772 12688 20774 12708
rect 20810 12280 20866 12336
rect 20718 8200 20774 8256
rect 20810 5208 20866 5264
rect 20718 4256 20774 4312
rect 20534 3848 20590 3904
rect 20442 3052 20498 3088
rect 20442 3032 20444 3052
rect 20444 3032 20496 3052
rect 20496 3032 20498 3052
rect 4986 176 5042 232
rect 20810 584 20866 640
rect 20626 176 20682 232
<< metal3 >>
rect 0 22538 480 22568
rect 2957 22538 3023 22541
rect 0 22536 3023 22538
rect 0 22480 2962 22536
rect 3018 22480 3023 22536
rect 0 22478 3023 22480
rect 0 22448 480 22478
rect 2957 22475 3023 22478
rect 17953 22538 18019 22541
rect 22320 22538 22800 22568
rect 17953 22536 22800 22538
rect 17953 22480 17958 22536
rect 18014 22480 22800 22536
rect 17953 22478 22800 22480
rect 17953 22475 18019 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 2497 22130 2563 22133
rect 0 22128 2563 22130
rect 0 22072 2502 22128
rect 2558 22072 2563 22128
rect 0 22070 2563 22072
rect 0 22040 480 22070
rect 2497 22067 2563 22070
rect 19793 22130 19859 22133
rect 22320 22130 22800 22160
rect 19793 22128 22800 22130
rect 19793 22072 19798 22128
rect 19854 22072 22800 22128
rect 19793 22070 22800 22072
rect 19793 22067 19859 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 3417 21586 3483 21589
rect 0 21584 3483 21586
rect 0 21528 3422 21584
rect 3478 21528 3483 21584
rect 0 21526 3483 21528
rect 0 21496 480 21526
rect 3417 21523 3483 21526
rect 20345 21586 20411 21589
rect 22320 21586 22800 21616
rect 20345 21584 22800 21586
rect 20345 21528 20350 21584
rect 20406 21528 22800 21584
rect 20345 21526 22800 21528
rect 20345 21523 20411 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 2405 21178 2471 21181
rect 0 21176 2471 21178
rect 0 21120 2410 21176
rect 2466 21120 2471 21176
rect 0 21118 2471 21120
rect 0 21088 480 21118
rect 2405 21115 2471 21118
rect 20069 21178 20135 21181
rect 22320 21178 22800 21208
rect 20069 21176 22800 21178
rect 20069 21120 20074 21176
rect 20130 21120 22800 21176
rect 20069 21118 22800 21120
rect 20069 21115 20135 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 3877 20634 3943 20637
rect 0 20632 3943 20634
rect 0 20576 3882 20632
rect 3938 20576 3943 20632
rect 0 20574 3943 20576
rect 0 20544 480 20574
rect 3877 20571 3943 20574
rect 19149 20634 19215 20637
rect 22320 20634 22800 20664
rect 19149 20632 22800 20634
rect 19149 20576 19154 20632
rect 19210 20576 22800 20632
rect 19149 20574 22800 20576
rect 19149 20571 19215 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 480 20166
rect 2773 20163 2839 20166
rect 20989 20226 21055 20229
rect 22320 20226 22800 20256
rect 20989 20224 22800 20226
rect 20989 20168 20994 20224
rect 21050 20168 22800 20224
rect 20989 20166 22800 20168
rect 20989 20163 21055 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 480 19214
rect 1945 19211 2011 19214
rect 20805 19274 20871 19277
rect 22320 19274 22800 19304
rect 20805 19272 22800 19274
rect 20805 19216 20810 19272
rect 20866 19216 22800 19272
rect 20805 19214 22800 19216
rect 20805 19211 20871 19214
rect 22320 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 20713 18866 20779 18869
rect 22320 18866 22800 18896
rect 20713 18864 22800 18866
rect 20713 18808 20718 18864
rect 20774 18808 22800 18864
rect 20713 18806 22800 18808
rect 20713 18803 20779 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 0 18232 480 18262
rect 1669 18259 1735 18262
rect 19425 18322 19491 18325
rect 22320 18322 22800 18352
rect 19425 18320 22800 18322
rect 19425 18264 19430 18320
rect 19486 18264 22800 18320
rect 19425 18262 22800 18264
rect 19425 18259 19491 18262
rect 22320 18232 22800 18262
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 480 17854
rect 1945 17851 2011 17854
rect 20713 17914 20779 17917
rect 22320 17914 22800 17944
rect 20713 17912 22800 17914
rect 20713 17856 20718 17912
rect 20774 17856 22800 17912
rect 20713 17854 22800 17856
rect 20713 17851 20779 17854
rect 22320 17824 22800 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1853 17370 1919 17373
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 480 17310
rect 1853 17307 1919 17310
rect 20437 17370 20503 17373
rect 22320 17370 22800 17400
rect 20437 17368 22800 17370
rect 20437 17312 20442 17368
rect 20498 17312 22800 17368
rect 20437 17310 22800 17312
rect 20437 17307 20503 17310
rect 22320 17280 22800 17310
rect 0 16962 480 16992
rect 3325 16962 3391 16965
rect 0 16960 3391 16962
rect 0 16904 3330 16960
rect 3386 16904 3391 16960
rect 0 16902 3391 16904
rect 0 16872 480 16902
rect 3325 16899 3391 16902
rect 17861 16962 17927 16965
rect 22320 16962 22800 16992
rect 17861 16960 22800 16962
rect 17861 16904 17866 16960
rect 17922 16904 22800 16960
rect 17861 16902 22800 16904
rect 17861 16899 17927 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 20161 16554 20227 16557
rect 22320 16554 22800 16584
rect 20161 16552 22800 16554
rect 20161 16496 20166 16552
rect 20222 16496 22800 16552
rect 20161 16494 22800 16496
rect 20161 16491 20227 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 20437 16010 20503 16013
rect 22320 16010 22800 16040
rect 20437 16008 22800 16010
rect 20437 15952 20442 16008
rect 20498 15952 22800 16008
rect 20437 15950 22800 15952
rect 20437 15947 20503 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 480 15542
rect 2773 15539 2839 15542
rect 19149 15602 19215 15605
rect 22320 15602 22800 15632
rect 19149 15600 22800 15602
rect 19149 15544 19154 15600
rect 19210 15544 22800 15600
rect 19149 15542 22800 15544
rect 19149 15539 19215 15542
rect 22320 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 19609 15194 19675 15197
rect 20437 15194 20503 15197
rect 19609 15192 20503 15194
rect 19609 15136 19614 15192
rect 19670 15136 20442 15192
rect 20498 15136 20503 15192
rect 19609 15134 20503 15136
rect 19609 15131 19675 15134
rect 20437 15131 20503 15134
rect 0 15058 480 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 480 14998
rect 1945 14995 2011 14998
rect 19609 15058 19675 15061
rect 22320 15058 22800 15088
rect 19609 15056 22800 15058
rect 19609 15000 19614 15056
rect 19670 15000 22800 15056
rect 19609 14998 22800 15000
rect 19609 14995 19675 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 19333 14650 19399 14653
rect 22320 14650 22800 14680
rect 19333 14648 22800 14650
rect 19333 14592 19338 14648
rect 19394 14592 22800 14648
rect 19333 14590 22800 14592
rect 19333 14587 19399 14590
rect 22320 14560 22800 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 480 14046
rect 1577 14043 1643 14046
rect 19885 14106 19951 14109
rect 22320 14106 22800 14136
rect 19885 14104 22800 14106
rect 19885 14048 19890 14104
rect 19946 14048 22800 14104
rect 19885 14046 22800 14048
rect 19885 14043 19951 14046
rect 22320 14016 22800 14046
rect 0 13698 480 13728
rect 3509 13698 3575 13701
rect 0 13696 3575 13698
rect 0 13640 3514 13696
rect 3570 13640 3575 13696
rect 0 13638 3575 13640
rect 0 13608 480 13638
rect 3509 13635 3575 13638
rect 18873 13698 18939 13701
rect 22320 13698 22800 13728
rect 18873 13696 22800 13698
rect 18873 13640 18878 13696
rect 18934 13640 22800 13696
rect 18873 13638 22800 13640
rect 18873 13635 18939 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 3601 13290 3667 13293
rect 0 13288 3667 13290
rect 0 13232 3606 13288
rect 3662 13232 3667 13288
rect 0 13230 3667 13232
rect 0 13200 480 13230
rect 3601 13227 3667 13230
rect 7189 13290 7255 13293
rect 7833 13290 7899 13293
rect 7189 13288 7899 13290
rect 7189 13232 7194 13288
rect 7250 13232 7838 13288
rect 7894 13232 7899 13288
rect 7189 13230 7899 13232
rect 7189 13227 7255 13230
rect 7833 13227 7899 13230
rect 20621 13290 20687 13293
rect 22320 13290 22800 13320
rect 20621 13288 22800 13290
rect 20621 13232 20626 13288
rect 20682 13232 22800 13288
rect 20621 13230 22800 13232
rect 20621 13227 20687 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 3141 12882 3207 12885
rect 4429 12882 4495 12885
rect 3141 12880 4495 12882
rect 3141 12824 3146 12880
rect 3202 12824 4434 12880
rect 4490 12824 4495 12880
rect 3141 12822 4495 12824
rect 3141 12819 3207 12822
rect 4429 12819 4495 12822
rect 16389 12882 16455 12885
rect 20161 12882 20227 12885
rect 16389 12880 20227 12882
rect 16389 12824 16394 12880
rect 16450 12824 20166 12880
rect 20222 12824 20227 12880
rect 16389 12822 20227 12824
rect 16389 12819 16455 12822
rect 20161 12819 20227 12822
rect 0 12746 480 12776
rect 3969 12746 4035 12749
rect 0 12744 4035 12746
rect 0 12688 3974 12744
rect 4030 12688 4035 12744
rect 0 12686 4035 12688
rect 0 12656 480 12686
rect 3969 12683 4035 12686
rect 9673 12746 9739 12749
rect 16389 12746 16455 12749
rect 9673 12744 16455 12746
rect 9673 12688 9678 12744
rect 9734 12688 16394 12744
rect 16450 12688 16455 12744
rect 9673 12686 16455 12688
rect 9673 12683 9739 12686
rect 16389 12683 16455 12686
rect 20713 12746 20779 12749
rect 22320 12746 22800 12776
rect 20713 12744 22800 12746
rect 20713 12688 20718 12744
rect 20774 12688 22800 12744
rect 20713 12686 22800 12688
rect 20713 12683 20779 12686
rect 22320 12656 22800 12686
rect 15469 12610 15535 12613
rect 19793 12610 19859 12613
rect 15469 12608 19859 12610
rect 15469 12552 15474 12608
rect 15530 12552 19798 12608
rect 19854 12552 19859 12608
rect 15469 12550 19859 12552
rect 15469 12547 15535 12550
rect 19793 12547 19859 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 3601 12338 3667 12341
rect 0 12336 3667 12338
rect 0 12280 3606 12336
rect 3662 12280 3667 12336
rect 0 12278 3667 12280
rect 0 12248 480 12278
rect 3601 12275 3667 12278
rect 20805 12338 20871 12341
rect 22320 12338 22800 12368
rect 20805 12336 22800 12338
rect 20805 12280 20810 12336
rect 20866 12280 22800 12336
rect 20805 12278 22800 12280
rect 20805 12275 20871 12278
rect 22320 12248 22800 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 3969 11794 4035 11797
rect 0 11792 4035 11794
rect 0 11736 3974 11792
rect 4030 11736 4035 11792
rect 0 11734 4035 11736
rect 0 11704 480 11734
rect 3969 11731 4035 11734
rect 17585 11794 17651 11797
rect 22320 11794 22800 11824
rect 17585 11792 22800 11794
rect 17585 11736 17590 11792
rect 17646 11736 22800 11792
rect 17585 11734 22800 11736
rect 17585 11731 17651 11734
rect 22320 11704 22800 11734
rect 19057 11658 19123 11661
rect 19425 11658 19491 11661
rect 19057 11656 19491 11658
rect 19057 11600 19062 11656
rect 19118 11600 19430 11656
rect 19486 11600 19491 11656
rect 19057 11598 19491 11600
rect 19057 11595 19123 11598
rect 19425 11595 19491 11598
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 12157 11386 12223 11389
rect 12801 11386 12867 11389
rect 0 11326 4906 11386
rect 0 11296 480 11326
rect 4846 11250 4906 11326
rect 12157 11384 12867 11386
rect 12157 11328 12162 11384
rect 12218 11328 12806 11384
rect 12862 11328 12867 11384
rect 12157 11326 12867 11328
rect 12157 11323 12223 11326
rect 12801 11323 12867 11326
rect 15745 11386 15811 11389
rect 22320 11386 22800 11416
rect 15745 11384 22800 11386
rect 15745 11328 15750 11384
rect 15806 11328 22800 11384
rect 15745 11326 22800 11328
rect 15745 11323 15811 11326
rect 22320 11296 22800 11326
rect 9489 11250 9555 11253
rect 4846 11248 9555 11250
rect 4846 11192 9494 11248
rect 9550 11192 9555 11248
rect 4846 11190 9555 11192
rect 9489 11187 9555 11190
rect 12157 11250 12223 11253
rect 18689 11250 18755 11253
rect 12157 11248 18755 11250
rect 12157 11192 12162 11248
rect 12218 11192 18694 11248
rect 18750 11192 18755 11248
rect 12157 11190 18755 11192
rect 12157 11187 12223 11190
rect 14046 10981 14106 11190
rect 18689 11187 18755 11190
rect 14046 10976 14155 10981
rect 14046 10920 14094 10976
rect 14150 10920 14155 10976
rect 14046 10918 14155 10920
rect 14089 10915 14155 10918
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3969 10842 4035 10845
rect 0 10840 4035 10842
rect 0 10784 3974 10840
rect 4030 10784 4035 10840
rect 0 10782 4035 10784
rect 0 10752 480 10782
rect 3969 10779 4035 10782
rect 19149 10842 19215 10845
rect 22320 10842 22800 10872
rect 19149 10840 22800 10842
rect 19149 10784 19154 10840
rect 19210 10784 22800 10840
rect 19149 10782 22800 10784
rect 19149 10779 19215 10782
rect 22320 10752 22800 10782
rect 7373 10570 7439 10573
rect 12617 10570 12683 10573
rect 7373 10568 12683 10570
rect 7373 10512 7378 10568
rect 7434 10512 12622 10568
rect 12678 10512 12683 10568
rect 7373 10510 12683 10512
rect 7373 10507 7439 10510
rect 12617 10507 12683 10510
rect 0 10434 480 10464
rect 3969 10434 4035 10437
rect 0 10432 4035 10434
rect 0 10376 3974 10432
rect 4030 10376 4035 10432
rect 0 10374 4035 10376
rect 0 10344 480 10374
rect 3969 10371 4035 10374
rect 10317 10434 10383 10437
rect 13905 10434 13971 10437
rect 10317 10432 13971 10434
rect 10317 10376 10322 10432
rect 10378 10376 13910 10432
rect 13966 10376 13971 10432
rect 10317 10374 13971 10376
rect 10317 10371 10383 10374
rect 13905 10371 13971 10374
rect 18689 10434 18755 10437
rect 22320 10434 22800 10464
rect 18689 10432 22800 10434
rect 18689 10376 18694 10432
rect 18750 10376 22800 10432
rect 18689 10374 22800 10376
rect 18689 10371 18755 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 10041 10298 10107 10301
rect 13261 10298 13327 10301
rect 10041 10296 13327 10298
rect 10041 10240 10046 10296
rect 10102 10240 13266 10296
rect 13322 10240 13327 10296
rect 10041 10238 13327 10240
rect 10041 10235 10107 10238
rect 13261 10235 13327 10238
rect 10869 10162 10935 10165
rect 16849 10162 16915 10165
rect 19241 10162 19307 10165
rect 10869 10160 19307 10162
rect 10869 10104 10874 10160
rect 10930 10104 16854 10160
rect 16910 10104 19246 10160
rect 19302 10104 19307 10160
rect 10869 10102 19307 10104
rect 10869 10099 10935 10102
rect 16849 10099 16915 10102
rect 19241 10099 19307 10102
rect 0 10026 480 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 480 9966
rect 4061 9963 4127 9966
rect 6085 10026 6151 10029
rect 14457 10026 14523 10029
rect 22320 10026 22800 10056
rect 6085 10024 22800 10026
rect 6085 9968 6090 10024
rect 6146 9968 14462 10024
rect 14518 9968 22800 10024
rect 6085 9966 22800 9968
rect 6085 9963 6151 9966
rect 14457 9963 14523 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 0 9482 480 9512
rect 4061 9482 4127 9485
rect 0 9480 4127 9482
rect 0 9424 4066 9480
rect 4122 9424 4127 9480
rect 0 9422 4127 9424
rect 0 9392 480 9422
rect 4061 9419 4127 9422
rect 11237 9482 11303 9485
rect 18781 9482 18847 9485
rect 11237 9480 18847 9482
rect 11237 9424 11242 9480
rect 11298 9424 18786 9480
rect 18842 9424 18847 9480
rect 11237 9422 18847 9424
rect 11237 9419 11303 9422
rect 18781 9419 18847 9422
rect 19149 9482 19215 9485
rect 22320 9482 22800 9512
rect 19149 9480 22800 9482
rect 19149 9424 19154 9480
rect 19210 9424 22800 9480
rect 19149 9422 22800 9424
rect 19149 9419 19215 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 9765 9210 9831 9213
rect 12893 9210 12959 9213
rect 9765 9208 12959 9210
rect 9765 9152 9770 9208
rect 9826 9152 12898 9208
rect 12954 9152 12959 9208
rect 9765 9150 12959 9152
rect 9765 9147 9831 9150
rect 12893 9147 12959 9150
rect 0 9074 480 9104
rect 9581 9074 9647 9077
rect 0 9072 9647 9074
rect 0 9016 9586 9072
rect 9642 9016 9647 9072
rect 0 9014 9647 9016
rect 0 8984 480 9014
rect 9581 9011 9647 9014
rect 10685 9074 10751 9077
rect 13077 9074 13143 9077
rect 10685 9072 13143 9074
rect 10685 9016 10690 9072
rect 10746 9016 13082 9072
rect 13138 9016 13143 9072
rect 10685 9014 13143 9016
rect 10685 9011 10751 9014
rect 13077 9011 13143 9014
rect 19190 9012 19196 9076
rect 19260 9074 19266 9076
rect 22320 9074 22800 9104
rect 19260 9014 22800 9074
rect 19260 9012 19266 9014
rect 22320 8984 22800 9014
rect 4797 8938 4863 8941
rect 9029 8938 9095 8941
rect 4797 8936 9095 8938
rect 4797 8880 4802 8936
rect 4858 8880 9034 8936
rect 9090 8880 9095 8936
rect 4797 8878 9095 8880
rect 4797 8875 4863 8878
rect 9029 8875 9095 8878
rect 9673 8938 9739 8941
rect 12157 8938 12223 8941
rect 9673 8936 12223 8938
rect 9673 8880 9678 8936
rect 9734 8880 12162 8936
rect 12218 8880 12223 8936
rect 9673 8878 12223 8880
rect 9673 8875 9739 8878
rect 12157 8875 12223 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 10910 8604 10916 8668
rect 10980 8666 10986 8668
rect 11053 8666 11119 8669
rect 10980 8664 11119 8666
rect 10980 8608 11058 8664
rect 11114 8608 11119 8664
rect 10980 8606 11119 8608
rect 10980 8604 10986 8606
rect 11053 8603 11119 8606
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 7833 8530 7899 8533
rect 9765 8530 9831 8533
rect 7833 8528 9831 8530
rect 7833 8472 7838 8528
rect 7894 8472 9770 8528
rect 9826 8472 9831 8528
rect 7833 8470 9831 8472
rect 7833 8467 7899 8470
rect 9765 8467 9831 8470
rect 12801 8530 12867 8533
rect 22320 8530 22800 8560
rect 12801 8528 22800 8530
rect 12801 8472 12806 8528
rect 12862 8472 22800 8528
rect 12801 8470 22800 8472
rect 12801 8467 12867 8470
rect 22320 8440 22800 8470
rect 5533 8394 5599 8397
rect 10501 8394 10567 8397
rect 5533 8392 10567 8394
rect 5533 8336 5538 8392
rect 5594 8336 10506 8392
rect 10562 8336 10567 8392
rect 5533 8334 10567 8336
rect 5533 8331 5599 8334
rect 10501 8331 10567 8334
rect 15837 8394 15903 8397
rect 17217 8394 17283 8397
rect 15837 8392 17283 8394
rect 15837 8336 15842 8392
rect 15898 8336 17222 8392
rect 17278 8336 17283 8392
rect 15837 8334 17283 8336
rect 15837 8331 15903 8334
rect 17217 8331 17283 8334
rect 16113 8258 16179 8261
rect 20713 8258 20779 8261
rect 16113 8256 20779 8258
rect 16113 8200 16118 8256
rect 16174 8200 20718 8256
rect 20774 8200 20779 8256
rect 16113 8198 20779 8200
rect 16113 8195 16179 8198
rect 20713 8195 20779 8198
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 10041 8122 10107 8125
rect 17585 8122 17651 8125
rect 22320 8122 22800 8152
rect 0 8062 4906 8122
rect 0 8032 480 8062
rect 4846 7986 4906 8062
rect 10041 8120 14290 8122
rect 10041 8064 10046 8120
rect 10102 8064 14290 8120
rect 10041 8062 14290 8064
rect 10041 8059 10107 8062
rect 11789 7986 11855 7989
rect 13997 7986 14063 7989
rect 4846 7984 14063 7986
rect 4846 7928 11794 7984
rect 11850 7928 14002 7984
rect 14058 7928 14063 7984
rect 4846 7926 14063 7928
rect 14230 7986 14290 8062
rect 17585 8120 22800 8122
rect 17585 8064 17590 8120
rect 17646 8064 22800 8120
rect 17585 8062 22800 8064
rect 17585 8059 17651 8062
rect 22320 8032 22800 8062
rect 16665 7986 16731 7989
rect 14230 7984 16731 7986
rect 14230 7928 16670 7984
rect 16726 7928 16731 7984
rect 14230 7926 16731 7928
rect 11789 7923 11855 7926
rect 13997 7923 14063 7926
rect 16665 7923 16731 7926
rect 4613 7850 4679 7853
rect 8661 7850 8727 7853
rect 4613 7848 8727 7850
rect 4613 7792 4618 7848
rect 4674 7792 8666 7848
rect 8722 7792 8727 7848
rect 4613 7790 8727 7792
rect 4613 7787 4679 7790
rect 8661 7787 8727 7790
rect 8845 7850 8911 7853
rect 19609 7850 19675 7853
rect 8845 7848 19675 7850
rect 8845 7792 8850 7848
rect 8906 7792 19614 7848
rect 19670 7792 19675 7848
rect 8845 7790 19675 7792
rect 8845 7787 8911 7790
rect 19609 7787 19675 7790
rect 5625 7714 5691 7717
rect 8477 7714 8543 7717
rect 5625 7712 8543 7714
rect 5625 7656 5630 7712
rect 5686 7656 8482 7712
rect 8538 7656 8543 7712
rect 5625 7654 8543 7656
rect 5625 7651 5691 7654
rect 8477 7651 8543 7654
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 480 7518
rect 4061 7515 4127 7518
rect 18781 7578 18847 7581
rect 22320 7578 22800 7608
rect 18781 7576 22800 7578
rect 18781 7520 18786 7576
rect 18842 7520 22800 7576
rect 18781 7518 22800 7520
rect 18781 7515 18847 7518
rect 22320 7488 22800 7518
rect 7649 7442 7715 7445
rect 19149 7442 19215 7445
rect 7649 7440 19215 7442
rect 7649 7384 7654 7440
rect 7710 7384 19154 7440
rect 19210 7384 19215 7440
rect 7649 7382 19215 7384
rect 7649 7379 7715 7382
rect 13494 7309 13554 7382
rect 19149 7379 19215 7382
rect 13445 7304 13554 7309
rect 13445 7248 13450 7304
rect 13506 7248 13554 7304
rect 13445 7246 13554 7248
rect 14414 7246 18706 7306
rect 13445 7243 13511 7246
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 10910 7108 10916 7172
rect 10980 7170 10986 7172
rect 11513 7170 11579 7173
rect 10980 7168 11579 7170
rect 10980 7112 11518 7168
rect 11574 7112 11579 7168
rect 10980 7110 11579 7112
rect 10980 7108 10986 7110
rect 11513 7107 11579 7110
rect 11973 7170 12039 7173
rect 14414 7170 14474 7246
rect 11973 7168 14474 7170
rect 11973 7112 11978 7168
rect 12034 7112 14474 7168
rect 11973 7110 14474 7112
rect 11973 7107 12039 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 11053 6898 11119 6901
rect 4846 6896 11119 6898
rect 4846 6840 11058 6896
rect 11114 6840 11119 6896
rect 4846 6838 11119 6840
rect 0 6762 480 6792
rect 4846 6762 4906 6838
rect 11053 6835 11119 6838
rect 0 6702 4906 6762
rect 0 6672 480 6702
rect 8334 6700 8340 6764
rect 8404 6762 8410 6764
rect 8477 6762 8543 6765
rect 8404 6760 8543 6762
rect 8404 6704 8482 6760
rect 8538 6704 8543 6760
rect 8404 6702 8543 6704
rect 18646 6762 18706 7246
rect 18781 7170 18847 7173
rect 22320 7170 22800 7200
rect 18781 7168 22800 7170
rect 18781 7112 18786 7168
rect 18842 7112 22800 7168
rect 18781 7110 22800 7112
rect 18781 7107 18847 7110
rect 22320 7080 22800 7110
rect 22320 6762 22800 6792
rect 18646 6702 22800 6762
rect 8404 6700 8410 6702
rect 8477 6699 8543 6702
rect 22320 6672 22800 6702
rect 6545 6626 6611 6629
rect 9305 6626 9371 6629
rect 6545 6624 9371 6626
rect 6545 6568 6550 6624
rect 6606 6568 9310 6624
rect 9366 6568 9371 6624
rect 6545 6566 9371 6568
rect 6545 6563 6611 6566
rect 9305 6563 9371 6566
rect 11973 6626 12039 6629
rect 15285 6626 15351 6629
rect 11973 6624 15351 6626
rect 11973 6568 11978 6624
rect 12034 6568 15290 6624
rect 15346 6568 15351 6624
rect 11973 6566 15351 6568
rect 11973 6563 12039 6566
rect 15285 6563 15351 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 13169 6354 13235 6357
rect 19885 6354 19951 6357
rect 13169 6352 19951 6354
rect 13169 6296 13174 6352
rect 13230 6296 19890 6352
rect 19946 6296 19951 6352
rect 13169 6294 19951 6296
rect 13169 6291 13235 6294
rect 19885 6291 19951 6294
rect 0 6218 480 6248
rect 8845 6218 8911 6221
rect 16389 6218 16455 6221
rect 22320 6218 22800 6248
rect 0 6216 8911 6218
rect 0 6160 8850 6216
rect 8906 6160 8911 6216
rect 0 6158 8911 6160
rect 0 6128 480 6158
rect 8845 6155 8911 6158
rect 12390 6216 16455 6218
rect 12390 6160 16394 6216
rect 16450 6160 16455 6216
rect 12390 6158 16455 6160
rect 9857 6082 9923 6085
rect 12390 6082 12450 6158
rect 16389 6155 16455 6158
rect 18646 6158 22800 6218
rect 9857 6080 12450 6082
rect 9857 6024 9862 6080
rect 9918 6024 12450 6080
rect 9857 6022 12450 6024
rect 9857 6019 9923 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 5809 5810 5875 5813
rect 0 5808 5875 5810
rect 0 5752 5814 5808
rect 5870 5752 5875 5808
rect 0 5750 5875 5752
rect 0 5720 480 5750
rect 5809 5747 5875 5750
rect 6729 5810 6795 5813
rect 9397 5810 9463 5813
rect 6729 5808 9463 5810
rect 6729 5752 6734 5808
rect 6790 5752 9402 5808
rect 9458 5752 9463 5808
rect 6729 5750 9463 5752
rect 6729 5747 6795 5750
rect 9397 5747 9463 5750
rect 10133 5810 10199 5813
rect 18646 5810 18706 6158
rect 22320 6128 22800 6158
rect 22320 5810 22800 5840
rect 10133 5808 18706 5810
rect 10133 5752 10138 5808
rect 10194 5752 18706 5808
rect 10133 5750 18706 5752
rect 18830 5750 22800 5810
rect 10133 5747 10199 5750
rect 10041 5676 10107 5677
rect 9990 5612 9996 5676
rect 10060 5674 10107 5676
rect 10869 5674 10935 5677
rect 10060 5672 10935 5674
rect 10102 5616 10874 5672
rect 10930 5616 10935 5672
rect 10060 5614 10935 5616
rect 10060 5612 10107 5614
rect 10041 5611 10107 5612
rect 10869 5611 10935 5614
rect 16297 5674 16363 5677
rect 17033 5674 17099 5677
rect 16297 5672 17099 5674
rect 16297 5616 16302 5672
rect 16358 5616 17038 5672
rect 17094 5616 17099 5672
rect 16297 5614 17099 5616
rect 16297 5611 16363 5614
rect 17033 5611 17099 5614
rect 17953 5674 18019 5677
rect 18830 5674 18890 5750
rect 22320 5720 22800 5750
rect 17953 5672 18890 5674
rect 17953 5616 17958 5672
rect 18014 5616 18890 5672
rect 17953 5614 18890 5616
rect 17953 5611 18019 5614
rect 12065 5538 12131 5541
rect 13905 5538 13971 5541
rect 12065 5536 13971 5538
rect 12065 5480 12070 5536
rect 12126 5480 13910 5536
rect 13966 5480 13971 5536
rect 12065 5478 13971 5480
rect 12065 5475 12131 5478
rect 13905 5475 13971 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 12341 5402 12407 5405
rect 13629 5402 13695 5405
rect 12341 5400 13695 5402
rect 12341 5344 12346 5400
rect 12402 5344 13634 5400
rect 13690 5344 13695 5400
rect 12341 5342 13695 5344
rect 12341 5339 12407 5342
rect 13629 5339 13695 5342
rect 0 5266 480 5296
rect 5993 5266 6059 5269
rect 0 5264 6059 5266
rect 0 5208 5998 5264
rect 6054 5208 6059 5264
rect 0 5206 6059 5208
rect 0 5176 480 5206
rect 5993 5203 6059 5206
rect 11053 5266 11119 5269
rect 11513 5266 11579 5269
rect 15929 5266 15995 5269
rect 11053 5264 15995 5266
rect 11053 5208 11058 5264
rect 11114 5208 11518 5264
rect 11574 5208 15934 5264
rect 15990 5208 15995 5264
rect 11053 5206 15995 5208
rect 11053 5203 11119 5206
rect 11513 5203 11579 5206
rect 15929 5203 15995 5206
rect 20805 5266 20871 5269
rect 22320 5266 22800 5296
rect 20805 5264 22800 5266
rect 20805 5208 20810 5264
rect 20866 5208 22800 5264
rect 20805 5206 22800 5208
rect 20805 5203 20871 5206
rect 22320 5176 22800 5206
rect 9029 5130 9095 5133
rect 17953 5130 18019 5133
rect 9029 5128 18019 5130
rect 9029 5072 9034 5128
rect 9090 5072 17958 5128
rect 18014 5072 18019 5128
rect 9029 5070 18019 5072
rect 9029 5067 9095 5070
rect 17953 5067 18019 5070
rect 8385 4994 8451 4997
rect 9581 4994 9647 4997
rect 13997 4994 14063 4997
rect 8385 4992 14063 4994
rect 8385 4936 8390 4992
rect 8446 4936 9586 4992
rect 9642 4936 14002 4992
rect 14058 4936 14063 4992
rect 8385 4934 14063 4936
rect 8385 4931 8451 4934
rect 9581 4931 9647 4934
rect 13997 4931 14063 4934
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 480 4798
rect 3969 4795 4035 4798
rect 9949 4858 10015 4861
rect 12617 4858 12683 4861
rect 22320 4858 22800 4888
rect 9949 4856 12683 4858
rect 9949 4800 9954 4856
rect 10010 4800 12622 4856
rect 12678 4800 12683 4856
rect 9949 4798 12683 4800
rect 9949 4795 10015 4798
rect 12617 4795 12683 4798
rect 15150 4798 22800 4858
rect 6729 4722 6795 4725
rect 9029 4722 9095 4725
rect 6729 4720 9095 4722
rect 6729 4664 6734 4720
rect 6790 4664 9034 4720
rect 9090 4664 9095 4720
rect 6729 4662 9095 4664
rect 6729 4659 6795 4662
rect 9029 4659 9095 4662
rect 9990 4660 9996 4724
rect 10060 4722 10066 4724
rect 11329 4722 11395 4725
rect 10060 4720 11395 4722
rect 10060 4664 11334 4720
rect 11390 4664 11395 4720
rect 10060 4662 11395 4664
rect 10060 4660 10066 4662
rect 11329 4659 11395 4662
rect 12617 4722 12683 4725
rect 15150 4722 15210 4798
rect 22320 4768 22800 4798
rect 12617 4720 15210 4722
rect 12617 4664 12622 4720
rect 12678 4664 15210 4720
rect 12617 4662 15210 4664
rect 12617 4659 12683 4662
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 20713 4314 20779 4317
rect 22320 4314 22800 4344
rect 20713 4312 22800 4314
rect 20713 4256 20718 4312
rect 20774 4256 22800 4312
rect 20713 4254 22800 4256
rect 20713 4251 20779 4254
rect 22320 4224 22800 4254
rect 5809 4178 5875 4181
rect 17217 4178 17283 4181
rect 5809 4176 17283 4178
rect 5809 4120 5814 4176
rect 5870 4120 17222 4176
rect 17278 4120 17283 4176
rect 5809 4118 17283 4120
rect 5809 4115 5875 4118
rect 6686 4045 6746 4118
rect 17217 4115 17283 4118
rect 6637 4040 6746 4045
rect 6637 3984 6642 4040
rect 6698 3984 6746 4040
rect 6637 3982 6746 3984
rect 7925 4042 7991 4045
rect 14181 4042 14247 4045
rect 7925 4040 14247 4042
rect 7925 3984 7930 4040
rect 7986 3984 14186 4040
rect 14242 3984 14247 4040
rect 7925 3982 14247 3984
rect 6637 3979 6703 3982
rect 7925 3979 7991 3982
rect 14181 3979 14247 3982
rect 0 3906 480 3936
rect 6453 3906 6519 3909
rect 0 3904 6519 3906
rect 0 3848 6458 3904
rect 6514 3848 6519 3904
rect 0 3846 6519 3848
rect 0 3816 480 3846
rect 6453 3843 6519 3846
rect 8661 3906 8727 3909
rect 13169 3906 13235 3909
rect 8661 3904 13235 3906
rect 8661 3848 8666 3904
rect 8722 3848 13174 3904
rect 13230 3848 13235 3904
rect 8661 3846 13235 3848
rect 8661 3843 8727 3846
rect 13169 3843 13235 3846
rect 17493 3906 17559 3909
rect 19190 3906 19196 3908
rect 17493 3904 19196 3906
rect 17493 3848 17498 3904
rect 17554 3848 19196 3904
rect 17493 3846 19196 3848
rect 17493 3843 17559 3846
rect 19190 3844 19196 3846
rect 19260 3844 19266 3908
rect 20529 3906 20595 3909
rect 22320 3906 22800 3936
rect 20529 3904 22800 3906
rect 20529 3848 20534 3904
rect 20590 3848 22800 3904
rect 20529 3846 22800 3848
rect 20529 3843 20595 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 11053 3770 11119 3773
rect 10918 3768 11119 3770
rect 10918 3712 11058 3768
rect 11114 3712 11119 3768
rect 10918 3710 11119 3712
rect 2865 3634 2931 3637
rect 8937 3634 9003 3637
rect 2865 3632 9003 3634
rect 2865 3576 2870 3632
rect 2926 3576 8942 3632
rect 8998 3576 9003 3632
rect 2865 3574 9003 3576
rect 2865 3571 2931 3574
rect 8937 3571 9003 3574
rect 0 3498 480 3528
rect 2773 3498 2839 3501
rect 0 3496 2839 3498
rect 0 3440 2778 3496
rect 2834 3440 2839 3496
rect 0 3438 2839 3440
rect 0 3408 480 3438
rect 2773 3435 2839 3438
rect 6269 3498 6335 3501
rect 10918 3498 10978 3710
rect 11053 3707 11119 3710
rect 6269 3496 10978 3498
rect 6269 3440 6274 3496
rect 6330 3440 10978 3496
rect 6269 3438 10978 3440
rect 17217 3498 17283 3501
rect 22320 3498 22800 3528
rect 17217 3496 22800 3498
rect 17217 3440 17222 3496
rect 17278 3440 22800 3496
rect 17217 3438 22800 3440
rect 6269 3435 6335 3438
rect 17217 3435 17283 3438
rect 22320 3408 22800 3438
rect 5809 3362 5875 3365
rect 9990 3362 9996 3364
rect 5809 3360 9996 3362
rect 5809 3304 5814 3360
rect 5870 3304 9996 3360
rect 5809 3302 9996 3304
rect 5809 3299 5875 3302
rect 9990 3300 9996 3302
rect 10060 3300 10066 3364
rect 18965 3362 19031 3365
rect 19149 3362 19215 3365
rect 18965 3360 19215 3362
rect 18965 3304 18970 3360
rect 19026 3304 19154 3360
rect 19210 3304 19215 3360
rect 18965 3302 19215 3304
rect 18965 3299 19031 3302
rect 19149 3299 19215 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 7281 3226 7347 3229
rect 8937 3226 9003 3229
rect 7281 3224 9003 3226
rect 7281 3168 7286 3224
rect 7342 3168 8942 3224
rect 8998 3168 9003 3224
rect 7281 3166 9003 3168
rect 7281 3163 7347 3166
rect 8937 3163 9003 3166
rect 10685 3226 10751 3229
rect 11053 3226 11119 3229
rect 10685 3224 11119 3226
rect 10685 3168 10690 3224
rect 10746 3168 11058 3224
rect 11114 3168 11119 3224
rect 10685 3166 11119 3168
rect 10685 3163 10751 3166
rect 11053 3163 11119 3166
rect 10777 3090 10843 3093
rect 20437 3090 20503 3093
rect 10777 3088 20503 3090
rect 10777 3032 10782 3088
rect 10838 3032 20442 3088
rect 20498 3032 20503 3088
rect 10777 3030 20503 3032
rect 10777 3027 10843 3030
rect 20437 3027 20503 3030
rect 0 2954 480 2984
rect 8569 2954 8635 2957
rect 10910 2954 10916 2956
rect 0 2894 674 2954
rect 0 2864 480 2894
rect 614 2818 674 2894
rect 8569 2952 10916 2954
rect 8569 2896 8574 2952
rect 8630 2896 10916 2952
rect 8569 2894 10916 2896
rect 8569 2891 8635 2894
rect 10910 2892 10916 2894
rect 10980 2892 10986 2956
rect 18965 2954 19031 2957
rect 22320 2954 22800 2984
rect 18965 2952 22800 2954
rect 18965 2896 18970 2952
rect 19026 2896 22800 2952
rect 18965 2894 22800 2896
rect 18965 2891 19031 2894
rect 22320 2864 22800 2894
rect 2773 2818 2839 2821
rect 614 2816 2839 2818
rect 614 2760 2778 2816
rect 2834 2760 2839 2816
rect 614 2758 2839 2760
rect 2773 2755 2839 2758
rect 3417 2818 3483 2821
rect 6269 2818 6335 2821
rect 3417 2816 6335 2818
rect 3417 2760 3422 2816
rect 3478 2760 6274 2816
rect 6330 2760 6335 2816
rect 3417 2758 6335 2760
rect 3417 2755 3483 2758
rect 6269 2755 6335 2758
rect 8753 2818 8819 2821
rect 12065 2818 12131 2821
rect 8753 2816 12131 2818
rect 8753 2760 8758 2816
rect 8814 2760 12070 2816
rect 12126 2760 12131 2816
rect 8753 2758 12131 2760
rect 8753 2755 8819 2758
rect 12065 2755 12131 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 2681 2546 2747 2549
rect 0 2544 2747 2546
rect 0 2488 2686 2544
rect 2742 2488 2747 2544
rect 0 2486 2747 2488
rect 0 2456 480 2486
rect 2681 2483 2747 2486
rect 17769 2546 17835 2549
rect 22320 2546 22800 2576
rect 17769 2544 22800 2546
rect 17769 2488 17774 2544
rect 17830 2488 22800 2544
rect 17769 2486 22800 2488
rect 17769 2483 17835 2486
rect 22320 2456 22800 2486
rect 8201 2410 8267 2413
rect 8334 2410 8340 2412
rect 8201 2408 8340 2410
rect 8201 2352 8206 2408
rect 8262 2352 8340 2408
rect 8201 2350 8340 2352
rect 8201 2347 8267 2350
rect 8334 2348 8340 2350
rect 8404 2348 8410 2412
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 2221 2002 2287 2005
rect 5533 2002 5599 2005
rect 0 2000 5599 2002
rect 0 1944 2226 2000
rect 2282 1944 5538 2000
rect 5594 1944 5599 2000
rect 0 1942 5599 1944
rect 0 1912 480 1942
rect 2221 1939 2287 1942
rect 5533 1939 5599 1942
rect 19057 2002 19123 2005
rect 22320 2002 22800 2032
rect 19057 2000 22800 2002
rect 19057 1944 19062 2000
rect 19118 1944 22800 2000
rect 19057 1942 22800 1944
rect 19057 1939 19123 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 3049 1594 3115 1597
rect 0 1592 3115 1594
rect 0 1536 3054 1592
rect 3110 1536 3115 1592
rect 0 1534 3115 1536
rect 0 1504 480 1534
rect 3049 1531 3115 1534
rect 18597 1594 18663 1597
rect 22320 1594 22800 1624
rect 18597 1592 22800 1594
rect 18597 1536 18602 1592
rect 18658 1536 22800 1592
rect 18597 1534 22800 1536
rect 18597 1531 18663 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 3877 1050 3943 1053
rect 0 1048 3943 1050
rect 0 992 3882 1048
rect 3938 992 3943 1048
rect 0 990 3943 992
rect 0 960 480 990
rect 3877 987 3943 990
rect 18873 1050 18939 1053
rect 22320 1050 22800 1080
rect 18873 1048 22800 1050
rect 18873 992 18878 1048
rect 18934 992 22800 1048
rect 18873 990 22800 992
rect 18873 987 18939 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 3601 642 3667 645
rect 0 640 3667 642
rect 0 584 3606 640
rect 3662 584 3667 640
rect 0 582 3667 584
rect 0 552 480 582
rect 3601 579 3667 582
rect 20805 642 20871 645
rect 22320 642 22800 672
rect 20805 640 22800 642
rect 20805 584 20810 640
rect 20866 584 22800 640
rect 20805 582 22800 584
rect 20805 579 20871 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 4981 234 5047 237
rect 0 232 5047 234
rect 0 176 4986 232
rect 5042 176 5047 232
rect 0 174 5047 176
rect 0 144 480 174
rect 4981 171 5047 174
rect 20621 234 20687 237
rect 22320 234 22800 264
rect 20621 232 22800 234
rect 20621 176 20626 232
rect 20682 176 22800 232
rect 20621 174 22800 176
rect 20621 171 20687 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 19196 9012 19260 9076
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 10916 8604 10980 8668
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 10916 7108 10980 7172
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 8340 6700 8404 6764
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 9996 5672 10060 5676
rect 9996 5616 10046 5672
rect 10046 5616 10060 5672
rect 9996 5612 10060 5616
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 9996 4660 10060 4724
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 19196 3844 19260 3908
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 9996 3300 10060 3364
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 10916 2892 10980 2956
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 8340 2348 8404 2412
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 10915 8668 10981 8669
rect 10915 8604 10916 8668
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 10918 7173 10978 8603
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 10915 7172 10981 7173
rect 10915 7108 10916 7172
rect 10980 7108 10981 7172
rect 10915 7107 10981 7108
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 8339 6764 8405 6765
rect 8339 6700 8340 6764
rect 8404 6700 8405 6764
rect 8339 6699 8405 6700
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 8342 2413 8402 6699
rect 9995 5676 10061 5677
rect 9995 5612 9996 5676
rect 10060 5612 10061 5676
rect 9995 5611 10061 5612
rect 9998 4725 10058 5611
rect 9995 4724 10061 4725
rect 9995 4660 9996 4724
rect 10060 4660 10061 4724
rect 9995 4659 10061 4660
rect 9998 3365 10058 4659
rect 9995 3364 10061 3365
rect 9995 3300 9996 3364
rect 10060 3300 10061 3364
rect 9995 3299 10061 3300
rect 10918 2957 10978 7107
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 10915 2956 10981 2957
rect 10915 2892 10916 2956
rect 10980 2892 10981 2956
rect 10915 2891 10981 2892
rect 8339 2412 8405 2413
rect 8339 2348 8340 2412
rect 8404 2348 8405 2412
rect 8339 2347 8405 2348
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 19195 9076 19261 9077
rect 19195 9012 19196 9076
rect 19260 9012 19261 9076
rect 19195 9011 19261 9012
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 19198 3909 19258 9011
rect 19195 3908 19261 3909
rect 19195 3844 19196 3908
rect 19260 3844 19261 3908
rect 19195 3843 19261 3844
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _032_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3496 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_24 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1606256979
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1606256979
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1606256979
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606256979
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _115_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6164 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76
timestamp 1606256979
transform 1 0 8096 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1606256979
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1606256979
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10580 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8924 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86
timestamp 1606256979
transform 1 0 9016 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1606256979
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100
timestamp 1606256979
transform 1 0 10304 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1606256979
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_115
timestamp 1606256979
transform 1 0 11684 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606256979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1606256979
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13156 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13064 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13800 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1606256979
transform 1 0 12972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_136
timestamp 1606256979
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1606256979
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp 1606256979
transform 1 0 13708 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_149
timestamp 1606256979
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1606256979
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606256979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15364 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1606256979
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1606256979
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16100 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 16192 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1606256979
transform 1 0 16652 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1606256979
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_167
timestamp 1606256979
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606256979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18584 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1606256979
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_200
timestamp 1606256979
transform 1 0 19504 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606256979
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_218
timestamp 1606256979
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1606256979
transform 1 0 4876 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 5244 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1606256979
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1606256979
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606256979
transform 1 0 9016 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10488 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1606256979
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606256979
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_99
timestamp 1606256979
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1606256979
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1606256979
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 13616 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp 1606256979
transform 1 0 13340 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1606256979
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606256979
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_163
timestamp 1606256979
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1606256979
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19780 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1606256979
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_199
timestamp 1606256979
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1606256979
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1606256979
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1748 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4508 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1606256979
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_34
timestamp 1606256979
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_46
timestamp 1606256979
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606256979
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606256979
transform 1 0 6992 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7544 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1606256979
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10304 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 1606256979
transform 1 0 11776 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13800 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_132
timestamp 1606256979
transform 1 0 13248 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_154
timestamp 1606256979
transform 1 0 15272 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18124 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 16836 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1606256979
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1606256979
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19136 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20240 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_194
timestamp 1606256979
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp 1606256979
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606256979
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2116 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4324 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1606256979
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1606256979
transform 1 0 6808 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8280 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_66
timestamp 1606256979
transform 1 0 7176 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_76
timestamp 1606256979
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606256979
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606256979
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11684 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1606256979
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp 1606256979
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606256979
transform 1 0 12696 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13248 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1606256979
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 15824 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16376 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1606256979
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606256979
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1606256979
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_164
timestamp 1606256979
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606256979
transform 1 0 17388 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1606256979
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1606256979
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606256979
transform 1 0 20240 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18400 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1606256979
transform 1 0 19872 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606256979
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2024 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1606256979
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1606256979
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_31
timestamp 1606256979
transform 1 0 3956 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1606256979
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_71
timestamp 1606256979
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1606256979
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_90
timestamp 1606256979
transform 1 0 9384 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1606256979
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1606256979
transform 1 0 11040 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1606256979
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1606256979
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1606256979
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12880 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_126
timestamp 1606256979
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_137
timestamp 1606256979
transform 1 0 13708 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606256979
transform 1 0 15272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15732 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1606256979
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1606256979
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1606256979
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606256979
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19596 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1606256979
transform 1 0 19228 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 1606256979
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1656 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1606256979
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4876 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3312 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1606256979
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1606256979
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_33
timestamp 1606256979
transform 1 0 4140 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_50
timestamp 1606256979
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1606256979
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1606256979
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6900 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8188 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1606256979
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_71
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9844 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606256979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_102
timestamp 1606256979
transform 1 0 10488 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1606256979
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1606256979
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1606256979
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606256979
transform 1 0 11040 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1606256979
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1606256979
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606256979
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606256979
transform 1 0 14260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14352 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1606256979
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16100 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_147
timestamp 1606256979
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1606256979
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1606256979
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 17756 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1606256979
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_171
timestamp 1606256979
transform 1 0 16836 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19412 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 20148 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19136 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1606256979
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1606256979
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp 1606256979
transform 1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1606256979
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_216
timestamp 1606256979
transform 1 0 20976 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606256979
transform 1 0 1656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_9
timestamp 1606256979
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4692 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1606256979
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1606256979
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_55
timestamp 1606256979
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8464 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1606256979
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1606256979
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1606256979
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11040 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_105
timestamp 1606256979
transform 1 0 10764 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1606256979
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 12696 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1606256979
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1606256979
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15640 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 18032 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1606256979
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 17664 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 1606256979
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1606256979
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1606256979
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19596 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 18584 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1606256979
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1606256979
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1606256979
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2116 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1606256979
transform 1 0 2944 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3404 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 1606256979
transform 1 0 3312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_34
timestamp 1606256979
transform 1 0 4232 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_40
timestamp 1606256979
transform 1 0 4784 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1606256979
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1606256979
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8556 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1606256979
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1606256979
transform 1 0 8096 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1606256979
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10212 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1606256979
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11224 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1606256979
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1606256979
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12696 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_135
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1606256979
transform 1 0 16192 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1606256979
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_158
timestamp 1606256979
transform 1 0 15640 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 18216 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1606256979
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606256979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1606256979
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 18676 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1606256979
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1606256979
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 20700 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1606256979
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp 1606256979
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606256979
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1606256979
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1606256979
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606256979
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5244 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1606256979
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1606256979
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1606256979
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7452 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1606256979
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_78
timestamp 1606256979
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1606256979
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12604 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_122
timestamp 1606256979
transform 1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1606256979
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1606256979
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15640 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1606256979
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17296 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_174
timestamp 1606256979
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1606256979
transform 1 0 18768 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_196
timestamp 1606256979
transform 1 0 19136 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1606256979
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1606256979
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1606256979
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_24
timestamp 1606256979
transform 1 0 3312 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1606256979
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606256979
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1606256979
transform 1 0 5888 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 8188 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_71
timestamp 1606256979
transform 1 0 7636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_96
timestamp 1606256979
transform 1 0 9936 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606256979
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13432 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15824 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_150
timestamp 1606256979
transform 1 0 14904 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1606256979
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 16836 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1606256979
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1606256979
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1606256979
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp 1606256979
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1606256979
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1606256979
transform 1 0 2024 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1606256979
transform 1 0 1932 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1606256979
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1606256979
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1606256979
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606256979
transform 1 0 5520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6164 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1606256979
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1606256979
transform 1 0 5796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7820 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1606256979
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_82
timestamp 1606256979
transform 1 0 8648 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10672 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12512 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1606256979
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1606256979
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_181
timestamp 1606256979
transform 1 0 17756 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_187
timestamp 1606256979
transform 1 0 18308 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 20240 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18400 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_204
timestamp 1606256979
transform 1 0 19872 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1606256979
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1606256979
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp 1606256979
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1606256979
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4784 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_28
timestamp 1606256979
transform 1 0 3680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1606256979
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6440 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_49
timestamp 1606256979
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1606256979
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1606256979
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 8096 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1606256979
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1606256979
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1606256979
transform 1 0 8372 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1606256979
transform 1 0 8740 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8832 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1606256979
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1606256979
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606256979
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1606256979
transform 1 0 11500 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1606256979
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1606256979
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1606256979
transform 1 0 13892 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 16192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1606256979
transform 1 0 15180 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1606256979
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1606256979
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606256979
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1606256979
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16928 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1606256979
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_171
timestamp 1606256979
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606256979
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_171
timestamp 1606256979
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19688 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18584 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1606256979
transform 1 0 18860 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1606256979
transform 1 0 19596 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1606256979
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1606256979
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1606256979
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606256979
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1606256979
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606256979
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606256979
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606256979
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606256979
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_78
timestamp 1606256979
transform 1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9016 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1606256979
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1606256979
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_106
timestamp 1606256979
transform 1 0 10856 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_110
timestamp 1606256979
transform 1 0 11224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1606256979
transform 1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 15272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1606256979
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1606256979
transform 1 0 15548 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1606256979
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1606256979
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18676 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_190
timestamp 1606256979
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1606256979
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1606256979
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1606256979
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4324 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_24
timestamp 1606256979
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606256979
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5980 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1606256979
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1606256979
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1606256979
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_102
timestamp 1606256979
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11500 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_110
timestamp 1606256979
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13340 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1606256979
transform 1 0 12972 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606256979
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1606256979
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_185
timestamp 1606256979
transform 1 0 18124 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1606256979
transform 1 0 19228 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606256979
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2852 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1606256979
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_17
timestamp 1606256979
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3864 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1606256979
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_39
timestamp 1606256979
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1606256979
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606256979
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1606256979
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8740 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7452 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 8464 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_68
timestamp 1606256979
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1606256979
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10396 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1606256979
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1606256979
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14260 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13432 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_140
timestamp 1606256979
transform 1 0 13984 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_159
timestamp 1606256979
transform 1 0 15732 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606256979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19044 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606256979
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 20700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1606256979
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1606256979
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1606256979
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1606256979
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6072 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_48
timestamp 1606256979
transform 1 0 5520 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8096 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_70
timestamp 1606256979
transform 1 0 7544 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9844 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1606256979
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606256979
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1606256979
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10856 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12512 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1606256979
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1606256979
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_138
timestamp 1606256979
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15548 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606256979
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18308 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp 1606256979
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_184
timestamp 1606256979
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19964 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1606256979
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1606256979
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606256979
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1606256979
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1606256979
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1606256979
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606256979
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1606256979
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1606256979
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1606256979
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1606256979
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4784 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6256 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1606256979
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1606256979
transform 1 0 5520 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7268 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1606256979
transform 1 0 8648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1606256979
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_83
timestamp 1606256979
transform 1 0 8740 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1606256979
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1606256979
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10948 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1606256979
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1606256979
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1606256979
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_132
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1606256979
transform 1 0 13800 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1606256979
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 15824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_148
timestamp 1606256979
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_146
timestamp 1606256979
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606256979
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16928 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16836 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1606256979
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1606256979
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_169
timestamp 1606256979
transform 1 0 16652 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18584 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1606256979
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1606256979
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1606256979
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1606256979
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20332 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1606256979
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1606256979
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2392 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1606256979
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1606256979
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_48
timestamp 1606256979
transform 1 0 5520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1606256979
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606256979
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_76
timestamp 1606256979
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10028 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1606256979
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1606256979
transform 1 0 11500 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606256979
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13340 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1606256979
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14996 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1606256979
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16652 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1606256979
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1606256979
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606256979
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18768 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19872 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1606256979
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_198
timestamp 1606256979
transform 1 0 19320 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20608 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1606256979
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606256979
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 1472 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_8
timestamp 1606256979
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_16
timestamp 1606256979
transform 1 0 2576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1606256979
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_36
timestamp 1606256979
transform 1 0 4416 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_48
timestamp 1606256979
transform 1 0 5520 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_60
timestamp 1606256979
transform 1 0 6624 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606256979
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10028 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1606256979
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1606256979
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1606256979
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1606256979
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_132
timestamp 1606256979
transform 1 0 13248 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_138
timestamp 1606256979
transform 1 0 13800 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15732 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1606256979
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606256979
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1606256979
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1606256979
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606256979
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19688 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1606256979
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp 1606256979
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1606256979
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2944 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1606256979
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_17
timestamp 1606256979
transform 1 0 2668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1606256979
transform 1 0 4416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_48
timestamp 1606256979
transform 1 0 5520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1606256979
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1606256979
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1606256979
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1606256979
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1606256979
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_163
timestamp 1606256979
transform 1 0 16100 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1606256979
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1606256979
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 19412 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_196
timestamp 1606256979
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1606256979
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1606256979
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606256979
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606256979
transform 1 0 2300 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1606256979
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_17
timestamp 1606256979
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606256979
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_38
timestamp 1606256979
transform 1 0 4600 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1606256979
transform 1 0 5704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1606256979
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1606256979
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1606256979
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12512 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606256979
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_117
timestamp 1606256979
transform 1 0 11868 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_123
timestamp 1606256979
transform 1 0 12420 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1606256979
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1606256979
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606256979
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606256979
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606256979
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1606256979
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606256979
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606256979
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1606256979
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_17
timestamp 1606256979
transform 1 0 2668 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1606256979
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_26
timestamp 1606256979
transform 1 0 3496 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_38
timestamp 1606256979
transform 1 0 4600 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_50
timestamp 1606256979
transform 1 0 5704 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1606256979
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606256979
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606256979
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606256979
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 13340 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1606256979
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1606256979
transform 1 0 13708 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1606256979
transform 1 0 14812 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_161
timestamp 1606256979
transform 1 0 15916 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1606256979
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1606256979
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1606256979
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1606256979
transform 1 0 19872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1606256979
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606256979
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606256979
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606256979
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606256979
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1606256979
transform 1 0 2116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1606256979
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1606256979
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1606256979
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606256979
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_47
timestamp 1606256979
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606256979
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606256979
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606256979
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1606256979
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1606256979
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1606256979
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606256979
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606256979
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1606256979
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1606256979
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606256979
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1606256979
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1606256979
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606256979
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1606256979
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_202
timestamp 1606256979
transform 1 0 19688 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606256979
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_208
timestamp 1606256979
transform 1 0 20240 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1606256979
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606256979
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606256979
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606256979
transform 1 0 1564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1606256979
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_17
timestamp 1606256979
transform 1 0 2668 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1606256979
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606256979
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1606256979
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606256979
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1606256979
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1606256979
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1606256979
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1606256979
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606256979
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606256979
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_190
timestamp 1606256979
transform 1 0 18584 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_198
timestamp 1606256979
transform 1 0 19320 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_207
timestamp 1606256979
transform 1 0 20148 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1606256979
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606256979
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1606256979
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1606256979
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_47
timestamp 1606256979
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1606256979
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1606256979
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1606256979
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1606256979
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606256979
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606256979
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_208
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606256979
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606256979
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_11
timestamp 1606256979
transform 1 0 2116 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1606256979
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 5980 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_44
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_52
timestamp 1606256979
transform 1 0 5888 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_59
timestamp 1606256979
transform 1 0 6532 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1606256979
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1606256979
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1606256979
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1606256979
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1606256979
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1606256979
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1606256979
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1606256979
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18124 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_178
timestamp 1606256979
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_184
timestamp 1606256979
transform 1 0 18032 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_191
timestamp 1606256979
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_203
timestamp 1606256979
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1606256979
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606256979
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606256979
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606256979
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1606256979
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1606256979
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1606256979
transform 1 0 4876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606256979
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1606256979
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1606256979
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1606256979
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1606256979
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1606256979
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606256979
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606256979
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1606256979
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1606256979
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1606256979
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_198
timestamp 1606256979
transform 1 0 19320 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1606256979
transform 1 0 20424 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606256979
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606256979
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606256979
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606256979
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606256979
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606256979
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606256979
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606256979
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606256979
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 22098 0 22154 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 5722 22320 5778 22800 6 ccff_head
port 10 nsew default input
rlabel metal2 s 17130 22320 17186 22800 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[0]
port 92 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[10]
port 93 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[11]
port 94 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 95 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[13]
port 96 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[14]
port 97 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[15]
port 98 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[16]
port 99 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[17]
port 100 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[18]
port 101 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[19]
port 102 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[1]
port 103 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chany_bottom_in[2]
port 104 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[3]
port 105 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[4]
port 106 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[5]
port 107 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[6]
port 108 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[7]
port 109 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[8]
port 110 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[9]
port 111 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_out[0]
port 112 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[10]
port 113 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[11]
port 114 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[12]
port 115 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[13]
port 116 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[14]
port 117 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[15]
port 118 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[16]
port 119 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[17]
port 120 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[18]
port 121 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[19]
port 122 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[1]
port 123 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_out[2]
port 124 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 chany_bottom_out[3]
port 125 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_out[4]
port 126 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[5]
port 127 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[6]
port 128 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 129 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_out[8]
port 130 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 chany_bottom_out[9]
port 131 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 132 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 133 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 134 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 135 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 136 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 137 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 138 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 139 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 140 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_in
port 141 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 142 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 143 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 144 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 145 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 146 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 147 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 148 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 149 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 150 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 151 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 152 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
