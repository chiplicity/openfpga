magic
tech sky130A
magscale 1 2
timestamp 1606228449
<< locali >>
rect 2053 16643 2087 16745
rect 9413 12087 9447 12257
rect 9045 10591 9079 10761
rect 11529 7939 11563 8041
rect 10517 7803 10551 7905
rect 12265 6103 12299 6205
rect 6653 5559 6687 5661
rect 10609 2295 10643 2601
rect 10701 2295 10735 2533
<< viali >>
rect 1961 20009 1995 20043
rect 2513 20009 2547 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 1961 19465 1995 19499
rect 3065 19465 3099 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 2881 19261 2915 19295
rect 2513 19125 2547 19159
rect 1869 18921 1903 18955
rect 3249 18853 3283 18887
rect 1685 18785 1719 18819
rect 2237 18785 2271 18819
rect 2973 18785 3007 18819
rect 2421 18717 2455 18751
rect 1961 18377 1995 18411
rect 3249 18377 3283 18411
rect 2513 18241 2547 18275
rect 10609 18241 10643 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 3065 18173 3099 18207
rect 10425 18173 10459 18207
rect 1961 17833 1995 17867
rect 11069 17833 11103 17867
rect 2605 17765 2639 17799
rect 3341 17765 3375 17799
rect 7389 17765 7423 17799
rect 9965 17765 9999 17799
rect 11529 17765 11563 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 3065 17697 3099 17731
rect 7113 17697 7147 17731
rect 9689 17697 9723 17731
rect 11437 17697 11471 17731
rect 12081 17697 12115 17731
rect 11713 17629 11747 17663
rect 1685 17289 1719 17323
rect 3709 17289 3743 17323
rect 10333 17289 10367 17323
rect 2329 17153 2363 17187
rect 5089 17153 5123 17187
rect 10977 17153 11011 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 2789 17085 2823 17119
rect 3065 17085 3099 17119
rect 3525 17085 3559 17119
rect 8677 17085 8711 17119
rect 8944 17017 8978 17051
rect 4445 16949 4479 16983
rect 4813 16949 4847 16983
rect 4905 16949 4939 16983
rect 10057 16949 10091 16983
rect 10701 16949 10735 16983
rect 10793 16949 10827 16983
rect 1869 16745 1903 16779
rect 2053 16745 2087 16779
rect 5641 16745 5675 16779
rect 7757 16745 7791 16779
rect 10149 16745 10183 16779
rect 11989 16745 12023 16779
rect 13645 16745 13679 16779
rect 2513 16677 2547 16711
rect 4528 16677 4562 16711
rect 6377 16677 6411 16711
rect 8217 16677 8251 16711
rect 12510 16677 12544 16711
rect 1685 16609 1719 16643
rect 2053 16609 2087 16643
rect 2226 16609 2260 16643
rect 6837 16609 6871 16643
rect 6929 16609 6963 16643
rect 8125 16609 8159 16643
rect 8769 16609 8803 16643
rect 10609 16609 10643 16643
rect 10876 16609 10910 16643
rect 12265 16609 12299 16643
rect 4261 16541 4295 16575
rect 7021 16541 7055 16575
rect 8401 16541 8435 16575
rect 6469 16405 6503 16439
rect 2973 16201 3007 16235
rect 6469 16201 6503 16235
rect 9137 16201 9171 16235
rect 11161 16201 11195 16235
rect 2237 16065 2271 16099
rect 3341 16065 3375 16099
rect 9781 16065 9815 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2789 15997 2823 16031
rect 5089 15997 5123 16031
rect 5356 15997 5390 16031
rect 7757 15997 7791 16031
rect 3608 15929 3642 15963
rect 8024 15929 8058 15963
rect 10048 15929 10082 15963
rect 1685 15861 1719 15895
rect 4721 15861 4755 15895
rect 6837 15861 6871 15895
rect 2881 15657 2915 15691
rect 4721 15657 4755 15691
rect 5089 15657 5123 15691
rect 8861 15657 8895 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 11437 15657 11471 15691
rect 6000 15589 6034 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 3249 15521 3283 15555
rect 4077 15521 4111 15555
rect 5181 15521 5215 15555
rect 7748 15521 7782 15555
rect 10057 15521 10091 15555
rect 11805 15521 11839 15555
rect 11897 15521 11931 15555
rect 3341 15453 3375 15487
rect 3525 15453 3559 15487
rect 4629 15453 4663 15487
rect 5273 15453 5307 15487
rect 5733 15453 5767 15487
rect 7481 15453 7515 15487
rect 10241 15453 10275 15487
rect 11345 15453 11379 15487
rect 12081 15453 12115 15487
rect 1961 15317 1995 15351
rect 2513 15317 2547 15351
rect 7113 15317 7147 15351
rect 10609 15317 10643 15351
rect 3985 15113 4019 15147
rect 4445 15113 4479 15147
rect 5733 15113 5767 15147
rect 7757 15113 7791 15147
rect 10149 15113 10183 15147
rect 10609 15113 10643 15147
rect 2145 14977 2179 15011
rect 4813 14977 4847 15011
rect 6377 14977 6411 15011
rect 8401 14977 8435 15011
rect 11161 14977 11195 15011
rect 1869 14909 1903 14943
rect 2605 14909 2639 14943
rect 4261 14909 4295 14943
rect 6193 14909 6227 14943
rect 8125 14909 8159 14943
rect 8769 14909 8803 14943
rect 2872 14841 2906 14875
rect 6101 14841 6135 14875
rect 9036 14841 9070 14875
rect 10517 14841 10551 14875
rect 8217 14773 8251 14807
rect 10977 14773 11011 14807
rect 11069 14773 11103 14807
rect 4077 14569 4111 14603
rect 7665 14569 7699 14603
rect 7941 14569 7975 14603
rect 8585 14569 8619 14603
rect 10149 14569 10183 14603
rect 4445 14501 4479 14535
rect 6368 14501 6402 14535
rect 1593 14433 1627 14467
rect 2596 14433 2630 14467
rect 4537 14433 4571 14467
rect 6101 14433 6135 14467
rect 7849 14433 7883 14467
rect 8953 14433 8987 14467
rect 10333 14433 10367 14467
rect 1777 14365 1811 14399
rect 2329 14365 2363 14399
rect 4629 14365 4663 14399
rect 5089 14365 5123 14399
rect 9045 14365 9079 14399
rect 9229 14365 9263 14399
rect 9689 14365 9723 14399
rect 3709 14297 3743 14331
rect 7481 14297 7515 14331
rect 8493 14297 8527 14331
rect 4997 14229 5031 14263
rect 3065 14025 3099 14059
rect 5733 14025 5767 14059
rect 10057 14025 10091 14059
rect 1685 13889 1719 13923
rect 2421 13889 2455 13923
rect 3709 13889 3743 13923
rect 6837 13889 6871 13923
rect 1409 13821 1443 13855
rect 2145 13821 2179 13855
rect 3525 13821 3559 13855
rect 4353 13821 4387 13855
rect 8677 13821 8711 13855
rect 4620 13753 4654 13787
rect 7104 13753 7138 13787
rect 8944 13753 8978 13787
rect 3433 13685 3467 13719
rect 6285 13685 6319 13719
rect 8217 13685 8251 13719
rect 3433 13481 3467 13515
rect 5457 13481 5491 13515
rect 5733 13481 5767 13515
rect 7573 13481 7607 13515
rect 8309 13481 8343 13515
rect 8953 13481 8987 13515
rect 11069 13481 11103 13515
rect 2053 13413 2087 13447
rect 7665 13413 7699 13447
rect 1777 13345 1811 13379
rect 2513 13345 2547 13379
rect 3249 13345 3283 13379
rect 4333 13345 4367 13379
rect 6101 13345 6135 13379
rect 6193 13345 6227 13379
rect 8493 13345 8527 13379
rect 9689 13345 9723 13379
rect 9956 13345 9990 13379
rect 2697 13277 2731 13311
rect 4077 13277 4111 13311
rect 6285 13277 6319 13311
rect 7757 13277 7791 13311
rect 9045 13277 9079 13311
rect 9229 13277 9263 13311
rect 8585 13209 8619 13243
rect 7205 13141 7239 13175
rect 1593 12937 1627 12971
rect 1961 12937 1995 12971
rect 3065 12937 3099 12971
rect 6469 12937 6503 12971
rect 6837 12937 6871 12971
rect 10149 12937 10183 12971
rect 4077 12869 4111 12903
rect 2605 12801 2639 12835
rect 3709 12801 3743 12835
rect 4721 12801 4755 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 1409 12733 1443 12767
rect 3525 12733 3559 12767
rect 5089 12733 5123 12767
rect 7205 12733 7239 12767
rect 8769 12733 8803 12767
rect 3433 12665 3467 12699
rect 5356 12665 5390 12699
rect 9036 12665 9070 12699
rect 2329 12597 2363 12631
rect 2421 12597 2455 12631
rect 4445 12597 4479 12631
rect 4537 12597 4571 12631
rect 3157 12393 3191 12427
rect 3617 12393 3651 12427
rect 4353 12393 4387 12427
rect 8585 12393 8619 12427
rect 9689 12393 9723 12427
rect 10701 12393 10735 12427
rect 7012 12325 7046 12359
rect 8953 12325 8987 12359
rect 1777 12257 1811 12291
rect 2044 12257 2078 12291
rect 3433 12257 3467 12291
rect 5080 12257 5114 12291
rect 6653 12257 6687 12291
rect 6745 12257 6779 12291
rect 9413 12257 9447 12291
rect 10057 12257 10091 12291
rect 4813 12189 4847 12223
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 6469 12121 6503 12155
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 6193 12053 6227 12087
rect 8125 12053 8159 12087
rect 9413 12053 9447 12087
rect 1777 11849 1811 11883
rect 6101 11849 6135 11883
rect 8309 11849 8343 11883
rect 10701 11849 10735 11883
rect 2329 11713 2363 11747
rect 4721 11713 4755 11747
rect 7481 11713 7515 11747
rect 7665 11713 7699 11747
rect 8953 11713 8987 11747
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 4629 11645 4663 11679
rect 6653 11645 6687 11679
rect 9321 11645 9355 11679
rect 20269 11645 20303 11679
rect 3056 11577 3090 11611
rect 4988 11577 5022 11611
rect 8677 11577 8711 11611
rect 9588 11577 9622 11611
rect 2145 11509 2179 11543
rect 4169 11509 4203 11543
rect 4445 11509 4479 11543
rect 6469 11509 6503 11543
rect 7021 11509 7055 11543
rect 7389 11509 7423 11543
rect 8769 11509 8803 11543
rect 20453 11509 20487 11543
rect 1869 11305 1903 11339
rect 3525 11305 3559 11339
rect 5457 11305 5491 11339
rect 11069 11305 11103 11339
rect 2789 11237 2823 11271
rect 4445 11237 4479 11271
rect 7012 11237 7046 11271
rect 2697 11169 2731 11203
rect 4537 11169 4571 11203
rect 5825 11169 5859 11203
rect 5917 11169 5951 11203
rect 6745 11169 6779 11203
rect 8769 11169 8803 11203
rect 9956 11169 9990 11203
rect 19717 11169 19751 11203
rect 2973 11101 3007 11135
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 8861 11101 8895 11135
rect 8953 11101 8987 11135
rect 9689 11101 9723 11135
rect 2329 11033 2363 11067
rect 4077 11033 4111 11067
rect 19901 11033 19935 11067
rect 8125 10965 8159 10999
rect 8401 10965 8435 10999
rect 3249 10761 3283 10795
rect 5733 10761 5767 10795
rect 9045 10761 9079 10795
rect 10793 10761 10827 10795
rect 3801 10625 3835 10659
rect 7021 10625 7055 10659
rect 1593 10557 1627 10591
rect 3617 10557 3651 10591
rect 4353 10557 4387 10591
rect 7481 10557 7515 10591
rect 7748 10557 7782 10591
rect 9045 10557 9079 10591
rect 9137 10557 9171 10591
rect 10977 10557 11011 10591
rect 19257 10557 19291 10591
rect 1860 10489 1894 10523
rect 4620 10489 4654 10523
rect 9382 10489 9416 10523
rect 2973 10421 3007 10455
rect 3709 10421 3743 10455
rect 6009 10421 6043 10455
rect 8861 10421 8895 10455
rect 10517 10421 10551 10455
rect 19441 10421 19475 10455
rect 2053 10217 2087 10251
rect 5457 10217 5491 10251
rect 5733 10217 5767 10251
rect 6101 10217 6135 10251
rect 6837 10217 6871 10251
rect 7205 10217 7239 10251
rect 7297 10217 7331 10251
rect 8585 10217 8619 10251
rect 11805 10217 11839 10251
rect 3341 10149 3375 10183
rect 4322 10149 4356 10183
rect 2421 10081 2455 10115
rect 2513 10081 2547 10115
rect 3065 10081 3099 10115
rect 8953 10081 8987 10115
rect 9689 10081 9723 10115
rect 10517 10081 10551 10115
rect 2697 10013 2731 10047
rect 4077 10013 4111 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 7481 10013 7515 10047
rect 9045 10013 9079 10047
rect 9229 10013 9263 10047
rect 3433 9673 3467 9707
rect 8769 9673 8803 9707
rect 3157 9605 3191 9639
rect 4537 9605 4571 9639
rect 5549 9605 5583 9639
rect 3985 9537 4019 9571
rect 5089 9537 5123 9571
rect 6101 9537 6135 9571
rect 7757 9537 7791 9571
rect 9321 9537 9355 9571
rect 1777 9469 1811 9503
rect 4905 9469 4939 9503
rect 2044 9401 2078 9435
rect 6009 9401 6043 9435
rect 9137 9401 9171 9435
rect 3801 9333 3835 9367
rect 3893 9333 3927 9367
rect 4997 9333 5031 9367
rect 5917 9333 5951 9367
rect 7205 9333 7239 9367
rect 7573 9333 7607 9367
rect 7665 9333 7699 9367
rect 9229 9333 9263 9367
rect 1961 9129 1995 9163
rect 2973 9129 3007 9163
rect 4261 9129 4295 9163
rect 4721 9129 4755 9163
rect 8585 9129 8619 9163
rect 9045 9129 9079 9163
rect 2329 9061 2363 9095
rect 8953 9061 8987 9095
rect 3341 8993 3375 9027
rect 4629 8993 4663 9027
rect 5540 8993 5574 9027
rect 6929 8993 6963 9027
rect 7196 8993 7230 9027
rect 9689 8993 9723 9027
rect 9956 8993 9990 9027
rect 2421 8925 2455 8959
rect 2605 8925 2639 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 4905 8925 4939 8959
rect 5273 8925 5307 8959
rect 9229 8925 9263 8959
rect 6653 8789 6687 8823
rect 8309 8789 8343 8823
rect 11069 8789 11103 8823
rect 2789 8585 2823 8619
rect 4445 8585 4479 8619
rect 5733 8585 5767 8619
rect 7849 8585 7883 8619
rect 11161 8585 11195 8619
rect 6285 8449 6319 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8309 8449 8343 8483
rect 8493 8449 8527 8483
rect 9781 8449 9815 8483
rect 1409 8381 1443 8415
rect 1676 8381 1710 8415
rect 3065 8381 3099 8415
rect 5641 8381 5675 8415
rect 9689 8381 9723 8415
rect 3332 8313 3366 8347
rect 8217 8313 8251 8347
rect 10048 8313 10082 8347
rect 5457 8245 5491 8279
rect 6101 8245 6135 8279
rect 6193 8245 6227 8279
rect 6837 8245 6871 8279
rect 7205 8245 7239 8279
rect 9505 8245 9539 8279
rect 11437 8245 11471 8279
rect 1961 8041 1995 8075
rect 2329 8041 2363 8075
rect 2973 8041 3007 8075
rect 4077 8041 4111 8075
rect 6653 8041 6687 8075
rect 8585 8041 8619 8075
rect 10057 8041 10091 8075
rect 11069 8041 11103 8075
rect 11529 8041 11563 8075
rect 13645 8041 13679 8075
rect 5264 7973 5298 8007
rect 3341 7905 3375 7939
rect 4997 7905 5031 7939
rect 7941 7905 7975 7939
rect 8769 7905 8803 7939
rect 10149 7905 10183 7939
rect 10517 7905 10551 7939
rect 11161 7905 11195 7939
rect 11529 7905 11563 7939
rect 11897 7905 11931 7939
rect 12265 7905 12299 7939
rect 12532 7905 12566 7939
rect 17969 7905 18003 7939
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 10333 7837 10367 7871
rect 11345 7837 11379 7871
rect 18245 7837 18279 7871
rect 7573 7769 7607 7803
rect 9689 7769 9723 7803
rect 10517 7769 10551 7803
rect 6377 7701 6411 7735
rect 10701 7701 10735 7735
rect 11713 7701 11747 7735
rect 3617 7497 3651 7531
rect 8401 7497 8435 7531
rect 13829 7497 13863 7531
rect 14105 7429 14139 7463
rect 2513 7361 2547 7395
rect 4169 7361 4203 7395
rect 7941 7361 7975 7395
rect 8953 7361 8987 7395
rect 14657 7361 14691 7395
rect 3985 7293 4019 7327
rect 5089 7293 5123 7327
rect 7849 7293 7883 7327
rect 9597 7293 9631 7327
rect 9864 7293 9898 7327
rect 12449 7293 12483 7327
rect 12716 7293 12750 7327
rect 5356 7225 5390 7259
rect 8861 7225 8895 7259
rect 14565 7225 14599 7259
rect 1961 7157 1995 7191
rect 2329 7157 2363 7191
rect 2421 7157 2455 7191
rect 2973 7157 3007 7191
rect 4077 7157 4111 7191
rect 6469 7157 6503 7191
rect 7389 7157 7423 7191
rect 7757 7157 7791 7191
rect 8769 7157 8803 7191
rect 10977 7157 11011 7191
rect 11253 7157 11287 7191
rect 11897 7157 11931 7191
rect 14473 7157 14507 7191
rect 3617 6953 3651 6987
rect 7113 6953 7147 6987
rect 9045 6953 9079 6987
rect 12541 6953 12575 6987
rect 16681 6953 16715 6987
rect 4445 6885 4479 6919
rect 6000 6885 6034 6919
rect 7656 6885 7690 6919
rect 10416 6885 10450 6919
rect 1501 6817 1535 6851
rect 2504 6817 2538 6851
rect 5733 6817 5767 6851
rect 7389 6817 7423 6851
rect 13452 6817 13486 6851
rect 15568 6817 15602 6851
rect 17417 6817 17451 6851
rect 1685 6749 1719 6783
rect 2237 6749 2271 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 10149 6749 10183 6783
rect 12633 6749 12667 6783
rect 12817 6749 12851 6783
rect 13185 6749 13219 6783
rect 15301 6749 15335 6783
rect 17693 6749 17727 6783
rect 4077 6681 4111 6715
rect 8769 6681 8803 6715
rect 12173 6681 12207 6715
rect 11529 6613 11563 6647
rect 14565 6613 14599 6647
rect 2789 6409 2823 6443
rect 13829 6409 13863 6443
rect 6837 6341 6871 6375
rect 11345 6341 11379 6375
rect 5917 6273 5951 6307
rect 7389 6273 7423 6307
rect 8401 6273 8435 6307
rect 10701 6273 10735 6307
rect 11989 6273 12023 6307
rect 14657 6273 14691 6307
rect 1409 6205 1443 6239
rect 3433 6205 3467 6239
rect 7297 6205 7331 6239
rect 8668 6205 8702 6239
rect 10425 6205 10459 6239
rect 11805 6205 11839 6239
rect 12265 6205 12299 6239
rect 12449 6205 12483 6239
rect 14565 6205 14599 6239
rect 15117 6205 15151 6239
rect 15853 6205 15887 6239
rect 16589 6205 16623 6239
rect 18337 6205 18371 6239
rect 1676 6137 1710 6171
rect 3700 6137 3734 6171
rect 5641 6137 5675 6171
rect 7205 6137 7239 6171
rect 11713 6137 11747 6171
rect 12694 6137 12728 6171
rect 15393 6137 15427 6171
rect 16129 6137 16163 6171
rect 16865 6137 16899 6171
rect 4813 6069 4847 6103
rect 5273 6069 5307 6103
rect 5733 6069 5767 6103
rect 6285 6069 6319 6103
rect 9781 6069 9815 6103
rect 10057 6069 10091 6103
rect 10517 6069 10551 6103
rect 12265 6069 12299 6103
rect 14105 6069 14139 6103
rect 14473 6069 14507 6103
rect 18521 6069 18555 6103
rect 1961 5865 1995 5899
rect 2973 5865 3007 5899
rect 3341 5865 3375 5899
rect 3433 5865 3467 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 6101 5865 6135 5899
rect 8493 5865 8527 5899
rect 9965 5865 9999 5899
rect 10701 5865 10735 5899
rect 12817 5865 12851 5899
rect 13645 5865 13679 5899
rect 6193 5797 6227 5831
rect 10793 5797 10827 5831
rect 11704 5797 11738 5831
rect 15669 5797 15703 5831
rect 2329 5729 2363 5763
rect 6929 5729 6963 5763
rect 7369 5729 7403 5763
rect 10149 5729 10183 5763
rect 13277 5729 13311 5763
rect 15761 5729 15795 5763
rect 16313 5729 16347 5763
rect 16865 5729 16899 5763
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 3617 5661 3651 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 7113 5661 7147 5695
rect 10977 5661 11011 5695
rect 11437 5661 11471 5695
rect 15853 5661 15887 5695
rect 5733 5593 5767 5627
rect 6653 5525 6687 5559
rect 6745 5525 6779 5559
rect 10333 5525 10367 5559
rect 13093 5525 13127 5559
rect 15301 5525 15335 5559
rect 16497 5525 16531 5559
rect 17049 5525 17083 5559
rect 2605 5321 2639 5355
rect 11805 5321 11839 5355
rect 16313 5321 16347 5355
rect 4629 5253 4663 5287
rect 6837 5253 6871 5287
rect 2237 5185 2271 5219
rect 3157 5185 3191 5219
rect 5181 5185 5215 5219
rect 6377 5185 6411 5219
rect 7389 5185 7423 5219
rect 7849 5185 7883 5219
rect 8769 5185 8803 5219
rect 10425 5185 10459 5219
rect 13093 5185 13127 5219
rect 16589 5185 16623 5219
rect 1961 5117 1995 5151
rect 6101 5117 6135 5151
rect 7205 5117 7239 5151
rect 12817 5117 12851 5151
rect 12909 5117 12943 5151
rect 13921 5117 13955 5151
rect 14933 5117 14967 5151
rect 2973 5049 3007 5083
rect 7297 5049 7331 5083
rect 9014 5049 9048 5083
rect 10692 5049 10726 5083
rect 14197 5049 14231 5083
rect 15200 5049 15234 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 3065 4981 3099 5015
rect 4997 4981 5031 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 6193 4981 6227 5015
rect 10149 4981 10183 5015
rect 12449 4981 12483 5015
rect 3065 4777 3099 4811
rect 3341 4777 3375 4811
rect 4077 4777 4111 4811
rect 7021 4777 7055 4811
rect 11897 4777 11931 4811
rect 15669 4777 15703 4811
rect 15761 4777 15795 4811
rect 16313 4777 16347 4811
rect 4445 4709 4479 4743
rect 13369 4709 13403 4743
rect 1952 4641 1986 4675
rect 5641 4641 5675 4675
rect 5908 4641 5942 4675
rect 8125 4641 8159 4675
rect 9689 4641 9723 4675
rect 9956 4641 9990 4675
rect 11805 4641 11839 4675
rect 12449 4641 12483 4675
rect 13093 4641 13127 4675
rect 13829 4641 13863 4675
rect 16681 4641 16715 4675
rect 1685 4573 1719 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 11989 4573 12023 4607
rect 14105 4573 14139 4607
rect 15945 4573 15979 4607
rect 16773 4573 16807 4607
rect 16865 4573 16899 4607
rect 11437 4505 11471 4539
rect 7757 4437 7791 4471
rect 11069 4437 11103 4471
rect 15301 4437 15335 4471
rect 1685 4233 1719 4267
rect 6837 4233 6871 4267
rect 7849 4233 7883 4267
rect 6377 4165 6411 4199
rect 15853 4165 15887 4199
rect 2329 4097 2363 4131
rect 4997 4097 5031 4131
rect 7389 4097 7423 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 9413 4097 9447 4131
rect 10057 4097 10091 4131
rect 13461 4097 13495 4131
rect 2697 4029 2731 4063
rect 7297 4029 7331 4063
rect 8217 4029 8251 4063
rect 13277 4029 13311 4063
rect 14473 4029 14507 4063
rect 17049 4029 17083 4063
rect 19625 4029 19659 4063
rect 19892 4029 19926 4063
rect 2964 3961 2998 3995
rect 5264 3961 5298 3995
rect 10324 3961 10358 3995
rect 13185 3961 13219 3995
rect 14740 3961 14774 3995
rect 17325 3961 17359 3995
rect 2053 3893 2087 3927
rect 2145 3893 2179 3927
rect 4077 3893 4111 3927
rect 7205 3893 7239 3927
rect 8861 3893 8895 3927
rect 9229 3893 9263 3927
rect 9321 3893 9355 3927
rect 11437 3893 11471 3927
rect 11897 3893 11931 3927
rect 12817 3893 12851 3927
rect 16129 3893 16163 3927
rect 21005 3893 21039 3927
rect 2881 3689 2915 3723
rect 13185 3689 13219 3723
rect 15669 3689 15703 3723
rect 4712 3621 4746 3655
rect 6469 3621 6503 3655
rect 9137 3621 9171 3655
rect 12050 3621 12084 3655
rect 13706 3621 13740 3655
rect 1501 3553 1535 3587
rect 1768 3553 1802 3587
rect 7481 3553 7515 3587
rect 7748 3553 7782 3587
rect 10149 3553 10183 3587
rect 10416 3553 10450 3587
rect 11805 3553 11839 3587
rect 15761 3553 15795 3587
rect 16313 3553 16347 3587
rect 17969 3553 18003 3587
rect 20269 3553 20303 3587
rect 4445 3485 4479 3519
rect 6561 3485 6595 3519
rect 6653 3485 6687 3519
rect 9689 3485 9723 3519
rect 13461 3485 13495 3519
rect 15853 3485 15887 3519
rect 16589 3485 16623 3519
rect 5825 3417 5859 3451
rect 11529 3417 11563 3451
rect 14841 3417 14875 3451
rect 6101 3349 6135 3383
rect 8861 3349 8895 3383
rect 15301 3349 15335 3383
rect 18153 3349 18187 3383
rect 20453 3349 20487 3383
rect 5181 3145 5215 3179
rect 5457 3145 5491 3179
rect 9045 3145 9079 3179
rect 11069 3145 11103 3179
rect 3433 3077 3467 3111
rect 10057 3077 10091 3111
rect 12449 3077 12483 3111
rect 2053 3009 2087 3043
rect 3801 3009 3835 3043
rect 6009 3009 6043 3043
rect 7389 3009 7423 3043
rect 9597 3009 9631 3043
rect 10517 3009 10551 3043
rect 10609 3009 10643 3043
rect 11621 3009 11655 3043
rect 13001 3009 13035 3043
rect 7656 2941 7690 2975
rect 9505 2941 9539 2975
rect 13461 2941 13495 2975
rect 14197 2941 14231 2975
rect 14749 2941 14783 2975
rect 15393 2941 15427 2975
rect 16129 2941 16163 2975
rect 16405 2941 16439 2975
rect 17049 2941 17083 2975
rect 18797 2941 18831 2975
rect 20545 2941 20579 2975
rect 2320 2873 2354 2907
rect 4068 2873 4102 2907
rect 5825 2873 5859 2907
rect 12817 2873 12851 2907
rect 13737 2873 13771 2907
rect 15669 2873 15703 2907
rect 20361 2873 20395 2907
rect 5917 2805 5951 2839
rect 8769 2805 8803 2839
rect 9413 2805 9447 2839
rect 10425 2805 10459 2839
rect 11437 2805 11471 2839
rect 11529 2805 11563 2839
rect 12909 2805 12943 2839
rect 14381 2805 14415 2839
rect 14933 2805 14967 2839
rect 17233 2805 17267 2839
rect 18981 2805 19015 2839
rect 20729 2805 20763 2839
rect 2421 2601 2455 2635
rect 4077 2601 4111 2635
rect 4537 2601 4571 2635
rect 5089 2601 5123 2635
rect 5641 2601 5675 2635
rect 6009 2601 6043 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8033 2601 8067 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 10609 2601 10643 2635
rect 10793 2601 10827 2635
rect 6101 2533 6135 2567
rect 8493 2533 8527 2567
rect 2789 2465 2823 2499
rect 4445 2465 4479 2499
rect 7297 2465 7331 2499
rect 8401 2465 8435 2499
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 4629 2397 4663 2431
rect 6285 2397 6319 2431
rect 7481 2397 7515 2431
rect 8677 2397 8711 2431
rect 10333 2397 10367 2431
rect 10609 2261 10643 2295
rect 10701 2533 10735 2567
rect 11161 2533 11195 2567
rect 12081 2533 12115 2567
rect 11253 2465 11287 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 13921 2465 13955 2499
rect 14473 2465 14507 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 11437 2397 11471 2431
rect 12909 2397 12943 2431
rect 16773 2329 16807 2363
rect 10701 2261 10735 2295
rect 13553 2261 13587 2295
rect 14105 2261 14139 2295
rect 14657 2261 14691 2295
rect 15669 2261 15703 2295
rect 16221 2261 16255 2295
rect 17325 2261 17359 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 2774 20040 2780 20052
rect 2547 20012 2780 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19904 2375 19907
rect 4798 19904 4804 19916
rect 2363 19876 4804 19904
rect 2363 19873 2375 19876
rect 2317 19867 2375 19873
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3050 19496 3056 19508
rect 3011 19468 3056 19496
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2130 19292 2136 19304
rect 1811 19264 2136 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 10594 19292 10600 19304
rect 2915 19264 10600 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2866 19156 2872 19168
rect 2547 19128 2872 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1854 18952 1860 18964
rect 1815 18924 1860 18952
rect 1854 18912 1860 18924
rect 1912 18912 1918 18964
rect 7190 18952 7196 18964
rect 2240 18924 7196 18952
rect 2240 18825 2268 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 2314 18844 2320 18896
rect 2372 18884 2378 18896
rect 3237 18887 3295 18893
rect 3237 18884 3249 18887
rect 2372 18856 3249 18884
rect 2372 18844 2378 18856
rect 3237 18853 3249 18856
rect 3283 18853 3295 18887
rect 3237 18847 3295 18853
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18785 2283 18819
rect 2225 18779 2283 18785
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 8386 18816 8392 18828
rect 3007 18788 8392 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 1688 18680 1716 18779
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2409 18751 2467 18757
rect 2409 18748 2421 18751
rect 1820 18720 2421 18748
rect 1820 18708 1826 18720
rect 2409 18717 2421 18720
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 3326 18680 3332 18692
rect 1688 18652 3332 18680
rect 3326 18640 3332 18652
rect 3384 18640 3390 18692
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 3234 18408 3240 18420
rect 3195 18380 3240 18408
rect 3234 18368 3240 18380
rect 3292 18368 3298 18420
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 2188 18244 2513 18272
rect 2188 18232 2194 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 10594 18272 10600 18284
rect 10555 18244 10600 18272
rect 2501 18235 2559 18241
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 1854 18204 1860 18216
rect 1811 18176 1860 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18204 2375 18207
rect 3053 18207 3111 18213
rect 2363 18176 3004 18204
rect 2363 18173 2375 18176
rect 2317 18167 2375 18173
rect 2976 18136 3004 18176
rect 3053 18173 3065 18207
rect 3099 18204 3111 18207
rect 8294 18204 8300 18216
rect 3099 18176 8300 18204
rect 3099 18173 3111 18176
rect 3053 18167 3111 18173
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 11054 18204 11060 18216
rect 10459 18176 11060 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 8662 18136 8668 18148
rect 2976 18108 8668 18136
rect 8662 18096 8668 18108
rect 8720 18096 8726 18148
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 1912 17768 2605 17796
rect 1912 17756 1918 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 3326 17796 3332 17808
rect 3287 17768 3332 17796
rect 2593 17759 2651 17765
rect 3326 17756 3332 17768
rect 3384 17756 3390 17808
rect 4798 17756 4804 17808
rect 4856 17796 4862 17808
rect 7377 17799 7435 17805
rect 7377 17796 7389 17799
rect 4856 17768 7389 17796
rect 4856 17756 4862 17768
rect 7377 17765 7389 17768
rect 7423 17765 7435 17799
rect 7377 17759 7435 17765
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 9953 17799 10011 17805
rect 9953 17796 9965 17799
rect 8352 17768 9965 17796
rect 8352 17756 8358 17768
rect 9953 17765 9965 17768
rect 9999 17765 10011 17799
rect 9953 17759 10011 17765
rect 11517 17799 11575 17805
rect 11517 17765 11529 17799
rect 11563 17796 11575 17799
rect 11606 17796 11612 17808
rect 11563 17768 11612 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 11606 17756 11612 17768
rect 11664 17756 11670 17808
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 3053 17731 3111 17737
rect 2363 17700 3004 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 1780 17660 1808 17691
rect 2866 17660 2872 17672
rect 1780 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 2976 17660 3004 17700
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 7101 17731 7159 17737
rect 3099 17700 7052 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 6270 17660 6276 17672
rect 2976 17632 6276 17660
rect 6270 17620 6276 17632
rect 6328 17620 6334 17672
rect 7024 17660 7052 17700
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7742 17728 7748 17740
rect 7147 17700 7748 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 10318 17728 10324 17740
rect 9723 17700 10324 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11471 17700 12081 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 9030 17660 9036 17672
rect 7024 17632 9036 17660
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 13630 17660 13636 17672
rect 11747 17632 13636 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 13630 17620 13636 17632
rect 13688 17620 13694 17672
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 3694 17320 3700 17332
rect 3655 17292 3700 17320
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 5718 17252 5724 17264
rect 2056 17224 5724 17252
rect 1486 17116 1492 17128
rect 1447 17088 1492 17116
rect 1486 17076 1492 17088
rect 1544 17076 1550 17128
rect 2056 17125 2084 17224
rect 5718 17212 5724 17224
rect 5776 17212 5782 17264
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 5074 17184 5080 17196
rect 2363 17156 3556 17184
rect 5035 17156 5080 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 2792 17048 2820 17079
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3528 17125 3556 17156
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11146 17184 11152 17196
rect 11011 17156 11152 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 3053 17119 3111 17125
rect 3053 17116 3065 17119
rect 2924 17088 3065 17116
rect 2924 17076 2930 17088
rect 3053 17085 3065 17088
rect 3099 17085 3111 17119
rect 3053 17079 3111 17085
rect 3513 17119 3571 17125
rect 3513 17085 3525 17119
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 9766 17116 9772 17128
rect 8711 17088 9772 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 6730 17048 6736 17060
rect 2792 17020 6736 17048
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 8932 17051 8990 17057
rect 8932 17017 8944 17051
rect 8978 17048 8990 17051
rect 9122 17048 9128 17060
rect 8978 17020 9128 17048
rect 8978 17017 8990 17020
rect 8932 17011 8990 17017
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 3844 16952 4445 16980
rect 3844 16940 3850 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4798 16980 4804 16992
rect 4759 16952 4804 16980
rect 4433 16943 4491 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 10042 16980 10048 16992
rect 4948 16952 4993 16980
rect 10003 16952 10048 16980
rect 4948 16940 4954 16952
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 10836 16952 10881 16980
rect 10836 16940 10842 16952
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2041 16779 2099 16785
rect 2041 16745 2053 16779
rect 2087 16776 2099 16779
rect 2087 16748 2728 16776
rect 2087 16745 2099 16748
rect 2041 16739 2099 16745
rect 1486 16668 1492 16720
rect 1544 16708 1550 16720
rect 2501 16711 2559 16717
rect 2501 16708 2513 16711
rect 1544 16680 2513 16708
rect 1544 16668 1550 16680
rect 2501 16677 2513 16680
rect 2547 16677 2559 16711
rect 2700 16708 2728 16748
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5350 16776 5356 16788
rect 5132 16748 5356 16776
rect 5132 16736 5138 16748
rect 5350 16736 5356 16748
rect 5408 16776 5414 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5408 16748 5641 16776
rect 5408 16736 5414 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 7742 16776 7748 16788
rect 7703 16748 7748 16776
rect 5629 16739 5687 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10686 16776 10692 16788
rect 10183 16748 10692 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16745 12035 16779
rect 13630 16776 13636 16788
rect 13543 16748 13636 16776
rect 11977 16739 12035 16745
rect 3786 16708 3792 16720
rect 2700 16680 3792 16708
rect 2501 16671 2559 16677
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4516 16711 4574 16717
rect 4516 16677 4528 16711
rect 4562 16708 4574 16711
rect 4706 16708 4712 16720
rect 4562 16680 4712 16708
rect 4562 16677 4574 16680
rect 4516 16671 4574 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 6365 16711 6423 16717
rect 6365 16677 6377 16711
rect 6411 16708 6423 16711
rect 8205 16711 8263 16717
rect 6411 16680 6960 16708
rect 6411 16677 6423 16680
rect 6365 16671 6423 16677
rect 6932 16652 6960 16680
rect 8205 16677 8217 16711
rect 8251 16708 8263 16711
rect 9582 16708 9588 16720
rect 8251 16680 9588 16708
rect 8251 16677 8263 16680
rect 8205 16671 8263 16677
rect 9582 16668 9588 16680
rect 9640 16668 9646 16720
rect 11992 16708 12020 16739
rect 13630 16736 13636 16748
rect 13688 16776 13694 16788
rect 17862 16776 17868 16788
rect 13688 16748 17868 16776
rect 13688 16736 13694 16748
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 12066 16708 12072 16720
rect 10612 16680 11284 16708
rect 11979 16680 12072 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2214 16643 2272 16649
rect 2214 16640 2226 16643
rect 2087 16612 2226 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2214 16609 2226 16612
rect 2260 16609 2272 16643
rect 2214 16603 2272 16609
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6696 16612 6837 16640
rect 6696 16600 6702 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 8113 16643 8171 16649
rect 6972 16612 7017 16640
rect 6972 16600 6978 16612
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 8159 16612 8769 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 8757 16609 8769 16612
rect 8803 16609 8815 16643
rect 8757 16603 8815 16609
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10612 16649 10640 16680
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 9824 16612 10609 16640
rect 9824 16600 9830 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10864 16643 10922 16649
rect 10864 16609 10876 16643
rect 10910 16640 10922 16643
rect 11146 16640 11152 16652
rect 10910 16612 11152 16640
rect 10910 16609 10922 16612
rect 10864 16603 10922 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 11256 16640 11284 16680
rect 12066 16668 12072 16680
rect 12124 16708 12130 16720
rect 12498 16711 12556 16717
rect 12498 16708 12510 16711
rect 12124 16680 12510 16708
rect 12124 16668 12130 16680
rect 12498 16677 12510 16680
rect 12544 16677 12556 16711
rect 12498 16671 12556 16677
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 11256 16612 12265 16640
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 3384 16544 4261 16572
rect 3384 16532 3390 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 7006 16572 7012 16584
rect 6967 16544 7012 16572
rect 4249 16535 4307 16541
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 9122 16572 9128 16584
rect 8435 16544 9128 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 6052 16204 6469 16232
rect 6052 16192 6058 16204
rect 6457 16201 6469 16204
rect 6503 16232 6515 16235
rect 7006 16232 7012 16244
rect 6503 16204 7012 16232
rect 6503 16201 6515 16204
rect 6457 16195 6515 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 9122 16232 9128 16244
rect 9083 16204 9128 16232
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 11146 16232 11152 16244
rect 11107 16204 11152 16232
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 1670 16056 1676 16108
rect 1728 16096 1734 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 1728 16068 2237 16096
rect 1728 16056 1734 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 3326 16096 3332 16108
rect 3287 16068 3332 16096
rect 2225 16059 2283 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 9766 16096 9772 16108
rect 9727 16068 9772 16096
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 2038 16028 2044 16040
rect 1999 16000 2044 16028
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 2866 16028 2872 16040
rect 2823 16000 2872 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3344 16028 3372 16056
rect 5350 16037 5356 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 3344 16000 5089 16028
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5344 16028 5356 16037
rect 5311 16000 5356 16028
rect 5077 15991 5135 15997
rect 5344 15991 5356 16000
rect 3596 15963 3654 15969
rect 3596 15929 3608 15963
rect 3642 15960 3654 15963
rect 3970 15960 3976 15972
rect 3642 15932 3976 15960
rect 3642 15929 3654 15932
rect 3596 15923 3654 15929
rect 3970 15920 3976 15932
rect 4028 15920 4034 15972
rect 5092 15960 5120 15991
rect 5350 15988 5356 15991
rect 5408 15988 5414 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7524 16000 7757 16028
rect 7524 15988 7530 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 5626 15960 5632 15972
rect 5092 15932 5632 15960
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 8012 15963 8070 15969
rect 8012 15929 8024 15963
rect 8058 15960 8070 15963
rect 8846 15960 8852 15972
rect 8058 15932 8852 15960
rect 8058 15929 8070 15932
rect 8012 15923 8070 15929
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 10042 15969 10048 15972
rect 10036 15960 10048 15969
rect 10003 15932 10048 15960
rect 10036 15923 10048 15932
rect 10042 15920 10048 15923
rect 10100 15920 10106 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 4706 15892 4712 15904
rect 4619 15864 4712 15892
rect 4706 15852 4712 15864
rect 4764 15892 4770 15904
rect 5258 15892 5264 15904
rect 4764 15864 5264 15892
rect 4764 15852 4770 15864
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2096 15660 2881 15688
rect 2096 15648 2102 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 2869 15651 2927 15657
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 4890 15688 4896 15700
rect 4755 15660 4896 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 5077 15691 5135 15697
rect 5077 15657 5089 15691
rect 5123 15688 5135 15691
rect 5166 15688 5172 15700
rect 5123 15660 5172 15688
rect 5123 15657 5135 15660
rect 5077 15651 5135 15657
rect 5166 15648 5172 15660
rect 5224 15688 5230 15700
rect 8846 15688 8852 15700
rect 5224 15660 7880 15688
rect 8807 15660 8852 15688
rect 5224 15648 5230 15660
rect 5994 15629 6000 15632
rect 5988 15620 6000 15629
rect 5955 15592 6000 15620
rect 5988 15583 6000 15592
rect 5994 15580 6000 15583
rect 6052 15580 6058 15632
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 2038 15552 2044 15564
rect 1811 15524 2044 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2314 15552 2320 15564
rect 2275 15524 2320 15552
rect 2314 15512 2320 15524
rect 2372 15512 2378 15564
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3283 15524 4077 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15552 5227 15555
rect 6362 15552 6368 15564
rect 5215 15524 6368 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 3326 15484 3332 15496
rect 3287 15456 3332 15484
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 3513 15487 3571 15493
rect 3513 15453 3525 15487
rect 3559 15484 3571 15487
rect 3970 15484 3976 15496
rect 3559 15456 3976 15484
rect 3559 15453 3571 15456
rect 3513 15447 3571 15453
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 5184 15484 5212 15515
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 7742 15561 7748 15564
rect 7736 15552 7748 15561
rect 7703 15524 7748 15552
rect 7736 15515 7748 15524
rect 7742 15512 7748 15515
rect 7800 15512 7806 15564
rect 7852 15552 7880 15660
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9640 15660 9689 15688
rect 9640 15648 9646 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 11146 15688 11152 15700
rect 10183 15660 11152 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 11606 15688 11612 15700
rect 11471 15660 11612 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 8864 15620 8892 15648
rect 8864 15592 10180 15620
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 7852 15524 10057 15552
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10152 15552 10180 15592
rect 11793 15555 11851 15561
rect 11793 15552 11805 15555
rect 10152 15524 10272 15552
rect 10045 15515 10103 15521
rect 4663 15456 5212 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 5316 15456 5361 15484
rect 5316 15444 5322 15456
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5684 15456 5733 15484
rect 5684 15444 5690 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 7466 15484 7472 15496
rect 5721 15447 5779 15453
rect 6748 15456 7472 15484
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 2501 15351 2559 15357
rect 2501 15317 2513 15351
rect 2547 15348 2559 15351
rect 2774 15348 2780 15360
rect 2547 15320 2780 15348
rect 2547 15317 2559 15320
rect 2501 15311 2559 15317
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 5736 15348 5764 15447
rect 6748 15348 6776 15456
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 10244 15493 10272 15524
rect 10336 15524 11805 15552
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 7098 15348 7104 15360
rect 5736 15320 6776 15348
rect 7059 15320 7104 15348
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 10336 15348 10364 15524
rect 11793 15521 11805 15524
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 12250 15552 12256 15564
rect 11931 15524 12256 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11900 15484 11928 15515
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 12066 15484 12072 15496
rect 11379 15456 11928 15484
rect 12027 15456 12072 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 7708 15320 10364 15348
rect 10597 15351 10655 15357
rect 7708 15308 7714 15320
rect 10597 15317 10609 15351
rect 10643 15348 10655 15351
rect 11146 15348 11152 15360
rect 10643 15320 11152 15348
rect 10643 15317 10655 15320
rect 10597 15311 10655 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2866 15144 2872 15156
rect 2148 15116 2872 15144
rect 2148 15017 2176 15116
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 3970 15144 3976 15156
rect 3931 15116 3976 15144
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4433 15147 4491 15153
rect 4433 15144 4445 15147
rect 4212 15116 4445 15144
rect 4212 15104 4218 15116
rect 4433 15113 4445 15116
rect 4479 15113 4491 15147
rect 5718 15144 5724 15156
rect 5679 15116 5724 15144
rect 4433 15107 4491 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7248 15116 7757 15144
rect 7248 15104 7254 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 7745 15107 7803 15113
rect 8772 15116 10149 15144
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 14977 2191 15011
rect 4798 15008 4804 15020
rect 4759 14980 4804 15008
rect 2133 14971 2191 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 7098 15008 7104 15020
rect 6411 14980 7104 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 7800 14980 8401 15008
rect 7800 14968 7806 14980
rect 8389 14977 8401 14980
rect 8435 15008 8447 15011
rect 8772 15008 8800 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10778 15144 10784 15156
rect 10643 15116 10784 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 8435 14980 8800 15008
rect 8435 14977 8447 14980
rect 8389 14971 8447 14977
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10100 14980 11161 15008
rect 10100 14968 10106 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 1854 14940 1860 14952
rect 1815 14912 1860 14940
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 2590 14940 2596 14952
rect 2551 14912 2596 14940
rect 2590 14900 2596 14912
rect 2648 14900 2654 14952
rect 2682 14900 2688 14952
rect 2740 14940 2746 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 2740 14912 4261 14940
rect 2740 14900 2746 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 6181 14943 6239 14949
rect 6181 14909 6193 14943
rect 6227 14940 6239 14943
rect 6454 14940 6460 14952
rect 6227 14912 6460 14940
rect 6227 14909 6239 14912
rect 6181 14903 6239 14909
rect 6454 14900 6460 14912
rect 6512 14900 6518 14952
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 8113 14943 8171 14949
rect 6696 14912 8055 14940
rect 6696 14900 6702 14912
rect 2860 14875 2918 14881
rect 2860 14841 2872 14875
rect 2906 14872 2918 14875
rect 3694 14872 3700 14884
rect 2906 14844 3700 14872
rect 2906 14841 2918 14844
rect 2860 14835 2918 14841
rect 3694 14832 3700 14844
rect 3752 14832 3758 14884
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6822 14872 6828 14884
rect 6135 14844 6828 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 8027 14872 8055 14912
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 8202 14940 8208 14952
rect 8159 14912 8208 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14940 8815 14943
rect 9766 14940 9772 14952
rect 8803 14912 9772 14940
rect 8803 14909 8815 14912
rect 8757 14903 8815 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 9024 14875 9082 14881
rect 8027 14844 8708 14872
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 8570 14804 8576 14816
rect 8251 14776 8576 14804
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8680 14804 8708 14844
rect 9024 14841 9036 14875
rect 9070 14872 9082 14875
rect 9306 14872 9312 14884
rect 9070 14844 9312 14872
rect 9070 14841 9082 14844
rect 9024 14835 9082 14841
rect 9306 14832 9312 14844
rect 9364 14832 9370 14884
rect 10505 14875 10563 14881
rect 10505 14841 10517 14875
rect 10551 14872 10563 14875
rect 10551 14844 11100 14872
rect 10551 14841 10563 14844
rect 10505 14835 10563 14841
rect 11072 14813 11100 14844
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 8680 14776 10977 14804
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 10965 14767 11023 14773
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11606 14804 11612 14816
rect 11103 14776 11612 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3384 14572 4077 14600
rect 3384 14560 3390 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7524 14572 7665 14600
rect 7524 14560 7530 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 7929 14603 7987 14609
rect 7929 14569 7941 14603
rect 7975 14600 7987 14603
rect 8202 14600 8208 14612
rect 7975 14572 8208 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9824 14572 10149 14600
rect 9824 14560 9830 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 3050 14532 3056 14544
rect 1596 14504 3056 14532
rect 1596 14473 1624 14504
rect 3050 14492 3056 14504
rect 3108 14492 3114 14544
rect 4433 14535 4491 14541
rect 4433 14501 4445 14535
rect 4479 14532 4491 14535
rect 6356 14535 6414 14541
rect 4479 14504 6316 14532
rect 4479 14501 4491 14504
rect 4433 14495 4491 14501
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14433 1639 14467
rect 1581 14427 1639 14433
rect 2584 14467 2642 14473
rect 2584 14433 2596 14467
rect 2630 14464 2642 14467
rect 3602 14464 3608 14476
rect 2630 14436 3608 14464
rect 2630 14433 2642 14436
rect 2584 14427 2642 14433
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 4571 14436 4752 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1544 14368 1777 14396
rect 1544 14356 1550 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 1765 14359 1823 14365
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 2332 14260 2360 14359
rect 3694 14328 3700 14340
rect 3655 14300 3700 14328
rect 3694 14288 3700 14300
rect 3752 14328 3758 14340
rect 4632 14328 4660 14359
rect 3752 14300 4660 14328
rect 3752 14288 3758 14300
rect 2590 14260 2596 14272
rect 2332 14232 2596 14260
rect 2590 14220 2596 14232
rect 2648 14260 2654 14272
rect 4246 14260 4252 14272
rect 2648 14232 4252 14260
rect 2648 14220 2654 14232
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4724 14260 4752 14436
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 6089 14467 6147 14473
rect 6089 14464 6101 14467
rect 5684 14436 6101 14464
rect 5684 14424 5690 14436
rect 6089 14433 6101 14436
rect 6135 14464 6147 14467
rect 6178 14464 6184 14476
rect 6135 14436 6184 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 6288 14464 6316 14504
rect 6356 14501 6368 14535
rect 6402 14532 6414 14535
rect 7098 14532 7104 14544
rect 6402 14504 7104 14532
rect 6402 14501 6414 14504
rect 6356 14495 6414 14501
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 8294 14532 8300 14544
rect 7852 14504 8300 14532
rect 7852 14473 7880 14504
rect 8294 14492 8300 14504
rect 8352 14532 8358 14544
rect 8352 14504 10364 14532
rect 8352 14492 8358 14504
rect 10336 14473 10364 14504
rect 7837 14467 7895 14473
rect 6288 14436 7788 14464
rect 5074 14396 5080 14408
rect 5035 14368 5080 14396
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 7760 14396 7788 14436
rect 7837 14433 7849 14467
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14433 10379 14467
rect 10321 14427 10379 14433
rect 8846 14396 8852 14408
rect 7760 14368 8852 14396
rect 8846 14356 8852 14368
rect 8904 14396 8910 14408
rect 8956 14396 8984 14427
rect 8904 14368 8984 14396
rect 9033 14399 9091 14405
rect 8904 14356 8910 14368
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9306 14396 9312 14408
rect 9263 14368 9312 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 7469 14331 7527 14337
rect 7469 14297 7481 14331
rect 7515 14328 7527 14331
rect 7742 14328 7748 14340
rect 7515 14300 7748 14328
rect 7515 14297 7527 14300
rect 7469 14291 7527 14297
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 8481 14331 8539 14337
rect 8481 14297 8493 14331
rect 8527 14328 8539 14331
rect 9048 14328 9076 14359
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10870 14328 10876 14340
rect 8527 14300 10876 14328
rect 8527 14297 8539 14300
rect 8481 14291 8539 14297
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 4985 14263 5043 14269
rect 4985 14260 4997 14263
rect 4724 14232 4997 14260
rect 4985 14229 4997 14232
rect 5031 14260 5043 14263
rect 7098 14260 7104 14272
rect 5031 14232 7104 14260
rect 5031 14229 5043 14232
rect 4985 14223 5043 14229
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1854 14016 1860 14068
rect 1912 14056 1918 14068
rect 3053 14059 3111 14065
rect 3053 14056 3065 14059
rect 1912 14028 3065 14056
rect 1912 14016 1918 14028
rect 3053 14025 3065 14028
rect 3099 14025 3111 14059
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 3053 14019 3111 14025
rect 3988 14028 5733 14056
rect 3234 13988 3240 14000
rect 1412 13960 3240 13988
rect 1412 13861 1440 13960
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 2314 13920 2320 13932
rect 1719 13892 2320 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 2682 13920 2688 13932
rect 2455 13892 2688 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3660 13892 3709 13920
rect 3660 13880 3666 13892
rect 3697 13889 3709 13892
rect 3743 13920 3755 13923
rect 3988 13920 4016 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 5721 14019 5779 14025
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9364 14028 10057 14056
rect 9364 14016 9370 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 3743 13892 4016 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 6546 13920 6552 13932
rect 6236 13892 6552 13920
rect 6236 13880 6242 13892
rect 6546 13880 6552 13892
rect 6604 13920 6610 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6604 13892 6837 13920
rect 6604 13880 6610 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1397 13815 1455 13821
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 3513 13855 3571 13861
rect 2179 13824 3464 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 3436 13784 3464 13824
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3559 13824 4292 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3786 13784 3792 13796
rect 3436 13756 3792 13784
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 4264 13784 4292 13824
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 5718 13852 5724 13864
rect 4396 13824 4441 13852
rect 4540 13824 5724 13852
rect 4396 13812 4402 13824
rect 4540 13784 4568 13824
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 9766 13852 9772 13864
rect 8711 13824 9772 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 4264 13756 4568 13784
rect 4608 13787 4666 13793
rect 4608 13753 4620 13787
rect 4654 13784 4666 13787
rect 5442 13784 5448 13796
rect 4654 13756 5448 13784
rect 4654 13753 4666 13756
rect 4608 13747 4666 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 7092 13787 7150 13793
rect 7092 13753 7104 13787
rect 7138 13784 7150 13787
rect 7742 13784 7748 13796
rect 7138 13756 7748 13784
rect 7138 13753 7150 13756
rect 7092 13747 7150 13753
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 8932 13787 8990 13793
rect 8932 13753 8944 13787
rect 8978 13784 8990 13787
rect 9214 13784 9220 13796
rect 8978 13756 9220 13784
rect 8978 13753 8990 13756
rect 8932 13747 8990 13753
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 3421 13719 3479 13725
rect 3421 13685 3433 13719
rect 3467 13716 3479 13719
rect 5074 13716 5080 13728
rect 3467 13688 5080 13716
rect 3467 13685 3479 13688
rect 3421 13679 3479 13685
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 7190 13716 7196 13728
rect 6319 13688 7196 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 3418 13512 3424 13524
rect 3379 13484 3424 13512
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 5442 13512 5448 13524
rect 5403 13484 5448 13512
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8941 13515 8999 13521
rect 8941 13481 8953 13515
rect 8987 13512 8999 13515
rect 9674 13512 9680 13524
rect 8987 13484 9680 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 2038 13444 2044 13456
rect 1999 13416 2044 13444
rect 2038 13404 2044 13416
rect 2096 13404 2102 13456
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 7576 13444 7604 13472
rect 2280 13416 7604 13444
rect 7653 13447 7711 13453
rect 2280 13404 2286 13416
rect 7653 13413 7665 13447
rect 7699 13444 7711 13447
rect 8570 13444 8576 13456
rect 7699 13416 8576 13444
rect 7699 13413 7711 13416
rect 7653 13407 7711 13413
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 11072 13444 11100 13475
rect 9600 13416 11100 13444
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2498 13376 2504 13388
rect 2459 13348 2504 13376
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 1670 13200 1676 13252
rect 1728 13240 1734 13252
rect 3252 13240 3280 13339
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4321 13379 4379 13385
rect 4321 13376 4333 13379
rect 4212 13348 4333 13376
rect 4212 13336 4218 13348
rect 4321 13345 4333 13348
rect 4367 13345 4379 13379
rect 6086 13376 6092 13388
rect 6047 13348 6092 13376
rect 4321 13339 4379 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6454 13376 6460 13388
rect 6227 13348 6460 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 8478 13376 8484 13388
rect 8439 13348 8484 13376
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 1728 13212 3280 13240
rect 1728 13200 1734 13212
rect 4080 13172 4108 13271
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 5500 13280 6285 13308
rect 5500 13268 5506 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 9033 13311 9091 13317
rect 7800 13280 7845 13308
rect 7800 13268 7806 13280
rect 9033 13277 9045 13311
rect 9079 13277 9091 13311
rect 9214 13308 9220 13320
rect 9127 13280 9220 13308
rect 9033 13271 9091 13277
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8573 13243 8631 13249
rect 8573 13240 8585 13243
rect 8444 13212 8585 13240
rect 8444 13200 8450 13212
rect 8573 13209 8585 13212
rect 8619 13209 8631 13243
rect 8573 13203 8631 13209
rect 5166 13172 5172 13184
rect 4080 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7282 13172 7288 13184
rect 7239 13144 7288 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 9048 13172 9076 13271
rect 9214 13268 9220 13280
rect 9272 13308 9278 13320
rect 9600 13308 9628 13416
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9766 13376 9772 13388
rect 9723 13348 9772 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 9950 13385 9956 13388
rect 9944 13339 9956 13385
rect 10008 13376 10014 13388
rect 10008 13348 10044 13376
rect 9950 13336 9956 13339
rect 10008 13336 10014 13348
rect 9272 13280 9628 13308
rect 9272 13268 9278 13280
rect 9674 13172 9680 13184
rect 9048 13144 9680 13172
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 1949 12971 2007 12977
rect 1949 12968 1961 12971
rect 1820 12940 1961 12968
rect 1820 12928 1826 12940
rect 1949 12937 1961 12940
rect 1995 12937 2007 12971
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 1949 12931 2007 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4154 12968 4160 12980
rect 3712 12940 4160 12968
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 3142 12832 3148 12844
rect 2639 12804 3148 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3712 12841 3740 12940
rect 4154 12928 4160 12940
rect 4212 12968 4218 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 4212 12940 6469 12968
rect 4212 12928 4218 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6788 12940 6837 12968
rect 6788 12928 6794 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8662 12968 8668 12980
rect 8444 12940 8668 12968
rect 8444 12928 8450 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10137 12971 10195 12977
rect 10137 12968 10149 12971
rect 10008 12940 10149 12968
rect 10008 12928 10014 12940
rect 10137 12937 10149 12940
rect 10183 12937 10195 12971
rect 10137 12931 10195 12937
rect 3786 12860 3792 12912
rect 3844 12900 3850 12912
rect 4065 12903 4123 12909
rect 4065 12900 4077 12903
rect 3844 12872 4077 12900
rect 3844 12860 3850 12872
rect 4065 12869 4077 12872
rect 4111 12869 4123 12903
rect 4065 12863 4123 12869
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 4982 12832 4988 12844
rect 4755 12804 4988 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7466 12832 7472 12844
rect 7379 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12832 7530 12844
rect 8202 12832 8208 12844
rect 7524 12804 8208 12832
rect 7524 12792 7530 12804
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2682 12764 2688 12776
rect 1443 12736 2688 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 4614 12764 4620 12776
rect 3559 12736 4620 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5166 12764 5172 12776
rect 5123 12736 5172 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 8757 12767 8815 12773
rect 8757 12733 8769 12767
rect 8803 12764 8815 12767
rect 9306 12764 9312 12776
rect 8803 12736 9312 12764
rect 8803 12733 8815 12736
rect 8757 12727 8815 12733
rect 9306 12724 9312 12736
rect 9364 12764 9370 12776
rect 9766 12764 9772 12776
rect 9364 12736 9772 12764
rect 9364 12724 9370 12736
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 3421 12699 3479 12705
rect 3421 12665 3433 12699
rect 3467 12696 3479 12699
rect 4338 12696 4344 12708
rect 3467 12668 4344 12696
rect 3467 12665 3479 12668
rect 3421 12659 3479 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 5344 12699 5402 12705
rect 5344 12665 5356 12699
rect 5390 12696 5402 12699
rect 6178 12696 6184 12708
rect 5390 12668 6184 12696
rect 5390 12665 5402 12668
rect 5344 12659 5402 12665
rect 6178 12656 6184 12668
rect 6236 12656 6242 12708
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 8846 12696 8852 12708
rect 8260 12668 8852 12696
rect 8260 12656 8266 12668
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 9024 12699 9082 12705
rect 9024 12665 9036 12699
rect 9070 12696 9082 12699
rect 9214 12696 9220 12708
rect 9070 12668 9220 12696
rect 9070 12665 9082 12668
rect 9024 12659 9082 12665
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 2314 12628 2320 12640
rect 2275 12600 2320 12628
rect 2314 12588 2320 12600
rect 2372 12588 2378 12640
rect 2409 12631 2467 12637
rect 2409 12597 2421 12631
rect 2455 12628 2467 12631
rect 2958 12628 2964 12640
rect 2455 12600 2964 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4433 12631 4491 12637
rect 4433 12628 4445 12631
rect 4212 12600 4445 12628
rect 4212 12588 4218 12600
rect 4433 12597 4445 12600
rect 4479 12597 4491 12631
rect 4433 12591 4491 12597
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 5534 12628 5540 12640
rect 4571 12600 5540 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6638 12628 6644 12640
rect 6512 12600 6644 12628
rect 6512 12588 6518 12600
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 10778 12628 10784 12640
rect 8536 12600 10784 12628
rect 8536 12588 8542 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 2314 12424 2320 12436
rect 1820 12396 2320 12424
rect 1820 12384 1826 12396
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 3142 12424 3148 12436
rect 3103 12396 3148 12424
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3602 12424 3608 12436
rect 3563 12396 3608 12424
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 4448 12396 6960 12424
rect 2774 12356 2780 12368
rect 1780 12328 2780 12356
rect 1780 12297 1808 12328
rect 2774 12316 2780 12328
rect 2832 12316 2838 12368
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4448 12356 4476 12396
rect 4120 12328 4476 12356
rect 4120 12316 4126 12328
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 6604 12328 6776 12356
rect 6604 12316 6610 12328
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 2032 12291 2090 12297
rect 2032 12257 2044 12291
rect 2078 12288 2090 12291
rect 2314 12288 2320 12300
rect 2078 12260 2320 12288
rect 2078 12257 2090 12260
rect 2032 12251 2090 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 5074 12297 5080 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3384 12260 3433 12288
rect 3384 12248 3390 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 5068 12288 5080 12297
rect 5035 12260 5080 12288
rect 3421 12251 3479 12257
rect 5068 12251 5080 12260
rect 5074 12248 5080 12251
rect 5132 12248 5138 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 6748 12297 6776 12328
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6512 12260 6653 12288
rect 6512 12248 6518 12260
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12257 6791 12291
rect 6932 12288 6960 12396
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8444 12396 8585 12424
rect 8444 12384 8450 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 8573 12387 8631 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 9876 12396 10701 12424
rect 7000 12359 7058 12365
rect 7000 12325 7012 12359
rect 7046 12356 7058 12359
rect 7466 12356 7472 12368
rect 7046 12328 7472 12356
rect 7046 12325 7058 12328
rect 7000 12319 7058 12325
rect 7466 12316 7472 12328
rect 7524 12316 7530 12368
rect 8941 12359 8999 12365
rect 8941 12325 8953 12359
rect 8987 12356 8999 12359
rect 9876 12356 9904 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 8987 12328 9904 12356
rect 8987 12325 8999 12328
rect 8941 12319 8999 12325
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10008 12328 10272 12356
rect 10008 12316 10014 12328
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 6932 12260 9413 12288
rect 6733 12251 6791 12257
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 4816 12152 4844 12183
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6546 12220 6552 12232
rect 6144 12192 6552 12220
rect 6144 12180 6150 12192
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 9033 12223 9091 12229
rect 9033 12220 9045 12223
rect 8352 12192 9045 12220
rect 8352 12180 8358 12192
rect 9033 12189 9045 12192
rect 9079 12189 9091 12223
rect 9214 12220 9220 12232
rect 9175 12192 9220 12220
rect 9033 12183 9091 12189
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 6457 12155 6515 12161
rect 6457 12152 6469 12155
rect 4764 12124 4844 12152
rect 5736 12124 6469 12152
rect 4764 12112 4770 12124
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5736 12084 5764 12124
rect 6457 12121 6469 12124
rect 6503 12152 6515 12155
rect 6730 12152 6736 12164
rect 6503 12124 6736 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 10060 12152 10088 12251
rect 10244 12229 10272 12328
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 7668 12124 10088 12152
rect 10152 12152 10180 12183
rect 10318 12152 10324 12164
rect 10152 12124 10324 12152
rect 4856 12056 5764 12084
rect 4856 12044 4862 12056
rect 6086 12044 6092 12096
rect 6144 12084 6150 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 6144 12056 6193 12084
rect 6144 12044 6150 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 7668 12084 7696 12124
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 6604 12056 7696 12084
rect 8113 12087 8171 12093
rect 6604 12044 6610 12056
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8938 12084 8944 12096
rect 8159 12056 8944 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 11698 12084 11704 12096
rect 9447 12056 11704 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1762 11880 1768 11892
rect 1723 11852 1768 11880
rect 1762 11840 1768 11852
rect 1820 11840 1826 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 6089 11883 6147 11889
rect 6089 11880 6101 11883
rect 5132 11852 6101 11880
rect 5132 11840 5138 11852
rect 6089 11849 6101 11852
rect 6135 11849 6147 11883
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 6089 11843 6147 11849
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 9272 11852 10701 11880
rect 9272 11840 9278 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 2314 11744 2320 11756
rect 2275 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11744 2378 11756
rect 2372 11716 2912 11744
rect 2372 11704 2378 11716
rect 2884 11688 2912 11716
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4304 11716 4721 11744
rect 4304 11704 4310 11716
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 2866 11636 2872 11688
rect 2924 11636 2930 11688
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11645 4675 11679
rect 4724 11676 4752 11707
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 7156 11716 7481 11744
rect 7156 11704 7162 11716
rect 7469 11713 7481 11716
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 8846 11744 8852 11756
rect 7699 11716 8852 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 8987 11716 9444 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 4798 11676 4804 11688
rect 4724 11648 4804 11676
rect 4617 11639 4675 11645
rect 3044 11611 3102 11617
rect 3044 11577 3056 11611
rect 3090 11608 3102 11611
rect 3142 11608 3148 11620
rect 3090 11580 3148 11608
rect 3090 11577 3102 11580
rect 3044 11571 3102 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3252 11580 4384 11608
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 1912 11512 2145 11540
rect 1912 11500 1918 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2133 11503 2191 11509
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3252 11540 3280 11580
rect 4356 11552 4384 11580
rect 2832 11512 3280 11540
rect 4157 11543 4215 11549
rect 2832 11500 2838 11512
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 4246 11540 4252 11552
rect 4203 11512 4252 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4396 11512 4445 11540
rect 4396 11500 4402 11512
rect 4433 11509 4445 11512
rect 4479 11540 4491 11543
rect 4522 11540 4528 11552
rect 4479 11512 4528 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4632 11540 4660 11639
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5258 11676 5264 11688
rect 4908 11648 5264 11676
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 4908 11608 4936 11648
rect 5258 11636 5264 11648
rect 5316 11676 5322 11688
rect 5994 11676 6000 11688
rect 5316 11648 6000 11676
rect 5316 11636 5322 11648
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 8478 11676 8484 11688
rect 6687 11648 8484 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 9306 11676 9312 11688
rect 9267 11648 9312 11676
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 4764 11580 4936 11608
rect 4976 11611 5034 11617
rect 4764 11568 4770 11580
rect 4976 11577 4988 11611
rect 5022 11608 5034 11611
rect 5626 11608 5632 11620
rect 5022 11580 5632 11608
rect 5022 11577 5034 11580
rect 4976 11571 5034 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 8662 11608 8668 11620
rect 5868 11580 8668 11608
rect 5868 11568 5874 11580
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 6454 11540 6460 11552
rect 4632 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 8754 11540 8760 11552
rect 8715 11512 8760 11540
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 9324 11540 9352 11636
rect 9416 11608 9444 11716
rect 20254 11676 20260 11688
rect 20215 11648 20260 11676
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 9576 11611 9634 11617
rect 9576 11608 9588 11611
rect 9416 11580 9588 11608
rect 9576 11577 9588 11580
rect 9622 11608 9634 11611
rect 11054 11608 11060 11620
rect 9622 11580 11060 11608
rect 9622 11577 9634 11580
rect 9576 11571 9634 11577
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 9766 11540 9772 11552
rect 9324 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 20441 11543 20499 11549
rect 20441 11509 20453 11543
rect 20487 11540 20499 11543
rect 20898 11540 20904 11552
rect 20487 11512 20904 11540
rect 20487 11509 20499 11512
rect 20441 11503 20499 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 4154 11336 4160 11348
rect 3559 11308 4160 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4706 11336 4712 11348
rect 4356 11308 4712 11336
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11268 2835 11271
rect 4356 11268 4384 11308
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4948 11308 5457 11336
rect 4948 11296 4954 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 9950 11336 9956 11348
rect 8812 11308 9956 11336
rect 8812 11296 8818 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 20254 11336 20260 11348
rect 11756 11308 20260 11336
rect 11756 11296 11762 11308
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 2823 11240 4384 11268
rect 4433 11271 4491 11277
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 4433 11237 4445 11271
rect 4479 11268 4491 11271
rect 5718 11268 5724 11280
rect 4479 11240 5724 11268
rect 4479 11237 4491 11240
rect 4433 11231 4491 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 7000 11271 7058 11277
rect 7000 11237 7012 11271
rect 7046 11268 7058 11271
rect 8938 11268 8944 11280
rect 7046 11240 8944 11268
rect 7046 11237 7058 11240
rect 7000 11231 7058 11237
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 9640 11240 12296 11268
rect 9640 11228 9646 11240
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 4525 11203 4583 11209
rect 2731 11172 4476 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3142 11132 3148 11144
rect 3007 11104 3148 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3292 11104 4108 11132
rect 3292 11092 3298 11104
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 3602 11064 3608 11076
rect 2363 11036 3608 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 4080 11073 4108 11104
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11033 4123 11067
rect 4448 11064 4476 11172
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4706 11200 4712 11212
rect 4571 11172 4712 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11200 5963 11203
rect 6178 11200 6184 11212
rect 5951 11172 6184 11200
rect 5951 11169 5963 11172
rect 5905 11163 5963 11169
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 8754 11200 8760 11212
rect 8715 11172 8760 11200
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9944 11203 10002 11209
rect 9944 11169 9956 11203
rect 9990 11200 10002 11203
rect 10410 11200 10416 11212
rect 9990 11172 10416 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 12268 11200 12296 11240
rect 12268 11172 12388 11200
rect 12360 11144 12388 11172
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 12492 11172 19717 11200
rect 12492 11160 12498 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4798 11132 4804 11144
rect 4663 11104 4804 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 6086 11132 6092 11144
rect 6047 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 8846 11132 8852 11144
rect 8807 11104 8852 11132
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 8996 11104 9041 11132
rect 8996 11092 9002 11104
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9732 11104 9777 11132
rect 9732 11092 9738 11104
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 5166 11064 5172 11076
rect 4448 11036 5172 11064
rect 4065 11027 4123 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 19889 11067 19947 11073
rect 7944 11036 8524 11064
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 7944 10996 7972 11036
rect 8110 10996 8116 11008
rect 4028 10968 7972 10996
rect 8071 10968 8116 10996
rect 4028 10956 4034 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8386 10996 8392 11008
rect 8347 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 8496 10996 8524 11036
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 20622 11064 20628 11076
rect 19935 11036 20628 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 11054 10996 11060 11008
rect 8496 10968 11060 10996
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3016 10764 3249 10792
rect 3016 10752 3022 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 3237 10755 3295 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5684 10764 5733 10792
rect 5684 10752 5690 10764
rect 5721 10761 5733 10764
rect 5767 10761 5779 10795
rect 5721 10755 5779 10761
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9766 10792 9772 10804
rect 9079 10764 9772 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 2924 10628 3801 10656
rect 2924 10616 2930 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7374 10656 7380 10668
rect 7055 10628 7380 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 8496 10628 9260 10656
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10588 1639 10591
rect 2774 10588 2780 10600
rect 1627 10560 2780 10588
rect 1627 10557 1639 10560
rect 1581 10551 1639 10557
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 3602 10588 3608 10600
rect 3563 10560 3608 10588
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 4890 10588 4896 10600
rect 4387 10560 4896 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 5132 10560 7481 10588
rect 5132 10548 5138 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7558 10548 7564 10600
rect 7616 10588 7622 10600
rect 7736 10591 7794 10597
rect 7736 10588 7748 10591
rect 7616 10560 7748 10588
rect 7616 10548 7622 10560
rect 7736 10557 7748 10560
rect 7782 10588 7794 10591
rect 8110 10588 8116 10600
rect 7782 10560 8116 10588
rect 7782 10557 7794 10560
rect 7736 10551 7794 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 1848 10523 1906 10529
rect 1848 10489 1860 10523
rect 1894 10520 1906 10523
rect 3142 10520 3148 10532
rect 1894 10492 3148 10520
rect 1894 10489 1906 10492
rect 1848 10483 1906 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 4608 10523 4666 10529
rect 4608 10489 4620 10523
rect 4654 10520 4666 10523
rect 4798 10520 4804 10532
rect 4654 10492 4804 10520
rect 4654 10489 4666 10492
rect 4608 10483 4666 10489
rect 4798 10480 4804 10492
rect 4856 10520 4862 10532
rect 5442 10520 5448 10532
rect 4856 10492 5448 10520
rect 4856 10480 4862 10492
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 8496 10520 8524 10628
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 9079 10560 9137 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9232 10588 9260 10628
rect 9232 10560 9536 10588
rect 9125 10551 9183 10557
rect 9306 10520 9312 10532
rect 5552 10492 8524 10520
rect 8864 10492 9312 10520
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2924 10424 2973 10452
rect 2924 10412 2930 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 3752 10424 3797 10452
rect 3752 10412 3758 10424
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 5552 10452 5580 10492
rect 4120 10424 5580 10452
rect 5997 10455 6055 10461
rect 4120 10412 4126 10424
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6086 10452 6092 10464
rect 6043 10424 6092 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 8864 10461 8892 10492
rect 9306 10480 9312 10492
rect 9364 10529 9370 10532
rect 9364 10523 9428 10529
rect 9364 10489 9382 10523
rect 9416 10489 9428 10523
rect 9508 10520 9536 10560
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10962 10588 10968 10600
rect 9732 10560 10968 10588
rect 9732 10548 9738 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 11112 10560 19257 10588
rect 11112 10548 11118 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 12526 10520 12532 10532
rect 9508 10492 12532 10520
rect 9364 10483 9428 10489
rect 9364 10480 9370 10483
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10468 10424 10517 10452
rect 10468 10412 10474 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 20162 10452 20168 10464
rect 19475 10424 20168 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2498 10248 2504 10260
rect 2087 10220 2504 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4430 10248 4436 10260
rect 4120 10220 4436 10248
rect 4120 10208 4126 10220
rect 4430 10208 4436 10220
rect 4488 10248 4494 10260
rect 5074 10248 5080 10260
rect 4488 10220 5080 10248
rect 4488 10208 4494 10220
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5718 10248 5724 10260
rect 5679 10220 5724 10248
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6328 10220 6837 10248
rect 6328 10208 6334 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 6825 10211 6883 10217
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 7064 10220 7205 10248
rect 7064 10208 7070 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 8386 10248 8392 10260
rect 7331 10220 8392 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9030 10248 9036 10260
rect 8619 10220 9036 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11020 10220 11805 10248
rect 11020 10208 11026 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 3326 10180 3332 10192
rect 3287 10152 3332 10180
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 4246 10140 4252 10192
rect 4304 10189 4310 10192
rect 4304 10183 4368 10189
rect 4304 10149 4322 10183
rect 4356 10180 4368 10183
rect 4356 10152 6224 10180
rect 4356 10149 4368 10152
rect 4304 10143 4368 10149
rect 4304 10140 4310 10143
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 2958 10112 2964 10124
rect 2547 10084 2964 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10112 3111 10115
rect 4154 10112 4160 10124
rect 3099 10084 4160 10112
rect 3099 10081 3111 10084
rect 3053 10075 3111 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 6196 10112 6224 10152
rect 8941 10115 8999 10121
rect 6196 10084 6316 10112
rect 2682 10044 2688 10056
rect 2643 10016 2688 10044
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 6288 10053 6316 10084
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8987 10084 9689 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10594 10112 10600 10124
rect 10551 10084 10600 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6196 9976 6224 10007
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7098 10044 7104 10056
rect 6880 10016 7104 10044
rect 6880 10004 6886 10016
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7558 10044 7564 10056
rect 7515 10016 7564 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 9030 10044 9036 10056
rect 8991 10016 9036 10044
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 10410 10044 10416 10056
rect 9263 10016 10416 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 7006 9976 7012 9988
rect 6196 9948 7012 9976
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 10042 9908 10048 9920
rect 3568 9880 10048 9908
rect 3568 9868 3574 9880
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3421 9707 3479 9713
rect 3421 9673 3433 9707
rect 3467 9704 3479 9707
rect 3694 9704 3700 9716
rect 3467 9676 3700 9704
rect 3467 9673 3479 9676
rect 3421 9667 3479 9673
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9030 9704 9036 9716
rect 8803 9676 9036 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 3142 9636 3148 9648
rect 3055 9608 3148 9636
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 4706 9636 4712 9648
rect 4571 9608 4712 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 5258 9636 5264 9648
rect 4948 9608 5264 9636
rect 4948 9596 4954 9608
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 5534 9636 5540 9648
rect 5495 9608 5540 9636
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 3160 9568 3188 9596
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3160 9540 3985 9568
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4304 9540 5089 9568
rect 4304 9528 4310 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 6089 9571 6147 9577
rect 6089 9568 6101 9571
rect 5684 9540 6101 9568
rect 5684 9528 5690 9540
rect 6089 9537 6101 9540
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 6328 9540 7757 9568
rect 6328 9528 6334 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 7745 9531 7803 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 1811 9472 1992 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 1964 9364 1992 9472
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 3844 9472 4905 9500
rect 3844 9460 3850 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 2032 9435 2090 9441
rect 2032 9401 2044 9435
rect 2078 9432 2090 9435
rect 2682 9432 2688 9444
rect 2078 9404 2688 9432
rect 2078 9401 2090 9404
rect 2032 9395 2090 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 3804 9404 5488 9432
rect 2222 9364 2228 9376
rect 1964 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 3804 9373 3832 9404
rect 5460 9376 5488 9404
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 5776 9404 6009 9432
rect 5776 9392 5782 9404
rect 5997 9401 6009 9404
rect 6043 9401 6055 9435
rect 9125 9435 9183 9441
rect 9125 9432 9137 9435
rect 5997 9395 6055 9401
rect 6104 9404 9137 9432
rect 3789 9367 3847 9373
rect 3789 9333 3801 9367
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 3881 9367 3939 9373
rect 3881 9333 3893 9367
rect 3927 9364 3939 9367
rect 4798 9364 4804 9376
rect 3927 9336 4804 9364
rect 3927 9333 3939 9336
rect 3881 9327 3939 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5166 9364 5172 9376
rect 5031 9336 5172 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5500 9336 5917 9364
rect 5500 9324 5506 9336
rect 5905 9333 5917 9336
rect 5951 9364 5963 9367
rect 6104 9364 6132 9404
rect 9125 9401 9137 9404
rect 9171 9401 9183 9435
rect 9125 9395 9183 9401
rect 7190 9364 7196 9376
rect 5951 9336 6132 9364
rect 7151 9336 7196 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7558 9364 7564 9376
rect 7519 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 9217 9367 9275 9373
rect 7708 9336 7753 9364
rect 7708 9324 7714 9336
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 9398 9364 9404 9376
rect 9263 9336 9404 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2406 9160 2412 9172
rect 1995 9132 2412 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4212 9132 4261 9160
rect 4212 9120 4218 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 7190 9160 7196 9172
rect 4755 9132 7196 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 7616 9132 8585 9160
rect 7616 9120 7622 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8720 9132 9045 9160
rect 8720 9120 8726 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 4062 9092 4068 9104
rect 2363 9064 4068 9092
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5258 9092 5264 9104
rect 5132 9064 5264 9092
rect 5132 9052 5138 9064
rect 5258 9052 5264 9064
rect 5316 9092 5322 9104
rect 5316 9064 6960 9092
rect 5316 9052 5322 9064
rect 3326 9024 3332 9036
rect 3287 8996 3332 9024
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 9024 4675 9027
rect 5350 9024 5356 9036
rect 4663 8996 5356 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5528 9027 5586 9033
rect 5528 8993 5540 9027
rect 5574 9024 5586 9027
rect 6270 9024 6276 9036
rect 5574 8996 6276 9024
rect 5574 8993 5586 8996
rect 5528 8987 5586 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 6932 9033 6960 9064
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 8260 9064 8953 9092
rect 8260 9052 8266 9064
rect 8941 9061 8953 9064
rect 8987 9061 8999 9095
rect 8941 9055 8999 9061
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 7184 9027 7242 9033
rect 7184 8993 7196 9027
rect 7230 9024 7242 9027
rect 9677 9027 9735 9033
rect 7230 8996 8524 9024
rect 7230 8993 7242 8996
rect 7184 8987 7242 8993
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 2004 8928 2421 8956
rect 2004 8916 2010 8928
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 2593 8919 2651 8925
rect 2608 8888 2636 8919
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 3694 8956 3700 8968
rect 3651 8928 3700 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 3620 8888 3648 8919
rect 3694 8916 3700 8928
rect 3752 8916 3758 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 4939 8928 5212 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 2608 8860 3648 8888
rect 5184 8820 5212 8928
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5316 8928 5361 8956
rect 5316 8916 5322 8928
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 6328 8860 6960 8888
rect 6328 8848 6334 8860
rect 5258 8820 5264 8832
rect 5171 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8820 5322 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 5316 8792 6653 8820
rect 5316 8780 5322 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6932 8820 6960 8860
rect 8496 8832 8524 8996
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 9944 9027 10002 9033
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 10318 9024 10324 9036
rect 9990 8996 10324 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9263 8928 9352 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 6932 8792 8309 8820
rect 6641 8783 6699 8789
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 8297 8783 8355 8789
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 9324 8820 9352 8928
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 12710 8888 12716 8900
rect 10744 8860 12716 8888
rect 10744 8848 10750 8860
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 10778 8820 10784 8832
rect 8536 8792 10784 8820
rect 8536 8780 8542 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 2777 8619 2835 8625
rect 2777 8616 2789 8619
rect 2740 8588 2789 8616
rect 2740 8576 2746 8588
rect 2777 8585 2789 8588
rect 2823 8585 2835 8619
rect 3694 8616 3700 8628
rect 2777 8579 2835 8585
rect 2976 8588 3700 8616
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 2976 8412 3004 8588
rect 3694 8576 3700 8588
rect 3752 8616 3758 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 3752 8588 4445 8616
rect 3752 8576 3758 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5408 8588 5733 8616
rect 5408 8576 5414 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 7374 8616 7380 8628
rect 7248 8588 7380 8616
rect 7248 8576 7254 8588
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 7708 8588 7849 8616
rect 7708 8576 7714 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 10686 8616 10692 8628
rect 7837 8579 7895 8585
rect 8312 8588 10692 8616
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 7098 8548 7104 8560
rect 4304 8520 7104 8548
rect 4304 8508 4310 8520
rect 7098 8508 7104 8520
rect 7156 8548 7162 8560
rect 7156 8520 7328 8548
rect 7156 8508 7162 8520
rect 6270 8480 6276 8492
rect 6231 8452 6276 8480
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 7300 8489 7328 8520
rect 8312 8489 8340 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 10836 8588 11161 8616
rect 10836 8576 10842 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8449 8355 8483
rect 8478 8480 8484 8492
rect 8439 8452 8484 8480
rect 8297 8443 8355 8449
rect 1710 8384 3004 8412
rect 3053 8415 3111 8421
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 4706 8412 4712 8424
rect 3099 8384 4712 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 1412 8344 1440 8375
rect 2222 8344 2228 8356
rect 1412 8316 2228 8344
rect 2222 8304 2228 8316
rect 2280 8344 2286 8356
rect 3068 8344 3096 8375
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 7374 8412 7380 8424
rect 5675 8384 7380 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7484 8412 7512 8443
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 8496 8412 8524 8440
rect 9674 8412 9680 8424
rect 7484 8384 8524 8412
rect 9635 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 2280 8316 3096 8344
rect 3320 8347 3378 8353
rect 2280 8304 2286 8316
rect 3320 8313 3332 8347
rect 3366 8344 3378 8347
rect 3602 8344 3608 8356
rect 3366 8316 3608 8344
rect 3366 8313 3378 8316
rect 3320 8307 3378 8313
rect 3602 8304 3608 8316
rect 3660 8304 3666 8356
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 3844 8316 8217 8344
rect 3844 8304 3850 8316
rect 8205 8313 8217 8316
rect 8251 8344 8263 8347
rect 8754 8344 8760 8356
rect 8251 8316 8760 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 10036 8347 10094 8353
rect 10036 8313 10048 8347
rect 10082 8344 10094 8347
rect 11054 8344 11060 8356
rect 10082 8316 11060 8344
rect 10082 8313 10094 8316
rect 10036 8307 10094 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5074 8276 5080 8288
rect 4764 8248 5080 8276
rect 4764 8236 4770 8248
rect 5074 8236 5080 8248
rect 5132 8276 5138 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5132 8248 5457 8276
rect 5132 8236 5138 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 6086 8276 6092 8288
rect 6047 8248 6092 8276
rect 5445 8239 5503 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6181 8279 6239 8285
rect 6181 8245 6193 8279
rect 6227 8276 6239 8279
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6227 8248 6837 8276
rect 6227 8245 6239 8248
rect 6181 8239 6239 8245
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 7064 8248 7205 8276
rect 7064 8236 7070 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 9490 8276 9496 8288
rect 9451 8248 9496 8276
rect 7193 8239 7251 8245
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 11422 8276 11428 8288
rect 11383 8248 11428 8276
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2188 8044 2329 8072
rect 2188 8032 2194 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3326 8072 3332 8084
rect 3007 8044 3332 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 4062 8072 4068 8084
rect 4023 8044 4068 8072
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5810 8072 5816 8084
rect 5092 8044 5816 8072
rect 5092 8004 5120 8044
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6144 8044 6653 8072
rect 6144 8032 6150 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7282 8072 7288 8084
rect 6972 8044 7288 8072
rect 6972 8032 6978 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 7432 8044 8585 8072
rect 7432 8032 7438 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 8573 8035 8631 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11422 8072 11428 8084
rect 11103 8044 11428 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 11563 8044 13645 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 5258 8013 5264 8016
rect 5252 8004 5264 8013
rect 3436 7976 5120 8004
rect 5219 7976 5264 8004
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 3326 7936 3332 7948
rect 2004 7908 3332 7936
rect 2004 7896 2010 7908
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 1912 7840 2421 7868
rect 1912 7828 1918 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2424 7732 2452 7831
rect 2608 7800 2636 7831
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3436 7877 3464 7976
rect 5252 7967 5264 7976
rect 5258 7964 5264 7967
rect 5316 7964 5322 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7392 8004 7420 8032
rect 9490 8004 9496 8016
rect 7248 7976 7420 8004
rect 8772 7976 9496 8004
rect 7248 7964 7254 7976
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4764 7908 4997 7936
rect 4764 7896 4770 7908
rect 4985 7905 4997 7908
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 8772 7945 8800 7976
rect 9490 7964 9496 7976
rect 9548 8004 9554 8016
rect 9548 7976 11928 8004
rect 9548 7964 9554 7976
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 6972 7908 7941 7936
rect 6972 7896 6978 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10226 7936 10232 7948
rect 10183 7908 10232 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11900 7945 11928 7976
rect 11992 7976 18000 8004
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10551 7908 11161 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11149 7899 11207 7905
rect 11256 7908 11529 7936
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 2832 7840 3433 7868
rect 2832 7828 2838 7840
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3421 7831 3479 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 6880 7840 8033 7868
rect 6880 7828 6886 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8478 7868 8484 7880
rect 8251 7840 8484 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 10318 7868 10324 7880
rect 10231 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7868 10382 7880
rect 11256 7868 11284 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 10376 7840 11284 7868
rect 11333 7871 11391 7877
rect 10376 7828 10382 7840
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11992 7868 12020 7976
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7936 12311 7939
rect 12342 7936 12348 7948
rect 12299 7908 12348 7936
rect 12299 7905 12311 7908
rect 12253 7899 12311 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12520 7939 12578 7945
rect 12520 7905 12532 7939
rect 12566 7936 12578 7939
rect 13814 7936 13820 7948
rect 12566 7908 13820 7936
rect 12566 7905 12578 7908
rect 12520 7899 12578 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 17972 7945 18000 7976
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 11333 7831 11391 7837
rect 11532 7840 12020 7868
rect 18233 7871 18291 7877
rect 3620 7800 3648 7828
rect 2608 7772 3648 7800
rect 7561 7803 7619 7809
rect 7561 7769 7573 7803
rect 7607 7800 7619 7803
rect 9677 7803 9735 7809
rect 7607 7772 9628 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 4246 7732 4252 7744
rect 2424 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 6365 7735 6423 7741
rect 6365 7732 6377 7735
rect 4764 7704 6377 7732
rect 4764 7692 4770 7704
rect 6365 7701 6377 7704
rect 6411 7701 6423 7735
rect 9600 7732 9628 7772
rect 9677 7769 9689 7803
rect 9723 7800 9735 7803
rect 10505 7803 10563 7809
rect 10505 7800 10517 7803
rect 9723 7772 10517 7800
rect 9723 7769 9735 7772
rect 9677 7763 9735 7769
rect 10505 7769 10517 7772
rect 10551 7769 10563 7803
rect 10505 7763 10563 7769
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11348 7800 11376 7831
rect 11112 7772 11376 7800
rect 11112 7760 11118 7772
rect 9950 7732 9956 7744
rect 9600 7704 9956 7732
rect 6365 7695 6423 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7732 10747 7735
rect 11532 7732 11560 7840
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18690 7868 18696 7880
rect 18279 7840 18696 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 10735 7704 11560 7732
rect 11701 7735 11759 7741
rect 10735 7701 10747 7704
rect 10689 7695 10747 7701
rect 11701 7701 11713 7735
rect 11747 7732 11759 7735
rect 11974 7732 11980 7744
rect 11747 7704 11980 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 3605 7531 3663 7537
rect 3605 7528 3617 7531
rect 3476 7500 3617 7528
rect 3476 7488 3482 7500
rect 3605 7497 3617 7500
rect 3651 7497 3663 7531
rect 3605 7491 3663 7497
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 7742 7528 7748 7540
rect 3936 7500 7748 7528
rect 3936 7488 3942 7500
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 13814 7528 13820 7540
rect 8435 7500 13676 7528
rect 13775 7500 13820 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3660 7364 4169 7392
rect 3660 7352 3666 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7708 7364 7941 7392
rect 7708 7352 7714 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 8938 7392 8944 7404
rect 8899 7364 8944 7392
rect 7929 7355 7987 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3844 7296 3985 7324
rect 3844 7284 3850 7296
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 5074 7324 5080 7336
rect 5035 7296 5080 7324
rect 3973 7287 4031 7293
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7524 7296 7849 7324
rect 7524 7284 7530 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 8444 7296 9597 7324
rect 8444 7284 8450 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9852 7327 9910 7333
rect 9852 7293 9864 7327
rect 9898 7324 9910 7327
rect 10686 7324 10692 7336
rect 9898 7296 10692 7324
rect 9898 7293 9910 7296
rect 9852 7287 9910 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12704 7327 12762 7333
rect 12704 7293 12716 7327
rect 12750 7324 12762 7327
rect 13648 7324 13676 7500
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7460 14151 7463
rect 16482 7460 16488 7472
rect 14139 7432 16488 7460
rect 14139 7429 14151 7432
rect 14093 7423 14151 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 13872 7364 14657 7392
rect 13872 7352 13878 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 16574 7324 16580 7336
rect 12750 7296 12848 7324
rect 13648 7296 16580 7324
rect 12750 7293 12762 7296
rect 12704 7287 12762 7293
rect 12820 7268 12848 7296
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 5344 7259 5402 7265
rect 5344 7225 5356 7259
rect 5390 7256 5402 7259
rect 5902 7256 5908 7268
rect 5390 7228 5908 7256
rect 5390 7225 5402 7228
rect 5344 7219 5402 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 7392 7228 8861 7256
rect 1486 7148 1492 7200
rect 1544 7188 1550 7200
rect 1949 7191 2007 7197
rect 1949 7188 1961 7191
rect 1544 7160 1961 7188
rect 1544 7148 1550 7160
rect 1949 7157 1961 7160
rect 1995 7157 2007 7191
rect 2314 7188 2320 7200
rect 2275 7160 2320 7188
rect 1949 7151 2007 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2774 7188 2780 7200
rect 2455 7160 2780 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4062 7188 4068 7200
rect 4023 7160 4068 7188
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 6454 7188 6460 7200
rect 6415 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7392 7197 7420 7228
rect 8849 7225 8861 7228
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 12618 7256 12624 7268
rect 10008 7228 12624 7256
rect 10008 7216 10014 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 12802 7216 12808 7268
rect 12860 7216 12866 7268
rect 12986 7216 12992 7268
rect 13044 7256 13050 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 13044 7228 14565 7256
rect 13044 7216 13050 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7157 7435 7191
rect 7742 7188 7748 7200
rect 7703 7160 7748 7188
rect 7377 7151 7435 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8754 7188 8760 7200
rect 8715 7160 8760 7188
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 10962 7188 10968 7200
rect 10923 7160 10968 7188
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 11112 7160 11253 7188
rect 11112 7148 11118 7160
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 11885 7191 11943 7197
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 11931 7160 14473 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 14461 7157 14473 7160
rect 14507 7157 14519 7191
rect 14461 7151 14519 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3602 6984 3608 6996
rect 3563 6956 3608 6984
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 5626 6984 5632 6996
rect 4028 6956 5632 6984
rect 4028 6944 4034 6956
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 1762 6876 1768 6928
rect 1820 6916 1826 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 1820 6888 4445 6916
rect 1820 6876 1826 6888
rect 4433 6885 4445 6888
rect 4479 6916 4491 6919
rect 5534 6916 5540 6928
rect 4479 6888 5540 6916
rect 4479 6885 4491 6888
rect 4433 6879 4491 6885
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 5988 6919 6046 6925
rect 5988 6885 6000 6919
rect 6034 6916 6046 6919
rect 6454 6916 6460 6928
rect 6034 6888 6460 6916
rect 6034 6885 6046 6888
rect 5988 6879 6046 6885
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 7116 6916 7144 6947
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8812 6956 9045 6984
rect 8812 6944 8818 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 10502 6984 10508 6996
rect 9033 6947 9091 6953
rect 9784 6956 10508 6984
rect 7650 6925 7656 6928
rect 7644 6916 7656 6925
rect 7116 6888 7656 6916
rect 7644 6879 7656 6888
rect 7650 6876 7656 6879
rect 7708 6876 7714 6928
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 2498 6857 2504 6860
rect 2492 6848 2504 6857
rect 2459 6820 2504 6848
rect 2492 6811 2504 6820
rect 2498 6808 2504 6811
rect 2556 6808 2562 6860
rect 4890 6848 4896 6860
rect 4540 6820 4896 6848
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 4540 6789 4568 6820
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5132 6820 5733 6848
rect 5132 6808 5138 6820
rect 5721 6817 5733 6820
rect 5767 6848 5779 6851
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 5767 6820 7389 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9784 6848 9812 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 13096 6956 16681 6984
rect 10404 6919 10462 6925
rect 10404 6885 10416 6919
rect 10450 6916 10462 6919
rect 10962 6916 10968 6928
rect 10450 6888 10968 6916
rect 10450 6885 10462 6888
rect 10404 6879 10462 6885
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 12802 6916 12808 6928
rect 12715 6888 12808 6916
rect 12802 6876 12808 6888
rect 12860 6916 12866 6928
rect 13096 6916 13124 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 16669 6947 16727 6953
rect 12860 6888 13124 6916
rect 12860 6876 12866 6888
rect 8260 6820 9812 6848
rect 8260 6808 8266 6820
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3252 6752 4537 6780
rect 3252 6712 3280 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4525 6743 4583 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 9950 6780 9956 6792
rect 9824 6752 9956 6780
rect 9824 6740 9830 6752
rect 9950 6740 9956 6752
rect 10008 6780 10014 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10008 6752 10149 6780
rect 10008 6740 10014 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 12820 6789 12848 6876
rect 13440 6851 13498 6857
rect 13440 6817 13452 6851
rect 13486 6848 13498 6851
rect 13814 6848 13820 6860
rect 13486 6820 13820 6848
rect 13486 6817 13498 6820
rect 13440 6811 13498 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 15556 6851 15614 6857
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 16114 6848 16120 6860
rect 15602 6820 16120 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16540 6820 17417 6848
rect 16540 6808 16546 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 11848 6752 12633 6780
rect 11848 6740 11854 6752
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 12805 6743 12863 6749
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 14366 6740 14372 6792
rect 14424 6780 14430 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 14424 6752 15301 6780
rect 14424 6740 14430 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 17678 6780 17684 6792
rect 17639 6752 17684 6780
rect 15289 6743 15347 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 3160 6684 3280 6712
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 3160 6644 3188 6684
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3384 6684 4077 6712
rect 3384 6672 3390 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 8938 6712 8944 6724
rect 8803 6684 8944 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 12161 6715 12219 6721
rect 12161 6681 12173 6715
rect 12207 6712 12219 6715
rect 12986 6712 12992 6724
rect 12207 6684 12992 6712
rect 12207 6681 12219 6684
rect 12161 6675 12219 6681
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 1544 6616 3188 6644
rect 1544 6604 1550 6616
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 4890 6644 4896 6656
rect 3292 6616 4896 6644
rect 3292 6604 3298 6616
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5902 6604 5908 6656
rect 5960 6644 5966 6656
rect 11517 6647 11575 6653
rect 11517 6644 11529 6647
rect 5960 6616 11529 6644
rect 5960 6604 5966 6616
rect 11517 6613 11529 6616
rect 11563 6613 11575 6647
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 11517 6607 11575 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2556 6412 2789 6440
rect 2556 6400 2562 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 12434 6440 12440 6452
rect 4948 6412 12440 6440
rect 4948 6400 4954 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 6914 6372 6920 6384
rect 6871 6344 6920 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 11238 6372 11244 6384
rect 10008 6344 11244 6372
rect 10008 6332 10014 6344
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 11333 6375 11391 6381
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 11379 6344 12480 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 5902 6304 5908 6316
rect 5863 6276 5908 6304
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7064 6276 7389 6304
rect 7064 6264 7070 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 8386 6304 8392 6316
rect 8347 6276 8392 6304
rect 7377 6267 7435 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 10686 6304 10692 6316
rect 10647 6276 10692 6304
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 12452 6304 12480 6344
rect 13832 6304 13860 6400
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 12452 6276 12572 6304
rect 13832 6276 14657 6304
rect 11977 6267 12035 6273
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 2280 6208 3433 6236
rect 2280 6196 2286 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 4028 6208 7297 6236
rect 4028 6196 4034 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8656 6239 8714 6245
rect 8656 6205 8668 6239
rect 8702 6236 8714 6239
rect 8938 6236 8944 6248
rect 8702 6208 8944 6236
rect 8702 6205 8714 6208
rect 8656 6199 8714 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9180 6208 10425 6236
rect 9180 6196 9186 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 11790 6236 11796 6248
rect 10560 6208 11796 6236
rect 10560 6196 10566 6208
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 1664 6171 1722 6177
rect 1664 6137 1676 6171
rect 1710 6168 1722 6171
rect 3688 6171 3746 6177
rect 1710 6140 3464 6168
rect 1710 6137 1722 6140
rect 1664 6131 1722 6137
rect 2498 6060 2504 6112
rect 2556 6100 2562 6112
rect 2866 6100 2872 6112
rect 2556 6072 2872 6100
rect 2556 6060 2562 6072
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3436 6100 3464 6140
rect 3688 6137 3700 6171
rect 3734 6168 3746 6171
rect 4706 6168 4712 6180
rect 3734 6140 4712 6168
rect 3734 6137 3746 6140
rect 3688 6131 3746 6137
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 5626 6168 5632 6180
rect 5587 6140 5632 6168
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 7193 6171 7251 6177
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 7742 6168 7748 6180
rect 7239 6140 7748 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 11701 6171 11759 6177
rect 11701 6168 11713 6171
rect 7892 6140 11713 6168
rect 7892 6128 7898 6140
rect 11701 6137 11713 6140
rect 11747 6137 11759 6171
rect 11992 6168 12020 6267
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12342 6236 12348 6248
rect 12299 6208 12348 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12400 6208 12449 6236
rect 12400 6196 12406 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12544 6236 12572 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 12544 6208 14565 6236
rect 12437 6199 12495 6205
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 15102 6236 15108 6248
rect 15063 6208 15108 6236
rect 14553 6199 14611 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 15838 6236 15844 6248
rect 15799 6208 15844 6236
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 16574 6236 16580 6248
rect 16535 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 17736 6208 18337 6236
rect 17736 6196 17742 6208
rect 18325 6205 18337 6208
rect 18371 6205 18383 6239
rect 18325 6199 18383 6205
rect 12682 6171 12740 6177
rect 12682 6168 12694 6171
rect 11992 6140 12694 6168
rect 11701 6131 11759 6137
rect 12682 6137 12694 6140
rect 12728 6168 12740 6171
rect 12802 6168 12808 6180
rect 12728 6140 12808 6168
rect 12728 6137 12740 6140
rect 12682 6131 12740 6137
rect 12802 6128 12808 6140
rect 12860 6128 12866 6180
rect 15381 6171 15439 6177
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 16022 6168 16028 6180
rect 15427 6140 16028 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 16117 6171 16175 6177
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16298 6168 16304 6180
rect 16163 6140 16304 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16298 6128 16304 6140
rect 16356 6128 16362 6180
rect 16850 6168 16856 6180
rect 16811 6140 16856 6168
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 3786 6100 3792 6112
rect 3436 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6100 3850 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 3844 6072 4813 6100
rect 3844 6060 3850 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 4801 6063 4859 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6144 6072 6285 6100
rect 6144 6060 6150 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 6273 6063 6331 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10045 6103 10103 6109
rect 10045 6069 10057 6103
rect 10091 6100 10103 6103
rect 10134 6100 10140 6112
rect 10091 6072 10140 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 10284 6072 10517 6100
rect 10284 6060 10290 6072
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 10505 6063 10563 6069
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 13170 6100 13176 6112
rect 12299 6072 13176 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 13964 6072 14105 6100
rect 13964 6060 13970 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 14458 6100 14464 6112
rect 14419 6072 14464 6100
rect 14093 6063 14151 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 19242 6100 19248 6112
rect 18555 6072 19248 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2314 5896 2320 5908
rect 1995 5868 2320 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2832 5868 2973 5896
rect 2832 5856 2838 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 3326 5896 3332 5908
rect 3287 5868 3332 5896
rect 2961 5859 3019 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3467 5868 4077 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 5350 5896 5356 5908
rect 4479 5868 5356 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 8478 5896 8484 5908
rect 6288 5868 7512 5896
rect 8439 5868 8484 5896
rect 3878 5788 3884 5840
rect 3936 5828 3942 5840
rect 3936 5800 4568 5828
rect 3936 5788 3942 5800
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2958 5760 2964 5772
rect 2363 5732 2964 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 4540 5760 4568 5800
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 6181 5831 6239 5837
rect 6181 5828 6193 5831
rect 5316 5800 6193 5828
rect 5316 5788 5322 5800
rect 6181 5797 6193 5800
rect 6227 5797 6239 5831
rect 6181 5791 6239 5797
rect 6288 5760 6316 5868
rect 7190 5828 7196 5840
rect 6932 5800 7196 5828
rect 6932 5769 6960 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 7484 5828 7512 5868
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 11054 5896 11060 5908
rect 10735 5868 11060 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 14458 5896 14464 5908
rect 13679 5868 14464 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 10152 5828 10180 5856
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 7484 5800 8156 5828
rect 10152 5800 10793 5828
rect 4540 5732 6316 5760
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 7357 5763 7415 5769
rect 7357 5760 7369 5763
rect 7064 5732 7369 5760
rect 7064 5720 7070 5732
rect 7357 5729 7369 5732
rect 7403 5729 7415 5763
rect 7357 5723 7415 5729
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 2639 5664 3617 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3605 5661 3617 5664
rect 3651 5692 3663 5695
rect 3786 5692 3792 5704
rect 3651 5664 3792 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4212 5664 4537 5692
rect 4212 5652 4218 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4525 5655 4583 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6454 5692 6460 5704
rect 6411 5664 6460 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6687 5664 7113 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 8128 5692 8156 5800
rect 10781 5797 10793 5800
rect 10827 5797 10839 5831
rect 11692 5831 11750 5837
rect 10781 5791 10839 5797
rect 11072 5800 11652 5828
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 11072 5760 11100 5800
rect 10183 5732 11100 5760
rect 11624 5760 11652 5800
rect 11692 5797 11704 5831
rect 11738 5828 11750 5831
rect 11790 5828 11796 5840
rect 11738 5800 11796 5828
rect 11738 5797 11750 5800
rect 11692 5791 11750 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 15657 5831 15715 5837
rect 15657 5797 15669 5831
rect 15703 5828 15715 5831
rect 16574 5828 16580 5840
rect 15703 5800 16580 5828
rect 15703 5797 15715 5800
rect 15657 5791 15715 5797
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 11974 5760 11980 5772
rect 11624 5732 11980 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 11974 5720 11980 5732
rect 12032 5760 12038 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 12032 5732 13277 5760
rect 12032 5720 12038 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 15749 5763 15807 5769
rect 15749 5760 15761 5763
rect 13265 5723 13323 5729
rect 13464 5732 15761 5760
rect 10778 5692 10784 5704
rect 8128 5664 10784 5692
rect 7101 5655 7159 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10962 5692 10968 5704
rect 10923 5664 10968 5692
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 11296 5664 11437 5692
rect 11296 5652 11302 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13464 5692 13492 5732
rect 15749 5729 15761 5732
rect 15795 5729 15807 5763
rect 16298 5760 16304 5772
rect 16259 5732 16304 5760
rect 15749 5723 15807 5729
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16850 5760 16856 5772
rect 16811 5732 16856 5760
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 15838 5692 15844 5704
rect 12492 5664 13492 5692
rect 15799 5664 15844 5692
rect 12492 5652 12498 5664
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 5721 5627 5779 5633
rect 5721 5593 5733 5627
rect 5767 5624 5779 5627
rect 15102 5624 15108 5636
rect 5767 5596 7144 5624
rect 5767 5593 5779 5596
rect 5721 5587 5779 5593
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 5684 5528 6653 5556
rect 5684 5516 5690 5528
rect 6641 5525 6653 5528
rect 6687 5556 6699 5559
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6687 5528 6745 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6733 5525 6745 5528
rect 6779 5556 6791 5559
rect 6914 5556 6920 5568
rect 6779 5528 6920 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7116 5556 7144 5596
rect 12728 5596 15108 5624
rect 10134 5556 10140 5568
rect 7116 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 12728 5556 12756 5596
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 10367 5528 12756 5556
rect 13081 5559 13139 5565
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13170 5556 13176 5568
rect 13127 5528 13176 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13170 5516 13176 5528
rect 13228 5556 13234 5568
rect 14366 5556 14372 5568
rect 13228 5528 14372 5556
rect 13228 5516 13234 5528
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 16482 5556 16488 5568
rect 16443 5528 16488 5556
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 16942 5516 16948 5568
rect 17000 5556 17006 5568
rect 17037 5559 17095 5565
rect 17037 5556 17049 5559
rect 17000 5528 17049 5556
rect 17000 5516 17006 5528
rect 17037 5525 17049 5528
rect 17083 5525 17095 5559
rect 17037 5519 17095 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 11790 5352 11796 5364
rect 2639 5324 11468 5352
rect 11751 5324 11796 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 4617 5287 4675 5293
rect 4617 5253 4629 5287
rect 4663 5284 4675 5287
rect 6454 5284 6460 5296
rect 4663 5256 6460 5284
rect 4663 5253 4675 5256
rect 4617 5247 4675 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6822 5284 6828 5296
rect 6783 5256 6828 5284
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 7190 5284 7196 5296
rect 6972 5256 7196 5284
rect 6972 5244 6978 5256
rect 7190 5244 7196 5256
rect 7248 5284 7254 5296
rect 7248 5256 8432 5284
rect 7248 5244 7254 5256
rect 8404 5228 8432 5256
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2866 5216 2872 5228
rect 2271 5188 2872 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 3142 5216 3148 5228
rect 3103 5188 3148 5216
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4764 5188 5181 5216
rect 4764 5176 4770 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 6362 5216 6368 5228
rect 6323 5188 6368 5216
rect 5169 5179 5227 5185
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7064 5188 7389 5216
rect 7064 5176 7070 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7800 5188 7849 5216
rect 7800 5176 7806 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8444 5188 8769 5216
rect 8444 5176 8450 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10008 5188 10425 5216
rect 10008 5176 10014 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 11440 5216 11468 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 13078 5352 13084 5364
rect 12676 5324 13084 5352
rect 12676 5312 12682 5324
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16172 5324 16313 5352
rect 16172 5312 16178 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 11756 5256 13124 5284
rect 11756 5244 11762 5256
rect 11974 5216 11980 5228
rect 11440 5188 11980 5216
rect 10413 5179 10471 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 13096 5225 13124 5256
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 16574 5216 16580 5228
rect 13081 5179 13139 5185
rect 13740 5188 15056 5216
rect 16535 5188 16580 5216
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5148 2007 5151
rect 3326 5148 3332 5160
rect 1995 5120 3332 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 5810 5148 5816 5160
rect 3844 5120 5816 5148
rect 3844 5108 3850 5120
rect 5810 5108 5816 5120
rect 5868 5148 5874 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5868 5120 6101 5148
rect 5868 5108 5874 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6880 5120 7205 5148
rect 6880 5108 6886 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 12584 5120 12817 5148
rect 12584 5108 12590 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13740 5148 13768 5188
rect 13906 5148 13912 5160
rect 12943 5120 13768 5148
rect 13867 5120 13912 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 2961 5083 3019 5089
rect 2961 5080 2973 5083
rect 1596 5052 2973 5080
rect 1596 5021 1624 5052
rect 2961 5049 2973 5052
rect 3007 5049 3019 5083
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 2961 5043 3019 5049
rect 5736 5052 7297 5080
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 4981 1639 5015
rect 1581 4975 1639 4981
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2096 4984 2141 5012
rect 2096 4972 2102 4984
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2372 4984 3065 5012
rect 2372 4972 2378 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 3053 4975 3111 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 5736 5021 5764 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 9002 5083 9060 5089
rect 9002 5080 9014 5083
rect 8536 5052 9014 5080
rect 8536 5040 8542 5052
rect 9002 5049 9014 5052
rect 9048 5049 9060 5083
rect 9002 5043 9060 5049
rect 10680 5083 10738 5089
rect 10680 5049 10692 5083
rect 10726 5049 10738 5083
rect 10680 5043 10738 5049
rect 5721 5015 5779 5021
rect 5132 4984 5177 5012
rect 5132 4972 5138 4984
rect 5721 4981 5733 5015
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6270 5012 6276 5024
rect 6227 4984 6276 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6270 4972 6276 4984
rect 6328 5012 6334 5024
rect 8202 5012 8208 5024
rect 6328 4984 8208 5012
rect 6328 4972 6334 4984
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10695 5012 10723 5043
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 12912 5080 12940 5111
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 14424 5120 14933 5148
rect 14424 5108 14430 5120
rect 14921 5117 14933 5120
rect 14967 5117 14979 5151
rect 15028 5148 15056 5188
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 16758 5148 16764 5160
rect 15028 5120 16764 5148
rect 14921 5111 14979 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 12676 5052 12940 5080
rect 14185 5083 14243 5089
rect 12676 5040 12682 5052
rect 14185 5049 14197 5083
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 15188 5083 15246 5089
rect 15188 5049 15200 5083
rect 15234 5080 15246 5083
rect 15838 5080 15844 5092
rect 15234 5052 15844 5080
rect 15234 5049 15246 5052
rect 15188 5043 15246 5049
rect 11698 5012 11704 5024
rect 10183 4984 11704 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 11940 4984 12449 5012
rect 11940 4972 11946 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 14200 5012 14228 5043
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 15470 5012 15476 5024
rect 14200 4984 15476 5012
rect 12437 4975 12495 4981
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3142 4808 3148 4820
rect 3099 4780 3148 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 5074 4808 5080 4820
rect 4111 4780 5080 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 9950 4768 9956 4820
rect 10008 4768 10014 4820
rect 11882 4808 11888 4820
rect 11843 4780 11888 4808
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 15795 4780 16313 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 4433 4743 4491 4749
rect 4433 4740 4445 4743
rect 3568 4712 4445 4740
rect 3568 4700 3574 4712
rect 4433 4709 4445 4712
rect 4479 4709 4491 4743
rect 8294 4740 8300 4752
rect 4433 4703 4491 4709
rect 4540 4712 8300 4740
rect 1940 4675 1998 4681
rect 1940 4641 1952 4675
rect 1986 4672 1998 4675
rect 2866 4672 2872 4684
rect 1986 4644 2872 4672
rect 1986 4641 1998 4644
rect 1940 4635 1998 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 3878 4672 3884 4684
rect 3384 4644 3884 4672
rect 3384 4632 3390 4644
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 1670 4604 1676 4616
rect 1452 4576 1676 4604
rect 1452 4564 1458 4576
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4540 4613 4568 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 9968 4740 9996 4768
rect 9692 4712 9996 4740
rect 13357 4743 13415 4749
rect 4890 4632 4896 4684
rect 4948 4672 4954 4684
rect 5626 4672 5632 4684
rect 4948 4644 5632 4672
rect 4948 4632 4954 4644
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 5896 4675 5954 4681
rect 5896 4641 5908 4675
rect 5942 4672 5954 4675
rect 6362 4672 6368 4684
rect 5942 4644 6368 4672
rect 5942 4641 5954 4644
rect 5896 4635 5954 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 8113 4675 8171 4681
rect 8113 4641 8125 4675
rect 8159 4672 8171 4675
rect 9122 4672 9128 4684
rect 8159 4644 9128 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9692 4681 9720 4712
rect 13357 4709 13369 4743
rect 13403 4740 13415 4743
rect 14550 4740 14556 4752
rect 13403 4712 14556 4740
rect 13403 4709 13415 4712
rect 13357 4703 13415 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9944 4675 10002 4681
rect 9944 4672 9956 4675
rect 9824 4644 9956 4672
rect 9824 4632 9830 4644
rect 9944 4641 9956 4644
rect 9990 4672 10002 4675
rect 10318 4672 10324 4684
rect 9990 4644 10324 4672
rect 9990 4641 10002 4644
rect 9944 4635 10002 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11839 4644 12449 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 12437 4635 12495 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4641 13875 4675
rect 16666 4672 16672 4684
rect 16627 4644 16672 4672
rect 13817 4635 13875 4641
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 3752 4576 4537 4604
rect 3752 4564 3758 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5534 4604 5540 4616
rect 4755 4576 5540 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8938 4604 8944 4616
rect 8435 4576 8944 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11940 4576 11989 4604
rect 11940 4564 11946 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 11425 4539 11483 4545
rect 11425 4505 11437 4539
rect 11471 4536 11483 4539
rect 13832 4536 13860 4635
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4604 14151 4607
rect 14458 4604 14464 4616
rect 14139 4576 14464 4604
rect 14139 4573 14151 4576
rect 14093 4567 14151 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16114 4604 16120 4616
rect 15979 4576 16120 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 11471 4508 13860 4536
rect 11471 4505 11483 4508
rect 11425 4499 11483 4505
rect 15838 4496 15844 4548
rect 15896 4536 15902 4548
rect 16868 4536 16896 4567
rect 15896 4508 16896 4536
rect 15896 4496 15902 4508
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 9582 4468 9588 4480
rect 7791 4440 9588 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 15289 4471 15347 4477
rect 15289 4437 15301 4471
rect 15335 4468 15347 4471
rect 17034 4468 17040 4480
rect 15335 4440 17040 4468
rect 15335 4437 15347 4440
rect 15289 4431 15347 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 2314 4264 2320 4276
rect 1719 4236 2320 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 2866 4264 2872 4276
rect 2424 4236 2872 4264
rect 2424 4196 2452 4236
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 6822 4264 6828 4276
rect 6783 4236 6828 4264
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 8202 4264 8208 4276
rect 7883 4236 8208 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 16666 4264 16672 4276
rect 8352 4236 16672 4264
rect 8352 4224 8358 4236
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 6362 4196 6368 4208
rect 2332 4168 2452 4196
rect 6275 4168 6368 4196
rect 2332 4137 2360 4168
rect 6362 4156 6368 4168
rect 6420 4196 6426 4208
rect 15838 4196 15844 4208
rect 6420 4168 7420 4196
rect 15799 4168 15844 4196
rect 6420 4156 6426 4168
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4246 4128 4252 4140
rect 4120 4100 4252 4128
rect 4120 4088 4126 4100
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4890 4128 4896 4140
rect 4488 4100 4896 4128
rect 4488 4088 4494 4100
rect 4890 4088 4896 4100
rect 4948 4128 4954 4140
rect 7392 4137 7420 4168
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4948 4100 4997 4128
rect 4948 4088 4954 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 7377 4091 7435 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8846 4128 8852 4140
rect 8527 4100 8852 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 8996 4100 9413 4128
rect 8996 4088 9002 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 13446 4128 13452 4140
rect 13407 4100 13452 4128
rect 10045 4091 10103 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 18046 4128 18052 4140
rect 15488 4100 18052 4128
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 1728 4032 2697 4060
rect 1728 4020 1734 4032
rect 2685 4029 2697 4032
rect 2731 4060 2743 4063
rect 4448 4060 4476 4088
rect 2731 4032 4476 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5132 4032 5948 4060
rect 5132 4020 5138 4032
rect 2952 3995 3010 4001
rect 2952 3961 2964 3995
rect 2998 3992 3010 3995
rect 3142 3992 3148 4004
rect 2998 3964 3148 3992
rect 2998 3961 3010 3964
rect 2952 3955 3010 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 5252 3995 5310 4001
rect 5252 3961 5264 3995
rect 5298 3992 5310 3995
rect 5810 3992 5816 4004
rect 5298 3964 5816 3992
rect 5298 3961 5310 3964
rect 5252 3955 5310 3961
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 4065 3927 4123 3933
rect 2188 3896 2233 3924
rect 2188 3884 2194 3896
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 5534 3924 5540 3936
rect 4111 3896 5540 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5920 3924 5948 4032
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6788 4032 7297 4060
rect 6788 4020 6794 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 8202 4060 8208 4072
rect 8163 4032 8208 4060
rect 7285 4023 7343 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8496 4032 10272 4060
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 5920 3896 7205 3924
rect 7193 3893 7205 3896
rect 7239 3924 7251 3927
rect 8496 3924 8524 4032
rect 9766 3992 9772 4004
rect 8864 3964 9772 3992
rect 8864 3933 8892 3964
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 7239 3896 8524 3924
rect 8849 3927 8907 3933
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 8849 3893 8861 3927
rect 8895 3893 8907 3927
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 8849 3887 8907 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9364 3896 9409 3924
rect 9364 3884 9370 3896
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10134 3924 10140 3936
rect 9732 3896 10140 3924
rect 9732 3884 9738 3896
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10244 3924 10272 4032
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 12158 4060 12164 4072
rect 10652 4032 12164 4060
rect 10652 4020 10658 4032
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12268 4032 13277 4060
rect 10312 3995 10370 4001
rect 10312 3961 10324 3995
rect 10358 3992 10370 3995
rect 11054 3992 11060 4004
rect 10358 3964 11060 3992
rect 10358 3961 10370 3964
rect 10312 3955 10370 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 12268 3992 12296 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 14366 4060 14372 4072
rect 13596 4032 14372 4060
rect 13596 4020 13602 4032
rect 14366 4020 14372 4032
rect 14424 4060 14430 4072
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 14424 4032 14473 4060
rect 14424 4020 14430 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 15488 4060 15516 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 17034 4060 17040 4072
rect 14461 4023 14519 4029
rect 14568 4032 15516 4060
rect 16995 4032 17040 4060
rect 13170 3992 13176 4004
rect 11164 3964 12296 3992
rect 13131 3964 13176 3992
rect 11164 3924 11192 3964
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14568 3992 14596 4032
rect 17034 4020 17040 4032
rect 17092 4020 17098 4072
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 19886 4069 19892 4072
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 17184 4032 19625 4060
rect 17184 4020 17190 4032
rect 19613 4029 19625 4032
rect 19659 4029 19671 4063
rect 19880 4060 19892 4069
rect 19847 4032 19892 4060
rect 19613 4023 19671 4029
rect 19880 4023 19892 4032
rect 19886 4020 19892 4023
rect 19944 4020 19950 4072
rect 13412 3964 14596 3992
rect 14728 3995 14786 4001
rect 13412 3952 13418 3964
rect 14728 3961 14740 3995
rect 14774 3992 14786 3995
rect 15010 3992 15016 4004
rect 14774 3964 15016 3992
rect 14774 3961 14786 3964
rect 14728 3955 14786 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 17313 3995 17371 4001
rect 15988 3964 16252 3992
rect 15988 3952 15994 3964
rect 10244 3896 11192 3924
rect 11425 3927 11483 3933
rect 11425 3893 11437 3927
rect 11471 3924 11483 3927
rect 11606 3924 11612 3936
rect 11471 3896 11612 3924
rect 11471 3893 11483 3896
rect 11425 3887 11483 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12805 3927 12863 3933
rect 12805 3893 12817 3927
rect 12851 3924 12863 3927
rect 15746 3924 15752 3936
rect 12851 3896 15752 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16224 3924 16252 3964
rect 17313 3961 17325 3995
rect 17359 3992 17371 3995
rect 17954 3992 17960 4004
rect 17359 3964 17960 3992
rect 17359 3961 17371 3964
rect 17313 3955 17371 3961
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 20993 3927 21051 3933
rect 20993 3924 21005 3927
rect 16224 3896 21005 3924
rect 20993 3893 21005 3896
rect 21039 3893 21051 3927
rect 20993 3887 21051 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2866 3720 2872 3732
rect 2827 3692 2872 3720
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3694 3720 3700 3732
rect 3568 3692 3700 3720
rect 3568 3680 3574 3692
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 13173 3723 13231 3729
rect 4120 3692 13124 3720
rect 4120 3680 4126 3692
rect 1670 3652 1676 3664
rect 1504 3624 1676 3652
rect 1504 3593 1532 3624
rect 1670 3612 1676 3624
rect 1728 3612 1734 3664
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 4154 3652 4160 3664
rect 2832 3624 4160 3652
rect 2832 3612 2838 3624
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 4706 3661 4712 3664
rect 4700 3652 4712 3661
rect 4667 3624 4712 3652
rect 4700 3615 4712 3624
rect 4706 3612 4712 3615
rect 4764 3612 4770 3664
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 5350 3652 5356 3664
rect 4948 3624 5356 3652
rect 4948 3612 4954 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 6454 3652 6460 3664
rect 6415 3624 6460 3652
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 7558 3652 7564 3664
rect 6604 3624 7564 3652
rect 6604 3612 6610 3624
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 9122 3652 9128 3664
rect 7668 3624 8984 3652
rect 9083 3624 9128 3652
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 1756 3587 1814 3593
rect 1756 3553 1768 3587
rect 1802 3584 1814 3587
rect 3418 3584 3424 3596
rect 1802 3556 3424 3584
rect 1802 3553 1814 3556
rect 1756 3547 1814 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 7006 3584 7012 3596
rect 4264 3556 7012 3584
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 4264 3516 4292 3556
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7374 3584 7380 3596
rect 7248 3556 7380 3584
rect 7248 3544 7254 3556
rect 7374 3544 7380 3556
rect 7432 3584 7438 3596
rect 7469 3587 7527 3593
rect 7469 3584 7481 3587
rect 7432 3556 7481 3584
rect 7432 3544 7438 3556
rect 7469 3553 7481 3556
rect 7515 3553 7527 3587
rect 7668 3584 7696 3624
rect 7469 3547 7527 3553
rect 7576 3556 7696 3584
rect 7736 3587 7794 3593
rect 4430 3516 4436 3528
rect 2556 3488 4292 3516
rect 4391 3488 4436 3516
rect 2556 3476 2562 3488
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 5500 3488 6561 3516
rect 5500 3476 5506 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 7576 3516 7604 3556
rect 7736 3553 7748 3587
rect 7782 3584 7794 3587
rect 8846 3584 8852 3596
rect 7782 3556 8852 3584
rect 7782 3553 7794 3556
rect 7736 3547 7794 3553
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 8956 3584 8984 3624
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 12066 3661 12072 3664
rect 12038 3655 12072 3661
rect 12038 3652 12050 3655
rect 10008 3624 10180 3652
rect 10008 3612 10014 3624
rect 10152 3593 10180 3624
rect 11716 3624 12050 3652
rect 10137 3587 10195 3593
rect 8956 3556 10088 3584
rect 6641 3479 6699 3485
rect 7484 3488 7604 3516
rect 8956 3516 8984 3556
rect 9122 3516 9128 3528
rect 8956 3488 9128 3516
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4448 3448 4476 3476
rect 5810 3448 5816 3460
rect 3752 3420 4476 3448
rect 5771 3420 5816 3448
rect 3752 3408 3758 3420
rect 5810 3408 5816 3420
rect 5868 3448 5874 3460
rect 6656 3448 6684 3479
rect 5868 3420 6684 3448
rect 5868 3408 5874 3420
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 7484 3448 7512 3488
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10060 3516 10088 3556
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10226 3544 10232 3596
rect 10284 3544 10290 3596
rect 10404 3587 10462 3593
rect 10404 3553 10416 3587
rect 10450 3584 10462 3587
rect 11606 3584 11612 3596
rect 10450 3556 11612 3584
rect 10450 3553 10462 3556
rect 10404 3547 10462 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 10244 3516 10272 3544
rect 11716 3516 11744 3624
rect 12038 3621 12050 3624
rect 12124 3652 12130 3664
rect 12124 3624 12186 3652
rect 12038 3615 12072 3621
rect 12066 3612 12072 3615
rect 12124 3612 12130 3624
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 13096 3584 13124 3692
rect 13173 3689 13185 3723
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 16114 3720 16120 3732
rect 15703 3692 16120 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 13188 3652 13216 3683
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 22462 3720 22468 3732
rect 16816 3692 22468 3720
rect 16816 3680 16822 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 13446 3652 13452 3664
rect 13188 3624 13452 3652
rect 13446 3612 13452 3624
rect 13504 3652 13510 3664
rect 13694 3655 13752 3661
rect 13694 3652 13706 3655
rect 13504 3624 13706 3652
rect 13504 3612 13510 3624
rect 13694 3621 13706 3624
rect 13740 3621 13752 3655
rect 13694 3615 13752 3621
rect 13832 3624 20300 3652
rect 13832 3584 13860 3624
rect 15746 3584 15752 3596
rect 11839 3556 13032 3584
rect 13096 3556 13860 3584
rect 15707 3556 15752 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 9732 3488 9777 3516
rect 10060 3488 10272 3516
rect 11532 3488 11744 3516
rect 13004 3516 13032 3556
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 16298 3584 16304 3596
rect 16259 3556 16304 3584
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 17954 3584 17960 3596
rect 17915 3556 17960 3584
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 20272 3593 20300 3624
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3553 20315 3587
rect 20257 3547 20315 3553
rect 13446 3516 13452 3528
rect 13004 3488 13452 3516
rect 9732 3476 9738 3488
rect 11532 3457 11560 3488
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 15841 3479 15899 3485
rect 11517 3451 11575 3457
rect 6880 3420 7512 3448
rect 8772 3420 9260 3448
rect 6880 3408 6886 3420
rect 658 3340 664 3392
rect 716 3380 722 3392
rect 2774 3380 2780 3392
rect 716 3352 2780 3380
rect 716 3340 722 3352
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 5994 3380 6000 3392
rect 4212 3352 6000 3380
rect 4212 3340 4218 3352
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6089 3383 6147 3389
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 8772 3380 8800 3420
rect 6135 3352 8800 3380
rect 8849 3383 8907 3389
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 8849 3349 8861 3383
rect 8895 3380 8907 3383
rect 8938 3380 8944 3392
rect 8895 3352 8944 3380
rect 8895 3349 8907 3352
rect 8849 3343 8907 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9232 3380 9260 3420
rect 11517 3417 11529 3451
rect 11563 3417 11575 3451
rect 11517 3411 11575 3417
rect 14829 3451 14887 3457
rect 14829 3417 14841 3451
rect 14875 3448 14887 3451
rect 15010 3448 15016 3460
rect 14875 3420 15016 3448
rect 14875 3417 14887 3420
rect 14829 3411 14887 3417
rect 15010 3408 15016 3420
rect 15068 3448 15074 3460
rect 15856 3448 15884 3479
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 15068 3420 15884 3448
rect 15068 3408 15074 3420
rect 13446 3380 13452 3392
rect 9232 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 15289 3383 15347 3389
rect 15289 3349 15301 3383
rect 15335 3380 15347 3383
rect 15378 3380 15384 3392
rect 15335 3352 15384 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3380 18199 3383
rect 18782 3380 18788 3392
rect 18187 3352 18788 3380
rect 18187 3349 18199 3352
rect 18141 3343 18199 3349
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 20441 3383 20499 3389
rect 20441 3349 20453 3383
rect 20487 3380 20499 3383
rect 22002 3380 22008 3392
rect 20487 3352 22008 3380
rect 20487 3349 20499 3352
rect 20441 3343 20499 3349
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 3694 3176 3700 3188
rect 2056 3148 3700 3176
rect 2056 3049 2084 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5169 3179 5227 3185
rect 5169 3176 5181 3179
rect 4764 3148 5181 3176
rect 4764 3136 4770 3148
rect 5169 3145 5181 3148
rect 5215 3145 5227 3179
rect 5442 3176 5448 3188
rect 5403 3148 5448 3176
rect 5169 3139 5227 3145
rect 3418 3108 3424 3120
rect 3379 3080 3424 3108
rect 3418 3068 3424 3080
rect 3476 3068 3482 3120
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3752 3012 3801 3040
rect 3752 3000 3758 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 5184 3040 5212 3139
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6822 3176 6828 3188
rect 6052 3148 6828 3176
rect 6052 3136 6058 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 9033 3179 9091 3185
rect 7248 3148 8432 3176
rect 7248 3136 7254 3148
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6086 3108 6092 3120
rect 5592 3080 6092 3108
rect 5592 3068 5598 3080
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5184 3012 6009 3040
rect 3789 3003 3847 3009
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 5997 3003 6055 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 8404 3040 8432 3148
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9306 3176 9312 3188
rect 9079 3148 9312 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 11057 3179 11115 3185
rect 9600 3148 10824 3176
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 9600 3108 9628 3148
rect 8904 3080 9628 3108
rect 8904 3068 8910 3080
rect 9600 3049 9628 3080
rect 10045 3111 10103 3117
rect 10045 3077 10057 3111
rect 10091 3108 10103 3111
rect 10091 3080 10732 3108
rect 10091 3077 10103 3080
rect 10045 3071 10103 3077
rect 9585 3043 9643 3049
rect 8404 3012 9168 3040
rect 2774 2972 2780 2984
rect 2148 2944 2780 2972
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 2148 2904 2176 2944
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 7644 2975 7702 2981
rect 3988 2944 7420 2972
rect 1176 2876 2176 2904
rect 2308 2907 2366 2913
rect 1176 2864 1182 2876
rect 2308 2873 2320 2907
rect 2354 2904 2366 2907
rect 3988 2904 4016 2944
rect 2354 2876 4016 2904
rect 4056 2907 4114 2913
rect 2354 2873 2366 2876
rect 2308 2867 2366 2873
rect 4056 2873 4068 2907
rect 4102 2904 4114 2907
rect 5534 2904 5540 2916
rect 4102 2876 5540 2904
rect 4102 2873 4114 2876
rect 4056 2867 4114 2873
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2904 5871 2907
rect 6914 2904 6920 2916
rect 5859 2876 6920 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 5626 2836 5632 2848
rect 1636 2808 5632 2836
rect 1636 2796 1642 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 7392 2836 7420 2944
rect 7644 2941 7656 2975
rect 7690 2972 7702 2975
rect 8938 2972 8944 2984
rect 7690 2944 8944 2972
rect 7690 2941 7702 2944
rect 7644 2935 7702 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9140 2972 9168 3012
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 9824 3012 10517 3040
rect 9824 3000 9830 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9140 2944 9505 2972
rect 9493 2941 9505 2944
rect 9539 2972 9551 2975
rect 9858 2972 9864 2984
rect 9539 2944 9864 2972
rect 9539 2941 9551 2944
rect 9493 2935 9551 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 10612 2904 10640 3003
rect 8772 2876 10640 2904
rect 10704 2904 10732 3080
rect 10796 2972 10824 3148
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 16298 3176 16304 3188
rect 11103 3148 16304 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3108 12495 3111
rect 12483 3080 16160 3108
rect 12483 3077 12495 3080
rect 12437 3071 12495 3077
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11112 3012 11621 3040
rect 11112 3000 11118 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 12066 3000 12072 3052
rect 12124 3040 12130 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12124 3012 13001 3040
rect 12124 3000 12130 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 15930 3040 15936 3052
rect 12989 3003 13047 3009
rect 13096 3012 15936 3040
rect 13096 2972 13124 3012
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 13446 2972 13452 2984
rect 10796 2944 13124 2972
rect 13407 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14608 2944 14749 2972
rect 14608 2932 14614 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 14737 2935 14795 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 16132 2981 16160 3080
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 16393 2975 16451 2981
rect 16393 2941 16405 2975
rect 16439 2972 16451 2975
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16439 2944 17049 2972
rect 16439 2941 16451 2944
rect 16393 2935 16451 2941
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18748 2944 18797 2972
rect 18748 2932 18754 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 11790 2904 11796 2916
rect 10704 2876 11796 2904
rect 8772 2845 8800 2876
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 11940 2876 12817 2904
rect 11940 2864 11946 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13906 2904 13912 2916
rect 13771 2876 13912 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 17126 2904 17132 2916
rect 15703 2876 17132 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 17126 2864 17132 2876
rect 17184 2864 17190 2916
rect 20346 2904 20352 2916
rect 20307 2876 20352 2904
rect 20346 2864 20352 2876
rect 20404 2904 20410 2916
rect 20548 2904 20576 2935
rect 20404 2876 20576 2904
rect 20404 2864 20410 2876
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 5960 2808 6005 2836
rect 7392 2808 8769 2836
rect 5960 2796 5966 2808
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8757 2799 8815 2805
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 9180 2808 9413 2836
rect 9180 2796 9186 2808
rect 9401 2805 9413 2808
rect 9447 2805 9459 2839
rect 9401 2799 9459 2805
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 9640 2808 10425 2836
rect 9640 2796 9646 2808
rect 10413 2805 10425 2808
rect 10459 2805 10471 2839
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 10413 2799 10471 2805
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 12894 2836 12900 2848
rect 11572 2808 11617 2836
rect 12855 2808 12900 2836
rect 11572 2796 11578 2808
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13630 2796 13636 2848
rect 13688 2836 13694 2848
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 13688 2808 14381 2836
rect 13688 2796 13694 2808
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 14369 2799 14427 2805
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 14608 2808 14933 2836
rect 14608 2796 14614 2808
rect 14921 2805 14933 2808
rect 14967 2805 14979 2839
rect 14921 2799 14979 2805
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17862 2836 17868 2848
rect 17267 2808 17868 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18969 2839 19027 2845
rect 18969 2805 18981 2839
rect 19015 2836 19027 2839
rect 19702 2836 19708 2848
rect 19015 2808 19708 2836
rect 19015 2805 19027 2808
rect 18969 2799 19027 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 21542 2836 21548 2848
rect 20763 2808 21548 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2188 2604 2421 2632
rect 2188 2592 2194 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 2409 2595 2467 2601
rect 2792 2604 4077 2632
rect 2038 2524 2044 2576
rect 2096 2564 2102 2576
rect 2792 2564 2820 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4212 2604 4537 2632
rect 4212 2592 4218 2604
rect 4525 2601 4537 2604
rect 4571 2632 4583 2635
rect 4571 2604 4936 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 2096 2536 2820 2564
rect 2096 2524 2102 2536
rect 3418 2524 3424 2576
rect 3476 2564 3482 2576
rect 4614 2564 4620 2576
rect 3476 2536 4620 2564
rect 3476 2524 3482 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3142 2496 3148 2508
rect 2823 2468 3148 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3142 2456 3148 2468
rect 3200 2496 3206 2508
rect 3786 2496 3792 2508
rect 3200 2468 3792 2496
rect 3200 2456 3206 2468
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4212 2468 4445 2496
rect 4212 2456 4218 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4908 2496 4936 2604
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 5040 2604 5089 2632
rect 5040 2592 5046 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 5810 2632 5816 2644
rect 5675 2604 5816 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 5994 2632 6000 2644
rect 5955 2604 6000 2632
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7466 2632 7472 2644
rect 7423 2604 7472 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 9214 2632 9220 2644
rect 8067 2604 9220 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2601 9827 2635
rect 10134 2632 10140 2644
rect 10095 2604 10140 2632
rect 9769 2595 9827 2601
rect 6089 2567 6147 2573
rect 6089 2533 6101 2567
rect 6135 2564 6147 2567
rect 7190 2564 7196 2576
rect 6135 2536 7196 2564
rect 6135 2533 6147 2536
rect 6089 2527 6147 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 7484 2564 7512 2592
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 7484 2536 8493 2564
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 9784 2564 9812 2595
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10275 2604 10609 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 12894 2632 12900 2644
rect 10827 2604 12900 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 10689 2567 10747 2573
rect 10689 2564 10701 2567
rect 9784 2536 10701 2564
rect 8481 2527 8539 2533
rect 10689 2533 10701 2536
rect 10735 2533 10747 2567
rect 10689 2527 10747 2533
rect 10962 2524 10968 2576
rect 11020 2564 11026 2576
rect 11149 2567 11207 2573
rect 11149 2564 11161 2567
rect 11020 2536 11161 2564
rect 11020 2524 11026 2536
rect 11149 2533 11161 2536
rect 11195 2533 11207 2567
rect 11149 2527 11207 2533
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12115 2536 13400 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 6730 2496 6736 2508
rect 4908 2468 6736 2496
rect 4433 2459 4491 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7064 2468 7297 2496
rect 7064 2456 7070 2468
rect 7285 2465 7297 2468
rect 7331 2496 7343 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7331 2468 8401 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8389 2465 8401 2468
rect 8435 2496 8447 2499
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 8435 2468 11253 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 11241 2465 11253 2468
rect 11287 2465 11299 2499
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 11241 2459 11299 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 13372 2505 13400 2536
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12032 2468 12633 2496
rect 12032 2456 12038 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2465 13415 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13357 2459 13415 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14458 2496 14464 2508
rect 14419 2468 14464 2496
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16022 2496 16028 2508
rect 15983 2468 16028 2496
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16574 2496 16580 2508
rect 16535 2468 16580 2496
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 198 2388 204 2440
rect 256 2428 262 2440
rect 2866 2428 2872 2440
rect 256 2400 2872 2428
rect 256 2388 262 2400
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3418 2428 3424 2440
rect 3099 2400 3424 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 6144 2400 6285 2428
rect 6144 2388 6150 2400
rect 6273 2397 6285 2400
rect 6319 2428 6331 2431
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6319 2400 7481 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 8846 2428 8852 2440
rect 8711 2400 8852 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 11606 2428 11612 2440
rect 11471 2400 11612 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 14182 2428 14188 2440
rect 12943 2400 14188 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 10962 2360 10968 2372
rect 2832 2332 10968 2360
rect 2832 2320 2838 2332
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 11514 2320 11520 2372
rect 11572 2320 11578 2372
rect 16761 2363 16819 2369
rect 16761 2329 16773 2363
rect 16807 2360 16819 2363
rect 17402 2360 17408 2372
rect 16807 2332 17408 2360
rect 16807 2329 16819 2332
rect 16761 2323 16819 2329
rect 17402 2320 17408 2332
rect 17460 2320 17466 2372
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 4154 2292 4160 2304
rect 3016 2264 4160 2292
rect 3016 2252 3022 2264
rect 4154 2252 4160 2264
rect 4212 2292 4218 2304
rect 5074 2292 5080 2304
rect 4212 2264 5080 2292
rect 4212 2252 4218 2264
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 7466 2292 7472 2304
rect 5684 2264 7472 2292
rect 5684 2252 5690 2264
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 7708 2264 10609 2292
rect 7708 2252 7714 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 10689 2295 10747 2301
rect 10689 2261 10701 2295
rect 10735 2292 10747 2295
rect 11532 2292 11560 2320
rect 10735 2264 11560 2292
rect 10735 2261 10747 2264
rect 10689 2255 10747 2261
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13228 2264 13553 2292
rect 13228 2252 13234 2264
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 14090 2292 14096 2304
rect 14051 2264 14096 2292
rect 13541 2255 13599 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14645 2295 14703 2301
rect 14645 2261 14657 2295
rect 14691 2292 14703 2295
rect 15010 2292 15016 2304
rect 14691 2264 15016 2292
rect 14691 2261 14703 2264
rect 14645 2255 14703 2261
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15620 2264 15669 2292
rect 15620 2252 15626 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16209 2295 16267 2301
rect 16209 2292 16221 2295
rect 16080 2264 16221 2292
rect 16080 2252 16086 2264
rect 16209 2261 16221 2264
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 17313 2295 17371 2301
rect 17313 2261 17325 2295
rect 17359 2292 17371 2295
rect 17954 2292 17960 2304
rect 17359 2264 17960 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 4062 2088 4068 2100
rect 2096 2060 4068 2088
rect 2096 2048 2102 2060
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 7282 1368 7288 1420
rect 7340 1408 7346 1420
rect 8110 1408 8116 1420
rect 7340 1380 8116 1408
rect 7340 1368 7346 1380
rect 8110 1368 8116 1380
rect 8168 1368 8174 1420
rect 3326 484 3332 536
rect 3384 524 3390 536
rect 4890 524 4896 536
rect 3384 496 4896 524
rect 3384 484 3390 496
rect 4890 484 4896 496
rect 4948 484 4954 536
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2780 20000 2832 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 4804 19864 4856 19916
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3056 19499 3108 19508
rect 3056 19465 3065 19499
rect 3065 19465 3099 19499
rect 3099 19465 3108 19499
rect 3056 19456 3108 19465
rect 2136 19252 2188 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 10600 19252 10652 19304
rect 2872 19116 2924 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1860 18955 1912 18964
rect 1860 18921 1869 18955
rect 1869 18921 1903 18955
rect 1903 18921 1912 18955
rect 1860 18912 1912 18921
rect 7196 18912 7248 18964
rect 2320 18844 2372 18896
rect 8392 18776 8444 18828
rect 1768 18708 1820 18760
rect 3332 18640 3384 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 3240 18411 3292 18420
rect 3240 18377 3249 18411
rect 3249 18377 3283 18411
rect 3283 18377 3292 18411
rect 3240 18368 3292 18377
rect 2136 18232 2188 18284
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 1860 18164 1912 18216
rect 8300 18164 8352 18216
rect 11060 18164 11112 18216
rect 8668 18096 8720 18148
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 1860 17756 1912 17808
rect 3332 17799 3384 17808
rect 3332 17765 3341 17799
rect 3341 17765 3375 17799
rect 3375 17765 3384 17799
rect 3332 17756 3384 17765
rect 4804 17756 4856 17808
rect 8300 17756 8352 17808
rect 11612 17756 11664 17808
rect 2872 17620 2924 17672
rect 6276 17620 6328 17672
rect 7748 17688 7800 17740
rect 10324 17688 10376 17740
rect 9036 17620 9088 17672
rect 13636 17620 13688 17672
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 5724 17212 5776 17264
rect 5080 17187 5132 17196
rect 2872 17076 2924 17128
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 11152 17144 11204 17196
rect 9772 17076 9824 17128
rect 6736 17008 6788 17060
rect 9128 17008 9180 17060
rect 3792 16940 3844 16992
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 10048 16983 10100 16992
rect 4896 16940 4948 16949
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 1492 16668 1544 16720
rect 5080 16736 5132 16788
rect 5356 16736 5408 16788
rect 7748 16779 7800 16788
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 10692 16736 10744 16788
rect 13636 16779 13688 16788
rect 3792 16668 3844 16720
rect 4712 16668 4764 16720
rect 9588 16668 9640 16720
rect 13636 16745 13645 16779
rect 13645 16745 13679 16779
rect 13679 16745 13688 16779
rect 13636 16736 13688 16745
rect 17868 16736 17920 16788
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 6644 16600 6696 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 9772 16600 9824 16652
rect 11152 16600 11204 16652
rect 12072 16668 12124 16720
rect 3332 16532 3384 16584
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 9128 16532 9180 16584
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 6000 16192 6052 16244
rect 7012 16192 7064 16244
rect 9128 16235 9180 16244
rect 9128 16201 9137 16235
rect 9137 16201 9171 16235
rect 9171 16201 9180 16235
rect 9128 16192 9180 16201
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 1676 16056 1728 16108
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 9772 16099 9824 16108
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 2872 15988 2924 16040
rect 5356 16031 5408 16040
rect 5356 15997 5390 16031
rect 5390 15997 5408 16031
rect 3976 15920 4028 15972
rect 5356 15988 5408 15997
rect 7472 15988 7524 16040
rect 5632 15920 5684 15972
rect 8852 15920 8904 15972
rect 10048 15963 10100 15972
rect 10048 15929 10082 15963
rect 10082 15929 10100 15963
rect 10048 15920 10100 15929
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 4712 15895 4764 15904
rect 4712 15861 4721 15895
rect 4721 15861 4755 15895
rect 4755 15861 4764 15895
rect 4712 15852 4764 15861
rect 5264 15852 5316 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 2044 15648 2096 15700
rect 4896 15648 4948 15700
rect 5172 15648 5224 15700
rect 8852 15691 8904 15700
rect 6000 15623 6052 15632
rect 6000 15589 6034 15623
rect 6034 15589 6052 15623
rect 6000 15580 6052 15589
rect 2044 15512 2096 15564
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 3976 15444 4028 15496
rect 6368 15512 6420 15564
rect 7748 15555 7800 15564
rect 7748 15521 7782 15555
rect 7782 15521 7800 15555
rect 7748 15512 7800 15521
rect 8852 15657 8861 15691
rect 8861 15657 8895 15691
rect 8895 15657 8904 15691
rect 8852 15648 8904 15657
rect 9588 15648 9640 15700
rect 11152 15648 11204 15700
rect 11612 15648 11664 15700
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 5632 15444 5684 15496
rect 7472 15487 7524 15496
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 2780 15308 2832 15360
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 7104 15351 7156 15360
rect 7104 15317 7113 15351
rect 7113 15317 7147 15351
rect 7147 15317 7156 15351
rect 7104 15308 7156 15317
rect 7656 15308 7708 15360
rect 12256 15512 12308 15564
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 11152 15308 11204 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2872 15104 2924 15156
rect 3976 15147 4028 15156
rect 3976 15113 3985 15147
rect 3985 15113 4019 15147
rect 4019 15113 4028 15147
rect 3976 15104 4028 15113
rect 4160 15104 4212 15156
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 7196 15104 7248 15156
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 7104 14968 7156 15020
rect 7748 14968 7800 15020
rect 10784 15104 10836 15156
rect 10048 14968 10100 15020
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 2688 14900 2740 14952
rect 6460 14900 6512 14952
rect 6644 14900 6696 14952
rect 3700 14832 3752 14884
rect 6828 14832 6880 14884
rect 8208 14900 8260 14952
rect 9772 14900 9824 14952
rect 8576 14764 8628 14816
rect 9312 14832 9364 14884
rect 11612 14764 11664 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 3332 14560 3384 14612
rect 7472 14560 7524 14612
rect 8208 14560 8260 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 9772 14560 9824 14612
rect 3056 14492 3108 14544
rect 3608 14424 3660 14476
rect 1492 14356 1544 14408
rect 3700 14331 3752 14340
rect 3700 14297 3709 14331
rect 3709 14297 3743 14331
rect 3743 14297 3752 14331
rect 3700 14288 3752 14297
rect 2596 14220 2648 14272
rect 4252 14220 4304 14272
rect 5632 14424 5684 14476
rect 6184 14424 6236 14476
rect 7104 14492 7156 14544
rect 8300 14492 8352 14544
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 8852 14356 8904 14408
rect 7748 14288 7800 14340
rect 9312 14356 9364 14408
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 10876 14288 10928 14340
rect 7104 14220 7156 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1860 14016 1912 14068
rect 3240 13948 3292 14000
rect 2320 13880 2372 13932
rect 2688 13880 2740 13932
rect 3608 13880 3660 13932
rect 9312 14016 9364 14068
rect 6184 13880 6236 13932
rect 6552 13880 6604 13932
rect 3792 13744 3844 13796
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 5724 13812 5776 13864
rect 9772 13812 9824 13864
rect 5448 13744 5500 13796
rect 7748 13744 7800 13796
rect 9220 13744 9272 13796
rect 5080 13676 5132 13728
rect 7196 13676 7248 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 9680 13472 9732 13524
rect 2044 13447 2096 13456
rect 2044 13413 2053 13447
rect 2053 13413 2087 13447
rect 2087 13413 2096 13447
rect 2044 13404 2096 13413
rect 2228 13404 2280 13456
rect 8576 13404 8628 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 1676 13200 1728 13252
rect 4160 13336 4212 13388
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 6460 13336 6512 13388
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 5448 13268 5500 13320
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 9220 13311 9272 13320
rect 8392 13200 8444 13252
rect 5172 13132 5224 13184
rect 7288 13132 7340 13184
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9772 13336 9824 13388
rect 9956 13379 10008 13388
rect 9956 13345 9990 13379
rect 9990 13345 10008 13379
rect 9956 13336 10008 13345
rect 9220 13268 9272 13277
rect 9680 13132 9732 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 1768 12928 1820 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3148 12792 3200 12844
rect 4160 12928 4212 12980
rect 6736 12928 6788 12980
rect 8392 12928 8444 12980
rect 8668 12928 8720 12980
rect 9956 12928 10008 12980
rect 3792 12860 3844 12912
rect 4988 12792 5040 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 8208 12792 8260 12844
rect 2688 12724 2740 12776
rect 4620 12724 4672 12776
rect 5172 12724 5224 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 9312 12724 9364 12776
rect 9772 12724 9824 12776
rect 4344 12656 4396 12708
rect 6184 12656 6236 12708
rect 8208 12656 8260 12708
rect 8852 12656 8904 12708
rect 9220 12656 9272 12708
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 2320 12588 2372 12597
rect 2964 12588 3016 12640
rect 4160 12588 4212 12640
rect 5540 12588 5592 12640
rect 6460 12588 6512 12640
rect 6644 12588 6696 12640
rect 8484 12588 8536 12640
rect 10784 12588 10836 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1768 12384 1820 12436
rect 2320 12384 2372 12436
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 2780 12316 2832 12368
rect 4068 12316 4120 12368
rect 6552 12316 6604 12368
rect 2320 12248 2372 12300
rect 3332 12248 3384 12300
rect 5080 12291 5132 12300
rect 5080 12257 5114 12291
rect 5114 12257 5132 12291
rect 5080 12248 5132 12257
rect 6460 12248 6512 12300
rect 8392 12384 8444 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 7472 12316 7524 12368
rect 9956 12316 10008 12368
rect 4712 12112 4764 12164
rect 6092 12180 6144 12232
rect 6552 12180 6604 12232
rect 8300 12180 8352 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 4804 12044 4856 12096
rect 6736 12112 6788 12164
rect 6092 12044 6144 12096
rect 6552 12044 6604 12096
rect 10324 12112 10376 12164
rect 8944 12044 8996 12096
rect 11704 12044 11756 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 5080 11840 5132 11892
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 9220 11840 9272 11892
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 4252 11704 4304 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 2872 11636 2924 11688
rect 7104 11704 7156 11756
rect 8852 11704 8904 11756
rect 3148 11568 3200 11620
rect 1860 11500 1912 11552
rect 2780 11500 2832 11552
rect 4252 11500 4304 11552
rect 4344 11500 4396 11552
rect 4528 11500 4580 11552
rect 4804 11636 4856 11688
rect 4712 11568 4764 11620
rect 5264 11636 5316 11688
rect 6000 11636 6052 11688
rect 8484 11636 8536 11688
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 5632 11568 5684 11620
rect 5816 11568 5868 11620
rect 8668 11611 8720 11620
rect 8668 11577 8677 11611
rect 8677 11577 8711 11611
rect 8711 11577 8720 11611
rect 8668 11568 8720 11577
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 11060 11568 11112 11620
rect 9772 11500 9824 11552
rect 20904 11500 20956 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 4160 11296 4212 11348
rect 4712 11296 4764 11348
rect 4896 11296 4948 11348
rect 8760 11296 8812 11348
rect 9956 11296 10008 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 11704 11296 11756 11348
rect 20260 11296 20312 11348
rect 5724 11228 5776 11280
rect 8944 11228 8996 11280
rect 9588 11228 9640 11280
rect 3148 11092 3200 11144
rect 3240 11092 3292 11144
rect 3608 11024 3660 11076
rect 4712 11160 4764 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6184 11160 6236 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 8760 11203 8812 11212
rect 8760 11169 8769 11203
rect 8769 11169 8803 11203
rect 8803 11169 8812 11203
rect 8760 11160 8812 11169
rect 10416 11160 10468 11212
rect 12440 11160 12492 11212
rect 4804 11092 4856 11144
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 8852 11135 8904 11144
rect 8852 11101 8861 11135
rect 8861 11101 8895 11135
rect 8895 11101 8904 11135
rect 8852 11092 8904 11101
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 12348 11092 12400 11144
rect 5172 11024 5224 11076
rect 3976 10956 4028 11008
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 20628 11024 20680 11076
rect 11060 10956 11112 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2964 10752 3016 10804
rect 5632 10752 5684 10804
rect 9772 10752 9824 10804
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 2872 10616 2924 10668
rect 7380 10616 7432 10668
rect 2780 10548 2832 10600
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 4896 10548 4948 10600
rect 5080 10548 5132 10600
rect 7564 10548 7616 10600
rect 8116 10548 8168 10600
rect 3148 10480 3200 10532
rect 4804 10480 4856 10532
rect 5448 10480 5500 10532
rect 2872 10412 2924 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 4068 10412 4120 10464
rect 6092 10412 6144 10464
rect 9312 10480 9364 10532
rect 9680 10548 9732 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11060 10548 11112 10600
rect 12532 10480 12584 10532
rect 10416 10412 10468 10464
rect 20168 10412 20220 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2504 10208 2556 10260
rect 4068 10208 4120 10260
rect 4436 10208 4488 10260
rect 5080 10208 5132 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 6276 10208 6328 10260
rect 7012 10208 7064 10260
rect 8392 10208 8444 10260
rect 9036 10208 9088 10260
rect 10968 10208 11020 10260
rect 3332 10183 3384 10192
rect 3332 10149 3341 10183
rect 3341 10149 3375 10183
rect 3375 10149 3384 10183
rect 3332 10140 3384 10149
rect 4252 10140 4304 10192
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 2964 10072 3016 10124
rect 4160 10072 4212 10124
rect 2688 10047 2740 10056
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 10600 10072 10652 10124
rect 6828 10004 6880 10056
rect 7104 10004 7156 10056
rect 7564 10004 7616 10056
rect 9036 10047 9088 10056
rect 9036 10013 9045 10047
rect 9045 10013 9079 10047
rect 9079 10013 9088 10047
rect 9036 10004 9088 10013
rect 10416 10004 10468 10056
rect 7012 9936 7064 9988
rect 3516 9868 3568 9920
rect 10048 9868 10100 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3700 9664 3752 9716
rect 9036 9664 9088 9716
rect 3148 9639 3200 9648
rect 3148 9605 3157 9639
rect 3157 9605 3191 9639
rect 3191 9605 3200 9639
rect 3148 9596 3200 9605
rect 4712 9596 4764 9648
rect 4896 9596 4948 9648
rect 5264 9596 5316 9648
rect 5540 9639 5592 9648
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 4252 9528 4304 9580
rect 5632 9528 5684 9580
rect 6276 9528 6328 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 3792 9460 3844 9512
rect 2688 9392 2740 9444
rect 2228 9324 2280 9376
rect 5724 9392 5776 9444
rect 4804 9324 4856 9376
rect 5172 9324 5224 9376
rect 5448 9324 5500 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 9404 9324 9456 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2412 9120 2464 9172
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 4160 9120 4212 9172
rect 7196 9120 7248 9172
rect 7564 9120 7616 9172
rect 8668 9120 8720 9172
rect 4068 9052 4120 9104
rect 5080 9052 5132 9104
rect 5264 9052 5316 9104
rect 3332 9027 3384 9036
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 3332 8984 3384 8993
rect 5356 8984 5408 9036
rect 6276 8984 6328 9036
rect 8208 9052 8260 9104
rect 1952 8916 2004 8968
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3700 8916 3752 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 6276 8848 6328 8900
rect 5264 8780 5316 8832
rect 9772 8984 9824 9036
rect 10324 8984 10376 9036
rect 8484 8780 8536 8832
rect 10692 8848 10744 8900
rect 12716 8848 12768 8900
rect 10784 8780 10836 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2688 8576 2740 8628
rect 3700 8576 3752 8628
rect 5356 8576 5408 8628
rect 7196 8576 7248 8628
rect 7380 8576 7432 8628
rect 7656 8576 7708 8628
rect 4252 8508 4304 8560
rect 7104 8508 7156 8560
rect 6276 8483 6328 8492
rect 6276 8449 6285 8483
rect 6285 8449 6319 8483
rect 6319 8449 6328 8483
rect 6276 8440 6328 8449
rect 10692 8576 10744 8628
rect 10784 8576 10836 8628
rect 8484 8483 8536 8492
rect 2228 8304 2280 8356
rect 4712 8372 4764 8424
rect 7380 8372 7432 8424
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 3608 8304 3660 8356
rect 3792 8304 3844 8356
rect 8760 8304 8812 8356
rect 11060 8304 11112 8356
rect 4712 8236 4764 8288
rect 5080 8236 5132 8288
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 7012 8236 7064 8288
rect 9496 8279 9548 8288
rect 9496 8245 9505 8279
rect 9505 8245 9539 8279
rect 9539 8245 9548 8279
rect 9496 8236 9548 8245
rect 11428 8279 11480 8288
rect 11428 8245 11437 8279
rect 11437 8245 11471 8279
rect 11471 8245 11480 8279
rect 11428 8236 11480 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 2136 8032 2188 8084
rect 3332 8032 3384 8084
rect 4068 8075 4120 8084
rect 4068 8041 4077 8075
rect 4077 8041 4111 8075
rect 4111 8041 4120 8075
rect 4068 8032 4120 8041
rect 5816 8032 5868 8084
rect 6092 8032 6144 8084
rect 6920 8032 6972 8084
rect 7288 8032 7340 8084
rect 7380 8032 7432 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 11428 8032 11480 8084
rect 5264 8007 5316 8016
rect 1952 7896 2004 7948
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 1860 7828 1912 7880
rect 2780 7828 2832 7880
rect 5264 7973 5298 8007
rect 5298 7973 5316 8007
rect 5264 7964 5316 7973
rect 7196 7964 7248 8016
rect 4712 7896 4764 7948
rect 6920 7896 6972 7948
rect 9496 7964 9548 8016
rect 10232 7896 10284 7948
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 6828 7828 6880 7880
rect 8484 7828 8536 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 12348 7896 12400 7948
rect 13820 7896 13872 7948
rect 4252 7692 4304 7744
rect 4712 7692 4764 7744
rect 11060 7760 11112 7812
rect 9956 7692 10008 7744
rect 18696 7828 18748 7880
rect 11980 7692 12032 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 3424 7488 3476 7540
rect 3884 7488 3936 7540
rect 7748 7488 7800 7540
rect 13820 7531 13872 7540
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 3608 7352 3660 7404
rect 7656 7352 7708 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 3792 7284 3844 7336
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 7472 7284 7524 7336
rect 8392 7284 8444 7336
rect 10692 7284 10744 7336
rect 12348 7284 12400 7336
rect 13820 7497 13829 7531
rect 13829 7497 13863 7531
rect 13863 7497 13872 7531
rect 13820 7488 13872 7497
rect 16488 7420 16540 7472
rect 13820 7352 13872 7404
rect 16580 7284 16632 7336
rect 5908 7216 5960 7268
rect 1492 7148 1544 7200
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 2780 7148 2832 7200
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 9956 7216 10008 7268
rect 12624 7216 12676 7268
rect 12808 7216 12860 7268
rect 12992 7216 13044 7268
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8760 7191 8812 7200
rect 8760 7157 8769 7191
rect 8769 7157 8803 7191
rect 8803 7157 8812 7191
rect 8760 7148 8812 7157
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 11060 7148 11112 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 3976 6944 4028 6996
rect 5632 6944 5684 6996
rect 1768 6876 1820 6928
rect 5540 6876 5592 6928
rect 6460 6876 6512 6928
rect 8760 6944 8812 6996
rect 7656 6919 7708 6928
rect 7656 6885 7690 6919
rect 7690 6885 7708 6919
rect 7656 6876 7708 6885
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 2504 6851 2556 6860
rect 2504 6817 2538 6851
rect 2538 6817 2556 6851
rect 2504 6808 2556 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 4896 6808 4948 6860
rect 5080 6808 5132 6860
rect 8208 6808 8260 6860
rect 10508 6944 10560 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 10968 6876 11020 6928
rect 12808 6876 12860 6928
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 9772 6740 9824 6792
rect 9956 6740 10008 6792
rect 11796 6740 11848 6792
rect 13820 6808 13872 6860
rect 16120 6808 16172 6860
rect 16488 6808 16540 6860
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 14372 6740 14424 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 1492 6604 1544 6656
rect 3332 6672 3384 6724
rect 8944 6672 8996 6724
rect 12992 6672 13044 6724
rect 3240 6604 3292 6656
rect 4896 6604 4948 6656
rect 5908 6604 5960 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2504 6400 2556 6452
rect 4896 6400 4948 6452
rect 12440 6400 12492 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 6920 6332 6972 6384
rect 9956 6332 10008 6384
rect 11244 6332 11296 6384
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 7012 6264 7064 6316
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2228 6196 2280 6248
rect 3976 6196 4028 6248
rect 8944 6196 8996 6248
rect 9128 6196 9180 6248
rect 10508 6196 10560 6248
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 2504 6060 2556 6112
rect 2872 6060 2924 6112
rect 4712 6128 4764 6180
rect 5632 6171 5684 6180
rect 5632 6137 5641 6171
rect 5641 6137 5675 6171
rect 5675 6137 5684 6171
rect 5632 6128 5684 6137
rect 7748 6128 7800 6180
rect 7840 6128 7892 6180
rect 12348 6196 12400 6248
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 17684 6196 17736 6248
rect 12808 6128 12860 6180
rect 16028 6128 16080 6180
rect 16304 6128 16356 6180
rect 16856 6171 16908 6180
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 3792 6060 3844 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 5816 6060 5868 6112
rect 6092 6060 6144 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10140 6060 10192 6112
rect 10232 6060 10284 6112
rect 13176 6060 13228 6112
rect 13912 6060 13964 6112
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 19248 6060 19300 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 2320 5856 2372 5908
rect 2780 5856 2832 5908
rect 3332 5899 3384 5908
rect 3332 5865 3341 5899
rect 3341 5865 3375 5899
rect 3375 5865 3384 5899
rect 3332 5856 3384 5865
rect 5356 5856 5408 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 8484 5899 8536 5908
rect 3884 5788 3936 5840
rect 2964 5720 3016 5772
rect 5264 5788 5316 5840
rect 7196 5788 7248 5840
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 10140 5856 10192 5908
rect 11060 5856 11112 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 14464 5856 14516 5908
rect 7012 5720 7064 5772
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3792 5652 3844 5704
rect 4160 5652 4212 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 6460 5652 6512 5704
rect 11796 5788 11848 5840
rect 16580 5788 16632 5840
rect 11980 5720 12032 5772
rect 10784 5652 10836 5704
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11244 5652 11296 5704
rect 12440 5652 12492 5704
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 5632 5516 5684 5568
rect 6920 5516 6972 5568
rect 10140 5516 10192 5568
rect 15108 5584 15160 5636
rect 13176 5516 13228 5568
rect 14372 5516 14424 5568
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 16948 5516 17000 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 11796 5355 11848 5364
rect 6460 5244 6512 5296
rect 6828 5287 6880 5296
rect 6828 5253 6837 5287
rect 6837 5253 6871 5287
rect 6871 5253 6880 5287
rect 6828 5244 6880 5253
rect 6920 5244 6972 5296
rect 7196 5244 7248 5296
rect 2872 5176 2924 5228
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 4712 5176 4764 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 7012 5176 7064 5228
rect 7748 5176 7800 5228
rect 8392 5176 8444 5228
rect 9956 5176 10008 5228
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12624 5312 12676 5364
rect 13084 5312 13136 5364
rect 16120 5312 16172 5364
rect 11704 5244 11756 5296
rect 11980 5176 12032 5228
rect 16580 5219 16632 5228
rect 3332 5108 3384 5160
rect 3792 5108 3844 5160
rect 5816 5108 5868 5160
rect 6828 5108 6880 5160
rect 12532 5108 12584 5160
rect 13912 5151 13964 5160
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2320 4972 2372 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 8484 5040 8536 5092
rect 5080 4972 5132 4981
rect 6276 4972 6328 5024
rect 8208 4972 8260 5024
rect 12624 5040 12676 5092
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14372 5108 14424 5160
rect 16580 5185 16589 5219
rect 16589 5185 16623 5219
rect 16623 5185 16632 5219
rect 16580 5176 16632 5185
rect 16764 5108 16816 5160
rect 11704 4972 11756 5024
rect 11888 4972 11940 5024
rect 15844 5040 15896 5092
rect 15476 4972 15528 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 3148 4768 3200 4820
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 5080 4768 5132 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 9956 4768 10008 4820
rect 11888 4811 11940 4820
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 15292 4768 15344 4820
rect 3516 4700 3568 4752
rect 2872 4632 2924 4684
rect 3332 4632 3384 4684
rect 3884 4632 3936 4684
rect 1400 4564 1452 4616
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 3700 4564 3752 4616
rect 8300 4700 8352 4752
rect 4896 4632 4948 4684
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 6368 4632 6420 4684
rect 9128 4632 9180 4684
rect 14556 4700 14608 4752
rect 9772 4632 9824 4684
rect 10324 4632 10376 4684
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 16672 4675 16724 4684
rect 5540 4564 5592 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8944 4564 8996 4616
rect 11888 4564 11940 4616
rect 16672 4641 16681 4675
rect 16681 4641 16715 4675
rect 16715 4641 16724 4675
rect 16672 4632 16724 4641
rect 14464 4564 14516 4616
rect 16120 4564 16172 4616
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 15844 4496 15896 4548
rect 9588 4428 9640 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 17040 4428 17092 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2320 4224 2372 4276
rect 2872 4224 2924 4276
rect 6828 4267 6880 4276
rect 6828 4233 6837 4267
rect 6837 4233 6871 4267
rect 6871 4233 6880 4267
rect 6828 4224 6880 4233
rect 8208 4224 8260 4276
rect 8300 4224 8352 4276
rect 16672 4224 16724 4276
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 15844 4199 15896 4208
rect 6368 4156 6420 4165
rect 4068 4088 4120 4140
rect 4252 4088 4304 4140
rect 4436 4088 4488 4140
rect 4896 4088 4948 4140
rect 15844 4165 15853 4199
rect 15853 4165 15887 4199
rect 15887 4165 15896 4199
rect 15844 4156 15896 4165
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8852 4088 8904 4140
rect 8944 4088 8996 4140
rect 9956 4088 10008 4140
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 1676 4020 1728 4072
rect 5080 4020 5132 4072
rect 3148 3952 3200 4004
rect 5816 3952 5868 4004
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 5540 3884 5592 3936
rect 6736 4020 6788 4072
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 9772 3952 9824 4004
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9680 3884 9732 3936
rect 10140 3884 10192 3936
rect 10600 4020 10652 4072
rect 12164 4020 12216 4072
rect 11060 3952 11112 4004
rect 13544 4020 13596 4072
rect 14372 4020 14424 4072
rect 18052 4088 18104 4140
rect 17040 4063 17092 4072
rect 13176 3995 13228 4004
rect 13176 3961 13185 3995
rect 13185 3961 13219 3995
rect 13219 3961 13228 3995
rect 13176 3952 13228 3961
rect 13360 3952 13412 4004
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 17132 4020 17184 4072
rect 19892 4063 19944 4072
rect 19892 4029 19926 4063
rect 19926 4029 19944 4063
rect 19892 4020 19944 4029
rect 15016 3952 15068 4004
rect 15936 3952 15988 4004
rect 11612 3884 11664 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 15752 3884 15804 3936
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17960 3952 18012 4004
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 3516 3680 3568 3732
rect 3700 3680 3752 3732
rect 4068 3680 4120 3732
rect 1676 3612 1728 3664
rect 2780 3612 2832 3664
rect 4160 3612 4212 3664
rect 4712 3655 4764 3664
rect 4712 3621 4746 3655
rect 4746 3621 4764 3655
rect 4712 3612 4764 3621
rect 4896 3612 4948 3664
rect 5356 3612 5408 3664
rect 6460 3655 6512 3664
rect 6460 3621 6469 3655
rect 6469 3621 6503 3655
rect 6503 3621 6512 3655
rect 6460 3612 6512 3621
rect 6552 3612 6604 3664
rect 7564 3612 7616 3664
rect 9128 3655 9180 3664
rect 3424 3544 3476 3596
rect 2504 3476 2556 3528
rect 7012 3544 7064 3596
rect 7196 3544 7248 3596
rect 7380 3544 7432 3596
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 5448 3476 5500 3528
rect 8852 3544 8904 3596
rect 9128 3621 9137 3655
rect 9137 3621 9171 3655
rect 9171 3621 9180 3655
rect 9128 3612 9180 3621
rect 9956 3612 10008 3664
rect 12072 3655 12124 3664
rect 3700 3408 3752 3460
rect 5816 3451 5868 3460
rect 5816 3417 5825 3451
rect 5825 3417 5859 3451
rect 5859 3417 5868 3451
rect 5816 3408 5868 3417
rect 6828 3408 6880 3460
rect 9128 3476 9180 3528
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 10232 3544 10284 3596
rect 11612 3544 11664 3596
rect 12072 3621 12084 3655
rect 12084 3621 12124 3655
rect 12072 3612 12124 3621
rect 16120 3680 16172 3732
rect 16764 3680 16816 3732
rect 22468 3680 22520 3732
rect 13452 3612 13504 3664
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 13452 3519 13504 3528
rect 9680 3476 9732 3485
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 16580 3519 16632 3528
rect 664 3340 716 3392
rect 2780 3340 2832 3392
rect 4160 3340 4212 3392
rect 6000 3340 6052 3392
rect 8944 3340 8996 3392
rect 15016 3408 15068 3460
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 13452 3340 13504 3392
rect 15384 3340 15436 3392
rect 18788 3340 18840 3392
rect 22008 3340 22060 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 3700 3136 3752 3188
rect 4712 3136 4764 3188
rect 5448 3179 5500 3188
rect 3424 3111 3476 3120
rect 3424 3077 3433 3111
rect 3433 3077 3467 3111
rect 3467 3077 3476 3111
rect 3424 3068 3476 3077
rect 3700 3000 3752 3052
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 6000 3136 6052 3188
rect 6828 3136 6880 3188
rect 7196 3136 7248 3188
rect 5540 3068 5592 3120
rect 6092 3068 6144 3120
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 9312 3136 9364 3188
rect 8852 3068 8904 3120
rect 1124 2864 1176 2916
rect 2780 2932 2832 2984
rect 5540 2864 5592 2916
rect 6920 2864 6972 2916
rect 1584 2796 1636 2848
rect 5632 2796 5684 2848
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 8944 2932 8996 2984
rect 9772 3000 9824 3052
rect 9864 2932 9916 2984
rect 16304 3136 16356 3188
rect 11060 3000 11112 3052
rect 12072 3000 12124 3052
rect 15936 3000 15988 3052
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 14556 2932 14608 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 18696 2932 18748 2984
rect 11796 2864 11848 2916
rect 11888 2864 11940 2916
rect 13912 2864 13964 2916
rect 17132 2864 17184 2916
rect 20352 2907 20404 2916
rect 20352 2873 20361 2907
rect 20361 2873 20395 2907
rect 20395 2873 20404 2907
rect 20352 2864 20404 2873
rect 5908 2796 5960 2805
rect 9128 2796 9180 2848
rect 9588 2796 9640 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 12900 2839 12952 2848
rect 11520 2796 11572 2805
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 13636 2796 13688 2848
rect 14556 2796 14608 2848
rect 17868 2796 17920 2848
rect 19708 2796 19760 2848
rect 21548 2796 21600 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2136 2592 2188 2644
rect 2044 2524 2096 2576
rect 4160 2592 4212 2644
rect 3424 2524 3476 2576
rect 4620 2524 4672 2576
rect 3148 2456 3200 2508
rect 3792 2456 3844 2508
rect 4160 2456 4212 2508
rect 4988 2592 5040 2644
rect 5816 2592 5868 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7472 2592 7524 2644
rect 9220 2592 9272 2644
rect 10140 2635 10192 2644
rect 7196 2524 7248 2576
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 12900 2592 12952 2644
rect 10968 2524 11020 2576
rect 6736 2456 6788 2508
rect 7012 2456 7064 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 11980 2456 12032 2508
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 14464 2499 14516 2508
rect 14464 2465 14473 2499
rect 14473 2465 14507 2499
rect 14507 2465 14516 2499
rect 14464 2456 14516 2465
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 204 2388 256 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3424 2388 3476 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 6092 2388 6144 2440
rect 8852 2388 8904 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11612 2388 11664 2440
rect 14188 2388 14240 2440
rect 2780 2320 2832 2372
rect 10968 2320 11020 2372
rect 11520 2320 11572 2372
rect 17408 2320 17460 2372
rect 2964 2252 3016 2304
rect 4160 2252 4212 2304
rect 5080 2252 5132 2304
rect 5632 2252 5684 2304
rect 7472 2252 7524 2304
rect 7656 2252 7708 2304
rect 13176 2252 13228 2304
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 15016 2252 15068 2304
rect 15568 2252 15620 2304
rect 16028 2252 16080 2304
rect 17960 2252 18012 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2044 2048 2096 2100
rect 4068 2048 4120 2100
rect 7288 1368 7340 1420
rect 8116 1368 8168 1420
rect 3332 484 3384 536
rect 4896 484 4948 536
<< metal2 >>
rect 3882 22536 3938 22545
rect 3882 22471 3938 22480
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2778 21176 2834 21185
rect 2778 21111 2834 21120
rect 1950 20632 2006 20641
rect 1950 20567 2006 20576
rect 1964 20058 1992 20567
rect 2792 20058 2820 21111
rect 2870 20224 2926 20233
rect 2870 20159 2926 20168
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 18766 1808 19858
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2136 19304 2188 19310
rect 1858 19272 1914 19281
rect 2136 19246 2188 19252
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 1858 19207 1914 19216
rect 1872 18970 1900 19207
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1950 18320 2006 18329
rect 2148 18290 2176 19246
rect 2332 18902 2360 19246
rect 2884 19174 2912 20159
rect 3068 19514 3096 22063
rect 3238 21584 3294 21593
rect 3238 21519 3294 21528
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 3252 18426 3280 21519
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 1950 18255 2006 18264
rect 2136 18284 2188 18290
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1872 17814 1900 18158
rect 1964 17882 1992 18255
rect 2136 18226 2188 18232
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 3344 17814 3372 18634
rect 3698 17912 3754 17921
rect 3698 17847 3754 17856
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 1674 17368 1730 17377
rect 1674 17303 1676 17312
rect 1728 17303 1730 17312
rect 1676 17274 1728 17280
rect 2884 17134 2912 17614
rect 3712 17338 3740 17847
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 1504 16726 1532 17070
rect 3792 16992 3844 16998
rect 1858 16960 1914 16969
rect 3792 16934 3844 16940
rect 1858 16895 1914 16904
rect 1872 16794 1900 16895
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 3804 16726 3832 16934
rect 1492 16720 1544 16726
rect 1492 16662 1544 16668
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1688 16114 1716 16594
rect 3332 16584 3384 16590
rect 2962 16552 3018 16561
rect 3332 16526 3384 16532
rect 2962 16487 3018 16496
rect 2976 16250 3004 16487
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3344 16114 3372 16526
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 1492 16040 1544 16046
rect 2044 16040 2096 16046
rect 1492 15982 1544 15988
rect 1674 16008 1730 16017
rect 1504 14414 1532 15982
rect 2044 15982 2096 15988
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 1674 15943 1730 15952
rect 1688 15910 1716 15943
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 2056 15706 2084 15982
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1582 14104 1638 14113
rect 1872 14074 1900 14894
rect 1964 14657 1992 15302
rect 1950 14648 2006 14657
rect 1950 14583 2006 14592
rect 1582 14039 1638 14048
rect 1860 14068 1912 14074
rect 1596 12986 1624 14039
rect 1860 14010 1912 14016
rect 2056 13462 2084 15506
rect 2332 13938 2360 15506
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 15065 2820 15302
rect 2884 15162 2912 15982
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2608 14278 2636 14894
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2700 13938 2728 14894
rect 3344 14618 3372 15438
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6866 1532 7142
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1688 6798 1716 13194
rect 1780 12986 1808 13330
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1780 11898 1808 12378
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 2240 11694 2268 13398
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2332 12442 2360 12582
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11762 2360 12242
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2228 11688 2280 11694
rect 2280 11636 2360 11642
rect 2228 11630 2360 11636
rect 2240 11614 2360 11630
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11354 1900 11494
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8090 1992 8910
rect 2240 8362 2268 9318
rect 2332 9058 2360 11614
rect 2516 10266 2544 13330
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12782 2728 13262
rect 3068 12986 3096 14486
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2792 11694 2820 12310
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2792 11558 2820 11630
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 10606 2820 11494
rect 2884 10674 2912 11630
rect 2976 10810 3004 12582
rect 3160 12442 3188 12786
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3160 11626 3188 12378
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3252 11150 3280 13942
rect 3620 13938 3648 14418
rect 3712 14346 3740 14826
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3436 13530 3464 13631
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3606 13288 3662 13297
rect 3606 13223 3662 13232
rect 3422 12744 3478 12753
rect 3422 12679 3478 12688
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2884 10470 2912 10610
rect 3160 10538 3188 11086
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2424 9178 2452 10066
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2700 9450 2728 9998
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2332 9030 2452 9058
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2134 8256 2190 8265
rect 2134 8191 2190 8200
rect 2148 8090 2176 8191
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 6928 1820 6934
rect 1768 6870 1820 6876
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 4622 1440 6190
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 664 3392 716 3398
rect 664 3334 716 3340
rect 204 2440 256 2446
rect 204 2382 256 2388
rect 216 480 244 2382
rect 676 480 704 3334
rect 1124 2916 1176 2922
rect 1124 2858 1176 2864
rect 1136 480 1164 2858
rect 1504 1057 1532 6598
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 4078 1716 4558
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 3670 1716 4014
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1490 1048 1546 1057
rect 1490 983 1546 992
rect 1596 480 1624 2790
rect 1780 2009 1808 6870
rect 1872 2553 1900 7822
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 1766 2000 1822 2009
rect 1766 1935 1822 1944
rect 1964 1601 1992 7890
rect 2148 6100 2176 8026
rect 2240 6798 2268 8298
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6254 2268 6734
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2148 6072 2268 6100
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4865 2084 4966
rect 2042 4856 2098 4865
rect 2042 4791 2098 4800
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2056 2582 2084 3878
rect 2148 2650 2176 3878
rect 2240 3505 2268 6072
rect 2332 5914 2360 7142
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2424 5710 2452 9030
rect 2700 8634 2728 9386
rect 2976 9178 3004 10066
rect 3160 9654 3188 10474
rect 3344 10198 3372 12242
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3238 10024 3294 10033
rect 3238 9959 3294 9968
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2870 9072 2926 9081
rect 2870 9007 2926 9016
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 6866 2544 7346
rect 2792 7290 2820 7822
rect 2700 7262 2820 7290
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4282 2360 4966
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2226 3496 2282 3505
rect 2226 3431 2282 3440
rect 2424 2961 2452 5646
rect 2516 3890 2544 6054
rect 2700 5794 2728 7262
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 5914 2820 7142
rect 2884 6118 2912 9007
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2700 5766 2912 5794
rect 2976 5778 3004 7142
rect 3252 6662 3280 9959
rect 3436 9738 3464 12679
rect 3620 12442 3648 13223
rect 3804 12918 3832 13738
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3896 12764 3924 22471
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4816 17814 4844 19858
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15502 4016 15914
rect 4724 15910 4752 16662
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4066 15600 4122 15609
rect 4122 15558 4200 15586
rect 4066 15535 4122 15544
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3988 15162 4016 15438
rect 4172 15162 4200 15558
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4816 15026 4844 16934
rect 4908 15706 4936 16934
rect 5092 16794 5120 17138
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5368 16046 5396 16730
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13954 4292 14214
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4264 13926 4384 13954
rect 4356 13870 4384 13926
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4356 13546 4384 13806
rect 5092 13734 5120 14350
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4264 13518 4384 13546
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12986 4200 13330
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3804 12736 3924 12764
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3514 10840 3570 10849
rect 3514 10775 3570 10784
rect 3528 9926 3556 10775
rect 3620 10606 3648 11018
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3436 9710 3648 9738
rect 3712 9722 3740 10406
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3344 8090 3372 8978
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3330 7984 3386 7993
rect 3330 7919 3332 7928
rect 3384 7919 3386 7928
rect 3332 7890 3384 7896
rect 3436 7546 3464 8910
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3528 6882 3556 9415
rect 3620 8514 3648 9710
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3804 9518 3832 12736
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4120 12336 4122 12345
rect 4066 12271 4122 12280
rect 3974 11384 4030 11393
rect 4172 11354 4200 12582
rect 4264 11762 4292 13518
rect 5184 13274 5212 15642
rect 5276 15502 5304 15846
rect 5644 15502 5672 15914
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5644 14482 5672 15438
rect 5736 15162 5764 17206
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6012 15638 6040 16186
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6196 13938 6224 14418
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5736 13530 5764 13806
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5460 13326 5488 13466
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5448 13320 5500 13326
rect 5184 13246 5304 13274
rect 5448 13262 5500 13268
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4356 12442 4384 12650
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4632 12322 4660 12718
rect 5000 12628 5028 12786
rect 5184 12782 5212 13126
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5000 12600 5120 12628
rect 4632 12294 4936 12322
rect 5092 12306 5120 12600
rect 4710 12200 4766 12209
rect 4710 12135 4712 12144
rect 4764 12135 4766 12144
rect 4712 12106 4764 12112
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4724 11880 4752 12106
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4540 11852 4752 11880
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4540 11558 4568 11852
rect 4816 11694 4844 12038
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 3974 11319 4030 11328
rect 4160 11348 4212 11354
rect 3988 11014 4016 11319
rect 4160 11290 4212 11296
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 4068 10464 4120 10470
rect 4066 10432 4068 10441
rect 4120 10432 4122 10441
rect 4066 10367 4122 10376
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 10062 4108 10202
rect 4264 10198 4292 11494
rect 4356 10996 4384 11494
rect 4724 11354 4752 11562
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4816 11234 4844 11630
rect 4908 11354 4936 12294
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11898 5120 12242
rect 5184 12209 5212 12718
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5276 12084 5304 13246
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5184 12056 5304 12084
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4712 11212 4764 11218
rect 4816 11206 4936 11234
rect 4712 11154 4764 11160
rect 4325 10968 4384 10996
rect 4325 10792 4353 10968
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4325 10764 4476 10792
rect 4448 10266 4476 10764
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3712 8634 3740 8910
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3620 8486 3740 8514
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3620 7886 3648 8298
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7410 3648 7822
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7002 3648 7346
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3528 6854 3648 6882
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3344 5914 3372 6666
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 2884 5658 2912 5766
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2884 5630 3004 5658
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4690 2912 5170
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 4282 2912 4626
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2516 3862 2636 3890
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2410 2952 2466 2961
rect 2410 2887 2466 2896
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 1950 1592 2006 1601
rect 1950 1527 2006 1536
rect 2056 480 2084 2042
rect 2516 480 2544 3470
rect 2608 2530 2636 3862
rect 2884 3738 2912 4218
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2792 3398 2820 3606
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2792 2689 2820 2926
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 2778 2680 2834 2689
rect 2778 2615 2834 2624
rect 2608 2502 2820 2530
rect 2792 2378 2820 2502
rect 2884 2446 2912 2751
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2976 2394 3004 5630
rect 3514 5264 3570 5273
rect 3148 5228 3200 5234
rect 3514 5199 3570 5208
rect 3148 5170 3200 5176
rect 3160 4826 3188 5170
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3344 4826 3372 5102
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3160 4010 3188 4762
rect 3528 4758 3556 5199
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3344 2961 3372 4626
rect 3620 4185 3648 6854
rect 3712 5522 3740 8486
rect 3804 8362 3832 9454
rect 4172 9178 4200 10066
rect 4264 9586 4292 10134
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9654 4752 11154
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10538 4844 11086
rect 4908 10606 4936 11206
rect 5184 11082 5212 12056
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 5092 10266 5120 10542
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 7342 3832 8298
rect 3882 8120 3938 8129
rect 4080 8090 4108 9046
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 3882 8055 3938 8064
rect 4068 8084 4120 8090
rect 3896 7546 3924 8055
rect 4068 8026 4120 8032
rect 4264 7750 4292 8502
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 8294 4752 8366
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 7954 4752 8230
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 3974 7576 4030 7585
rect 3884 7540 3936 7546
rect 4388 7568 4684 7588
rect 3974 7511 4030 7520
rect 3884 7482 3936 7488
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3988 7002 4016 7511
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3976 6248 4028 6254
rect 3882 6216 3938 6225
rect 3976 6190 4028 6196
rect 3882 6151 3938 6160
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5710 3832 6054
rect 3896 5846 3924 6151
rect 3884 5840 3936 5846
rect 3988 5817 4016 6190
rect 3884 5782 3936 5788
rect 3974 5808 4030 5817
rect 3974 5743 4030 5752
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3712 5494 3924 5522
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3712 3738 3740 4558
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3436 3126 3464 3538
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3330 2952 3386 2961
rect 3330 2887 3386 2896
rect 3146 2680 3202 2689
rect 3146 2615 3202 2624
rect 3160 2514 3188 2615
rect 3436 2582 3464 3062
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3436 2446 3464 2518
rect 3424 2440 3476 2446
rect 2780 2372 2832 2378
rect 2976 2366 3096 2394
rect 3424 2382 3476 2388
rect 2780 2314 2832 2320
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2976 480 3004 2246
rect 3068 649 3096 2366
rect 3528 2292 3556 3674
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3712 3194 3740 3402
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3712 3058 3740 3130
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3804 2514 3832 5102
rect 3896 4690 3924 5494
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 4080 4146 4108 7142
rect 4724 6798 4752 7686
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4724 6186 4752 6734
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5710 4752 6122
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4172 4026 4200 5646
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 3896 3998 4200 4026
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3436 2264 3556 2292
rect 3054 640 3110 649
rect 3054 575 3110 584
rect 3332 536 3384 542
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 2962 0 3018 480
rect 3332 478 3384 484
rect 3436 480 3464 2264
rect 3896 480 3924 3998
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 4080 3738 4108 3839
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4172 3398 4200 3606
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4160 2644 4212 2650
rect 4080 2604 4160 2632
rect 4080 2106 4108 2604
rect 4160 2586 4212 2592
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4172 2310 4200 2450
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4264 1442 4292 4082
rect 4448 3534 4476 4082
rect 4724 3670 4752 5170
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4724 3194 4752 3606
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 4632 2446 4660 2518
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4384 1442
rect 4356 480 4384 1414
rect 4816 480 4844 9318
rect 4908 6866 4936 9590
rect 5184 9500 5212 11018
rect 5276 9654 5304 11630
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 10266 5488 10474
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 9654 5580 12582
rect 6104 12238 6132 13330
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6092 12232 6144 12238
rect 6012 12180 6092 12186
rect 6012 12174 6144 12180
rect 6012 12158 6132 12174
rect 6012 11694 6040 12158
rect 6092 12096 6144 12102
rect 6196 12084 6224 12650
rect 6144 12056 6224 12084
rect 6092 12038 6144 12044
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5644 10810 5672 11562
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 9586 5672 10746
rect 5736 10266 5764 11222
rect 5828 11218 5856 11562
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5184 9472 5580 9500
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5092 8294 5120 9046
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7342 5120 8230
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 6866 5120 7278
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6458 4936 6598
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4146 4936 4626
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4908 542 4936 3606
rect 5000 2650 5028 4966
rect 5092 4826 5120 4966
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5092 2310 5120 4014
rect 5184 3448 5212 9318
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5276 8974 5304 9046
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8022 5304 8774
rect 5368 8634 5396 8978
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5846 5304 6054
rect 5356 5908 5408 5914
rect 5460 5896 5488 9318
rect 5552 6934 5580 9472
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5644 6186 5672 6938
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5408 5868 5488 5896
rect 5356 5850 5408 5856
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5368 3670 5396 5850
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 4690 5672 5510
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 3942 5580 4558
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5184 3420 5304 3448
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4896 536 4948 542
rect 3344 241 3372 478
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4342 0 4398 480
rect 4802 0 4858 480
rect 4896 478 4948 484
rect 5276 480 5304 3420
rect 5460 3194 5488 3470
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5552 3126 5580 3878
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5552 2922 5580 3062
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2310 5672 2790
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5736 480 5764 9386
rect 5828 8090 5856 11154
rect 6104 11150 6132 12038
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10266 6132 10406
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 8090 6132 8230
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 6662 5948 7210
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6322 5948 6598
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5828 5166 5856 6054
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5828 3466 5856 3946
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3194 6040 3334
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5920 2666 5948 2790
rect 5828 2650 5948 2666
rect 6012 2650 6040 3130
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 5816 2644 5948 2650
rect 5868 2638 5948 2644
rect 6000 2644 6052 2650
rect 5816 2586 5868 2592
rect 6000 2586 6052 2592
rect 6104 2446 6132 3062
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6196 480 6224 11154
rect 6288 10266 6316 17614
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 9042 6316 9522
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8906 6316 8978
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8498 6316 8842
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6380 7562 6408 15506
rect 6472 14958 6500 16390
rect 6656 14958 6684 16594
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 12646 6500 13330
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6564 12374 6592 13874
rect 6656 12866 6684 14894
rect 6748 12986 6776 17002
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 14890 6868 15846
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6656 12838 6776 12866
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11558 6500 12242
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 12102 6592 12174
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6380 7534 6592 7562
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6934 6500 7142
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6472 5710 6500 6870
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 2825 6316 4966
rect 6380 4690 6408 5170
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4214 6408 4626
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 3670 6500 5238
rect 6564 3670 6592 7534
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 6656 480 6684 12582
rect 6748 12288 6776 12838
rect 6748 12260 6868 12288
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 11218 6776 12106
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6840 10062 6868 12260
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6932 8090 6960 16594
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7024 16250 7052 16526
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7116 15026 7144 15302
rect 7208 15162 7236 18906
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8312 17814 8340 18158
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 16794 7788 17682
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7484 15502 7512 15982
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14550 7144 14962
rect 7484 14618 7512 15438
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 12628 7144 14214
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 12782 7236 13670
rect 7564 13524 7616 13530
rect 7668 13512 7696 15302
rect 7760 15026 7788 15506
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14618 8248 14894
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7760 13802 7788 14282
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7616 13484 7696 13512
rect 7564 13466 7616 13472
rect 7760 13326 7788 13738
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12850 7328 13126
rect 8220 12850 8248 13670
rect 8312 13530 8340 14486
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13258 8432 18770
rect 10612 18290 10640 19246
rect 17866 19136 17922 19145
rect 14684 19068 14980 19088
rect 17866 19071 17922 19080
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8588 14618 8616 14758
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7116 12600 7328 12628
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 10266 7052 11494
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7116 10146 7144 11698
rect 7024 10118 7144 10146
rect 7024 9994 7052 10118
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7024 8294 7052 9930
rect 7116 8566 7144 9998
rect 7300 9636 7328 12600
rect 7484 12374 7512 12786
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 10674 7420 11494
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 8128 10606 8156 10950
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 7576 10062 7604 10542
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7300 9608 7420 9636
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7392 8634 7420 9608
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7576 9178 7604 9318
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7668 8634 7696 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 9110 8248 12650
rect 8404 12442 8432 12922
rect 8496 12646 8524 13330
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8312 11898 8340 12174
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8496 11694 8524 12582
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10266 8432 10950
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7012 8288 7064 8294
rect 7010 8256 7012 8265
rect 7064 8256 7066 8265
rect 7010 8191 7066 8200
rect 7208 8106 7236 8570
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7116 8078 7236 8106
rect 7392 8090 7420 8366
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7288 8084 7340 8090
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 5302 6868 7822
rect 6932 6390 6960 7890
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 5778 7052 6258
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5302 6960 5510
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7024 5234 7052 5714
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4282 6868 5102
rect 7024 4826 7052 5170
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 2514 6776 4014
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 3194 6868 3402
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6932 2650 6960 2858
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7024 2514 7052 3538
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6748 2417 6776 2450
rect 6734 2408 6790 2417
rect 6734 2343 6790 2352
rect 7116 480 7144 8078
rect 7288 8026 7340 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7208 5846 7236 7958
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7208 3602 7236 5238
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7208 2582 7236 3130
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7300 1426 7328 8026
rect 8220 7993 8248 9046
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8498 8524 8774
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8206 7984 8262 7993
rect 8206 7919 8262 7928
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7392 3058 7420 3538
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7484 2650 7512 7278
rect 7668 6934 7696 7346
rect 7760 7206 7788 7482
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7838 6760 7894 6769
rect 7838 6695 7894 6704
rect 7852 6186 7880 6695
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7760 5234 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 8220 5030 8248 6802
rect 8404 6322 8432 7278
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8404 5234 8432 6258
rect 8496 5914 8524 7822
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8496 5098 8524 5850
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8220 4282 8248 4558
rect 8312 4282 8340 4694
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8312 4146 8340 4218
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 4072 8260 4078
rect 8206 4040 8208 4049
rect 8260 4040 8262 4049
rect 8206 3975 8262 3984
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7484 2310 7512 2586
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7288 1420 7340 1426
rect 7288 1362 7340 1368
rect 7576 480 7604 3606
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7654 2408 7710 2417
rect 7654 2343 7710 2352
rect 7668 2310 7696 2343
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 8128 480 8156 1362
rect 8588 480 8616 13398
rect 8680 12986 8708 18090
rect 11072 17882 11100 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8864 15706 8892 15914
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8864 12714 8892 14350
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8852 11756 8904 11762
rect 8956 11744 8984 12038
rect 8904 11716 8984 11744
rect 8852 11698 8904 11704
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8680 9178 8708 11562
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 11354 8800 11494
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8956 11286 8984 11716
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8772 8362 8800 11154
rect 8956 11150 8984 11222
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8864 7562 8892 11086
rect 9048 10266 9076 17614
rect 10336 17338 10364 17682
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9140 16590 9168 17002
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16250 9168 16526
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9600 15706 9628 16662
rect 9784 16658 9812 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 16114 9812 16594
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9784 14958 9812 16050
rect 10060 15978 10088 16934
rect 10704 16794 10732 16934
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10060 15026 10088 15914
rect 10796 15162 10824 16934
rect 11164 16658 11192 17138
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11164 16250 11192 16594
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11624 15706 11652 17750
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 16794 13676 17614
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 17880 16794 17908 19071
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11164 15366 11192 15642
rect 12084 15502 12112 16662
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9324 14414 9352 14826
rect 9784 14618 9812 14894
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9324 14074 9352 14350
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9232 13326 9260 13738
rect 9692 13530 9720 14350
rect 9784 13870 9812 14554
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9784 13394 9812 13806
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12238 9260 12650
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11898 9260 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11694 9352 12718
rect 9692 12442 9720 13126
rect 9784 12782 9812 13330
rect 9968 12986 9996 13330
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9968 12374 9996 12922
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9600 11286 9628 11727
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9680 11144 9732 11150
rect 9784 11098 9812 11494
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9732 11092 9812 11098
rect 9680 11086 9812 11092
rect 9692 11070 9812 11086
rect 9784 10810 9812 11070
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9722 9076 9998
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9324 9586 9352 10474
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 8864 7534 9076 7562
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 7002 8800 7142
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8956 6730 8984 7346
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6254 8984 6666
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 4146 8984 4558
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8864 3602 8892 4082
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8864 3126 8892 3538
rect 8956 3398 8984 4082
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8864 2446 8892 3062
rect 8956 2990 8984 3334
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9048 480 9076 7534
rect 9126 6896 9182 6905
rect 9126 6831 9182 6840
rect 9140 6254 9168 6831
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9416 4706 9444 9318
rect 9586 8528 9642 8537
rect 9586 8463 9642 8472
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9600 8242 9628 8463
rect 9692 8430 9720 10542
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8498 9812 8978
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9508 8022 9536 8230
rect 9600 8214 9720 8242
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9128 4684 9180 4690
rect 9416 4678 9536 4706
rect 9128 4626 9180 4632
rect 9140 3670 9168 4626
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 2854 9168 3470
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9232 2650 9260 3878
rect 9324 3194 9352 3878
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9508 480 9536 4678
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 2854 9628 4422
rect 9692 3942 9720 8214
rect 9784 6798 9812 8434
rect 9968 7834 9996 11290
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 8090 10088 9862
rect 10336 9160 10364 12106
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10470 10456 11154
rect 10796 10810 10824 12582
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10062 10456 10406
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10336 9132 10456 9160
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 9968 7806 10088 7834
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7274 9996 7686
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 6390 9996 6734
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 4690 9812 6054
rect 9968 5914 9996 6326
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9968 5234 9996 5850
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9968 4826 9996 5170
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9968 4146 9996 4762
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9692 3097 9720 3470
rect 9678 3088 9734 3097
rect 9784 3058 9812 3946
rect 9968 3670 9996 4082
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10060 3516 10088 7806
rect 10244 6118 10272 7890
rect 10336 7886 10364 8978
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10152 5914 10180 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10138 5808 10194 5817
rect 10138 5743 10194 5752
rect 10152 5574 10180 5743
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9968 3488 10088 3516
rect 9678 3023 9734 3032
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9588 2848 9640 2854
rect 9876 2825 9904 2926
rect 9588 2790 9640 2796
rect 9862 2816 9918 2825
rect 9862 2751 9918 2760
rect 9968 480 9996 3488
rect 10152 2650 10180 3878
rect 10244 3602 10272 6054
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10336 2446 10364 4626
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10428 480 10456 9132
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10520 6254 10548 6938
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10612 4078 10640 10066
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8634 10732 8842
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8634 10824 8774
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 6361 10732 7278
rect 10690 6352 10746 6361
rect 10690 6287 10692 6296
rect 10744 6287 10746 6296
rect 10692 6258 10744 6264
rect 10784 5704 10836 5710
rect 10782 5672 10784 5681
rect 10836 5672 10838 5681
rect 10782 5607 10838 5616
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10888 480 10916 14282
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11354 11100 11562
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10606 11100 10950
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10980 10266 11008 10542
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8362 11100 8774
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7818 11100 8298
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10980 6934 11008 7142
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10980 5710 11008 6870
rect 11072 5914 11100 7142
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4010 11100 4422
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11072 3058 11100 3946
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10980 2378 11008 2518
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11164 1442 11192 15302
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 8090 11468 8230
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5710 11284 6326
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11624 4434 11652 14758
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11354 11744 12038
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 6254 11836 6734
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5370 11836 5782
rect 11992 5778 12020 7686
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11716 5030 11744 5238
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11808 4604 11836 5306
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4826 11928 4966
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11888 4616 11940 4622
rect 11808 4576 11888 4604
rect 11888 4558 11940 4564
rect 11624 4406 11744 4434
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3602 11652 3878
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11426 3088 11482 3097
rect 11426 3023 11482 3032
rect 11440 2854 11468 3023
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11532 2378 11560 2790
rect 11624 2446 11652 3538
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11520 2372 11572 2378
rect 11520 2314 11572 2320
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1414 11376 1442
rect 11348 480 11376 1414
rect 11716 1034 11744 4406
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 2922 11928 3878
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11808 2514 11836 2858
rect 11992 2514 12020 5170
rect 12164 4072 12216 4078
rect 12162 4040 12164 4049
rect 12216 4040 12218 4049
rect 12162 3975 12218 3984
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12084 3058 12112 3606
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11716 1006 11836 1034
rect 11808 480 11836 1006
rect 12268 480 12296 15506
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19890 11520 19946 11529
rect 14684 11452 14980 11472
rect 19890 11455 19946 11464
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12348 11144 12400 11150
rect 12452 11098 12480 11154
rect 12400 11092 12480 11098
rect 12348 11086 12480 11092
rect 12360 11070 12480 11086
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7342 12388 7890
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 6254 12388 7278
rect 12544 7002 12572 10474
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12452 5710 12480 6394
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12544 5166 12572 5607
rect 12636 5370 12664 7210
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 2825 12664 5034
rect 12622 2816 12678 2825
rect 12622 2751 12678 2760
rect 12728 480 12756 8842
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13832 7546 13860 7890
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13832 7410 13860 7482
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12820 6934 12848 7210
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 13004 6730 13032 7210
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 16500 6866 16528 7414
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5914 12848 6122
rect 13188 6118 13216 6734
rect 13832 6458 13860 6802
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13188 5574 13216 6054
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13096 4690 13124 5306
rect 13924 5166 13952 6054
rect 14384 5574 14412 6734
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6361 14596 6598
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5914 14504 6054
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 15120 5642 15148 6190
rect 15856 5817 15884 6190
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15842 5808 15898 5817
rect 15842 5743 15898 5752
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 14384 5166 14412 5510
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13174 4176 13230 4185
rect 13174 4111 13230 4120
rect 13452 4140 13504 4146
rect 13188 4010 13216 4111
rect 13452 4082 13504 4088
rect 13358 4040 13414 4049
rect 13176 4004 13228 4010
rect 13358 3975 13360 3984
rect 13176 3946 13228 3952
rect 13412 3975 13414 3984
rect 13360 3946 13412 3952
rect 13464 3670 13492 4082
rect 14384 4078 14412 5102
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15304 4826 15332 5510
rect 15856 5098 15884 5646
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 13544 4072 13596 4078
rect 14372 4072 14424 4078
rect 13544 4014 13596 4020
rect 14370 4040 14372 4049
rect 14424 4040 14426 4049
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13452 3528 13504 3534
rect 13556 3516 13584 4014
rect 14370 3975 14426 3984
rect 13504 3488 13584 3516
rect 13452 3470 13504 3476
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 2990 13492 3334
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 12912 2650 12940 2790
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13188 480 13216 2246
rect 13648 480 13676 2790
rect 13924 2514 13952 2858
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14200 2446 14228 2926
rect 14476 2514 14504 4558
rect 14568 2990 14596 4694
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15028 3466 15056 3946
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15396 2990 15424 3334
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 480 14136 2246
rect 14568 480 14596 2790
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15488 2514 15516 4966
rect 15856 4554 15884 5034
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 4214 15884 4490
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3602 15792 3878
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15948 3058 15976 3946
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16040 2514 16068 6122
rect 16132 5370 16160 6802
rect 16592 6254 16620 7278
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17696 6254 17724 6734
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16316 5778 16344 6122
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16132 4622 16160 5306
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3738 16160 3878
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16316 3194 16344 3538
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 15028 480 15056 2246
rect 15580 480 15608 2246
rect 16040 480 16068 2246
rect 16500 480 16528 5510
rect 16592 5234 16620 5782
rect 16868 5778 16896 6122
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16684 4282 16712 4626
rect 16776 4622 16804 5102
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16776 3738 16804 4558
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 2514 16620 3470
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16960 480 16988 5510
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 4078 17080 4422
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17040 4072 17092 4078
rect 17132 4072 17184 4078
rect 17040 4014 17092 4020
rect 17130 4040 17132 4049
rect 17184 4040 17186 4049
rect 17130 3975 17186 3984
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17972 3602 18000 3946
rect 18064 3913 18092 4082
rect 18050 3904 18106 3913
rect 18050 3839 18106 3848
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18708 2990 18736 7822
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17144 2514 17172 2858
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 480 17448 2314
rect 17880 480 17908 2790
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18368 1170
rect 18340 480 18368 1142
rect 18800 480 18828 3334
rect 19260 480 19288 6054
rect 19904 4078 19932 11455
rect 20272 11354 20300 11630
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 480 19748 2790
rect 20180 480 20208 10406
rect 20350 2952 20406 2961
rect 20350 2887 20352 2896
rect 20404 2887 20406 2896
rect 20352 2858 20404 2864
rect 20640 480 20668 11018
rect 20916 626 20944 11494
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 20916 598 21128 626
rect 21100 480 21128 598
rect 21560 480 21588 2790
rect 22020 480 22048 3334
rect 22480 480 22508 3674
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9034 0 9090 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15566 0 15622 480
rect 16026 0 16082 480
rect 16486 0 16542 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18326 0 18382 480
rect 18786 0 18842 480
rect 19246 0 19302 480
rect 19706 0 19762 480
rect 20166 0 20222 480
rect 20626 0 20682 480
rect 21086 0 21142 480
rect 21546 0 21602 480
rect 22006 0 22062 480
rect 22466 0 22522 480
<< via2 >>
rect 3882 22480 3938 22536
rect 3054 22072 3110 22128
rect 2778 21120 2834 21176
rect 1950 20576 2006 20632
rect 2870 20168 2926 20224
rect 1950 19760 2006 19816
rect 1858 19216 1914 19272
rect 1950 18808 2006 18864
rect 1950 18264 2006 18320
rect 3238 21528 3294 21584
rect 3698 17856 3754 17912
rect 1674 17332 1730 17368
rect 1674 17312 1676 17332
rect 1676 17312 1728 17332
rect 1728 17312 1730 17332
rect 1858 16904 1914 16960
rect 2962 16496 3018 16552
rect 1674 15952 1730 16008
rect 1582 14048 1638 14104
rect 1950 14592 2006 14648
rect 2778 15000 2834 15056
rect 3422 13640 3478 13696
rect 3606 13232 3662 13288
rect 3422 12688 3478 12744
rect 2134 8200 2190 8256
rect 1490 992 1546 1048
rect 1858 2488 1914 2544
rect 1766 1944 1822 2000
rect 2042 4800 2098 4856
rect 3238 9968 3294 10024
rect 2870 9016 2926 9072
rect 2226 3440 2282 3496
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4066 15544 4122 15600
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3514 10784 3570 10840
rect 3514 9424 3570 9480
rect 3330 7948 3386 7984
rect 3330 7928 3332 7948
rect 3332 7928 3384 7948
rect 3384 7928 3386 7948
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 3974 11328 4030 11384
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4710 12164 4766 12200
rect 4710 12144 4712 12164
rect 4712 12144 4764 12164
rect 4764 12144 4766 12164
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 10412 4068 10432
rect 4068 10412 4120 10432
rect 4120 10412 4122 10432
rect 4066 10376 4122 10412
rect 5170 12144 5226 12200
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 2410 2896 2466 2952
rect 1950 1536 2006 1592
rect 2870 2760 2926 2816
rect 2778 2624 2834 2680
rect 3514 5208 3570 5264
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3882 8064 3938 8120
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 3974 7520 4030 7576
rect 3882 6160 3938 6216
rect 3974 5752 4030 5808
rect 3606 4120 3662 4176
rect 3330 2896 3386 2952
rect 3146 2624 3202 2680
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 3054 584 3110 640
rect 4066 3848 4122 3904
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 3330 176 3386 232
rect 6274 2760 6330 2816
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 17866 19080 17922 19136
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7010 8236 7012 8256
rect 7012 8236 7064 8256
rect 7064 8236 7066 8256
rect 7010 8200 7066 8236
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 6734 2352 6790 2408
rect 8206 7928 8262 7984
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7838 6704 7894 6760
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 8206 4020 8208 4040
rect 8208 4020 8260 4040
rect 8260 4020 8262 4040
rect 8206 3984 8262 4020
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 7654 2352 7710 2408
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 9586 11736 9642 11792
rect 9126 6840 9182 6896
rect 9586 8472 9642 8528
rect 9678 3032 9734 3088
rect 10138 5752 10194 5808
rect 9862 2760 9918 2816
rect 10690 6316 10746 6352
rect 10690 6296 10692 6316
rect 10692 6296 10744 6316
rect 10744 6296 10746 6316
rect 10782 5652 10784 5672
rect 10784 5652 10836 5672
rect 10836 5652 10838 5672
rect 10782 5616 10838 5652
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11426 3032 11482 3088
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12162 4020 12164 4040
rect 12164 4020 12216 4040
rect 12216 4020 12218 4040
rect 12162 3984 12218 4020
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 19890 11464 19946 11520
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 12530 5616 12586 5672
rect 12622 2760 12678 2816
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14554 6296 14610 6352
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15842 5752 15898 5808
rect 13174 4120 13230 4176
rect 13358 4004 13414 4040
rect 13358 3984 13360 4004
rect 13360 3984 13412 4004
rect 13412 3984 13414 4004
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14370 4020 14372 4040
rect 14372 4020 14424 4040
rect 14424 4020 14426 4040
rect 14370 3984 14426 4020
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17130 4020 17132 4040
rect 17132 4020 17184 4040
rect 17184 4020 17186 4040
rect 17130 3984 17186 4020
rect 18050 3848 18106 3904
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 20350 2916 20406 2952
rect 20350 2896 20352 2916
rect 20352 2896 20404 2916
rect 20404 2896 20406 2916
<< metal3 >>
rect 0 22538 480 22568
rect 3877 22538 3943 22541
rect 0 22536 3943 22538
rect 0 22480 3882 22536
rect 3938 22480 3943 22536
rect 0 22478 3943 22480
rect 0 22448 480 22478
rect 3877 22475 3943 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 0 21586 480 21616
rect 3233 21586 3299 21589
rect 0 21584 3299 21586
rect 0 21528 3238 21584
rect 3294 21528 3299 21584
rect 0 21526 3299 21528
rect 0 21496 480 21526
rect 3233 21523 3299 21526
rect 0 21178 480 21208
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 480 21118
rect 2773 21115 2839 21118
rect 0 20634 480 20664
rect 1945 20634 2011 20637
rect 0 20632 2011 20634
rect 0 20576 1950 20632
rect 2006 20576 2011 20632
rect 0 20574 2011 20576
rect 0 20544 480 20574
rect 1945 20571 2011 20574
rect 0 20226 480 20256
rect 2865 20226 2931 20229
rect 0 20224 2931 20226
rect 0 20168 2870 20224
rect 2926 20168 2931 20224
rect 0 20166 2931 20168
rect 0 20136 480 20166
rect 2865 20163 2931 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1853 19274 1919 19277
rect 0 19272 1919 19274
rect 0 19216 1858 19272
rect 1914 19216 1919 19272
rect 0 19214 1919 19216
rect 0 19184 480 19214
rect 1853 19211 1919 19214
rect 17861 19138 17927 19141
rect 22320 19138 22800 19168
rect 17861 19136 22800 19138
rect 17861 19080 17866 19136
rect 17922 19080 22800 19136
rect 17861 19078 22800 19080
rect 17861 19075 17927 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 22320 19048 22800 19078
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 480 18262
rect 1945 18259 2011 18262
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 3693 17914 3759 17917
rect 0 17912 3759 17914
rect 0 17856 3698 17912
rect 3754 17856 3759 17912
rect 0 17854 3759 17856
rect 0 17824 480 17854
rect 3693 17851 3759 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1669 17370 1735 17373
rect 0 17368 1735 17370
rect 0 17312 1674 17368
rect 1730 17312 1735 17368
rect 0 17310 1735 17312
rect 0 17280 480 17310
rect 1669 17307 1735 17310
rect 0 16962 480 16992
rect 1853 16962 1919 16965
rect 0 16960 1919 16962
rect 0 16904 1858 16960
rect 1914 16904 1919 16960
rect 0 16902 1919 16904
rect 0 16872 480 16902
rect 1853 16899 1919 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 2957 16554 3023 16557
rect 0 16552 3023 16554
rect 0 16496 2962 16552
rect 3018 16496 3023 16552
rect 0 16494 3023 16496
rect 0 16464 480 16494
rect 2957 16491 3023 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1669 16010 1735 16013
rect 0 16008 1735 16010
rect 0 15952 1674 16008
rect 1730 15952 1735 16008
rect 0 15950 1735 15952
rect 0 15920 480 15950
rect 1669 15947 1735 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 4061 15602 4127 15605
rect 0 15600 4127 15602
rect 0 15544 4066 15600
rect 4122 15544 4127 15600
rect 0 15542 4127 15544
rect 0 15512 480 15542
rect 4061 15539 4127 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 480 14998
rect 2773 14995 2839 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1945 14650 2011 14653
rect 0 14648 2011 14650
rect 0 14592 1950 14648
rect 2006 14592 2011 14648
rect 0 14590 2011 14592
rect 0 14560 480 14590
rect 1945 14587 2011 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 480 14046
rect 1577 14043 1643 14046
rect 0 13698 480 13728
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13608 480 13638
rect 3417 13635 3483 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 3601 13290 3667 13293
rect 0 13288 3667 13290
rect 0 13232 3606 13288
rect 3662 13232 3667 13288
rect 0 13230 3667 13232
rect 0 13200 480 13230
rect 3601 13227 3667 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 3417 12746 3483 12749
rect 0 12744 3483 12746
rect 0 12688 3422 12744
rect 3478 12688 3483 12744
rect 0 12686 3483 12688
rect 0 12656 480 12686
rect 3417 12683 3483 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 4705 12202 4771 12205
rect 5165 12202 5231 12205
rect 4705 12200 5231 12202
rect 4705 12144 4710 12200
rect 4766 12144 5170 12200
rect 5226 12144 5231 12200
rect 4705 12142 5231 12144
rect 4705 12139 4771 12142
rect 5165 12139 5231 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 9581 11794 9647 11797
rect 0 11792 9647 11794
rect 0 11736 9586 11792
rect 9642 11736 9647 11792
rect 0 11734 9647 11736
rect 0 11704 480 11734
rect 9581 11731 9647 11734
rect 19885 11522 19951 11525
rect 22320 11522 22800 11552
rect 19885 11520 22800 11522
rect 19885 11464 19890 11520
rect 19946 11464 22800 11520
rect 19885 11462 22800 11464
rect 19885 11459 19951 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22320 11432 22800 11462
rect 14672 11391 14992 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 480 11326
rect 3969 11323 4035 11326
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3509 10842 3575 10845
rect 0 10840 3575 10842
rect 0 10784 3514 10840
rect 3570 10784 3575 10840
rect 0 10782 3575 10784
rect 0 10752 480 10782
rect 3509 10779 3575 10782
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10026 480 10056
rect 3233 10026 3299 10029
rect 0 10024 3299 10026
rect 0 9968 3238 10024
rect 3294 9968 3299 10024
rect 0 9966 3299 9968
rect 0 9936 480 9966
rect 3233 9963 3299 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 0 9482 480 9512
rect 3509 9482 3575 9485
rect 0 9480 3575 9482
rect 0 9424 3514 9480
rect 3570 9424 3575 9480
rect 0 9422 3575 9424
rect 0 9392 480 9422
rect 3509 9419 3575 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 2865 9074 2931 9077
rect 0 9072 2931 9074
rect 0 9016 2870 9072
rect 2926 9016 2931 9072
rect 0 9014 2931 9016
rect 0 8984 480 9014
rect 2865 9011 2931 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 9581 8530 9647 8533
rect 0 8528 9647 8530
rect 0 8472 9586 8528
rect 9642 8472 9647 8528
rect 0 8470 9647 8472
rect 0 8440 480 8470
rect 9581 8467 9647 8470
rect 2129 8258 2195 8261
rect 7005 8258 7071 8261
rect 2129 8256 7071 8258
rect 2129 8200 2134 8256
rect 2190 8200 7010 8256
rect 7066 8200 7071 8256
rect 2129 8198 7071 8200
rect 2129 8195 2195 8198
rect 7005 8195 7071 8198
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 3877 8122 3943 8125
rect 0 8120 3943 8122
rect 0 8064 3882 8120
rect 3938 8064 3943 8120
rect 0 8062 3943 8064
rect 0 8032 480 8062
rect 3877 8059 3943 8062
rect 3325 7986 3391 7989
rect 8201 7986 8267 7989
rect 3325 7984 8267 7986
rect 3325 7928 3330 7984
rect 3386 7928 8206 7984
rect 8262 7928 8267 7984
rect 3325 7926 8267 7928
rect 3325 7923 3391 7926
rect 8201 7923 8267 7926
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3969 7578 4035 7581
rect 0 7576 4035 7578
rect 0 7520 3974 7576
rect 4030 7520 4035 7576
rect 0 7518 4035 7520
rect 0 7488 480 7518
rect 3969 7515 4035 7518
rect 0 7170 480 7200
rect 0 7110 4906 7170
rect 0 7080 480 7110
rect 4846 6898 4906 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 9121 6898 9187 6901
rect 4846 6896 9187 6898
rect 4846 6840 9126 6896
rect 9182 6840 9187 6896
rect 4846 6838 9187 6840
rect 9121 6835 9187 6838
rect 0 6762 480 6792
rect 7833 6762 7899 6765
rect 0 6760 7899 6762
rect 0 6704 7838 6760
rect 7894 6704 7899 6760
rect 0 6702 7899 6704
rect 0 6672 480 6702
rect 7833 6699 7899 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 10685 6354 10751 6357
rect 14549 6354 14615 6357
rect 10685 6352 14615 6354
rect 10685 6296 10690 6352
rect 10746 6296 14554 6352
rect 14610 6296 14615 6352
rect 10685 6294 14615 6296
rect 10685 6291 10751 6294
rect 14549 6291 14615 6294
rect 0 6218 480 6248
rect 3877 6218 3943 6221
rect 0 6216 3943 6218
rect 0 6160 3882 6216
rect 3938 6160 3943 6216
rect 0 6158 3943 6160
rect 0 6128 480 6158
rect 3877 6155 3943 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 3969 5810 4035 5813
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 0 5720 480 5750
rect 3969 5747 4035 5750
rect 10133 5810 10199 5813
rect 15837 5810 15903 5813
rect 10133 5808 15903 5810
rect 10133 5752 10138 5808
rect 10194 5752 15842 5808
rect 15898 5752 15903 5808
rect 10133 5750 15903 5752
rect 10133 5747 10199 5750
rect 15837 5747 15903 5750
rect 10777 5674 10843 5677
rect 12525 5674 12591 5677
rect 10777 5672 12591 5674
rect 10777 5616 10782 5672
rect 10838 5616 12530 5672
rect 12586 5616 12591 5672
rect 10777 5614 12591 5616
rect 10777 5611 10843 5614
rect 12525 5611 12591 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 3509 5266 3575 5269
rect 0 5264 3575 5266
rect 0 5208 3514 5264
rect 3570 5208 3575 5264
rect 0 5206 3575 5208
rect 0 5176 480 5206
rect 3509 5203 3575 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 2037 4858 2103 4861
rect 0 4856 2103 4858
rect 0 4800 2042 4856
rect 2098 4800 2103 4856
rect 0 4798 2103 4800
rect 0 4768 480 4798
rect 2037 4795 2103 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 0 4254 3434 4314
rect 0 4224 480 4254
rect 3374 4042 3434 4254
rect 3601 4178 3667 4181
rect 13169 4178 13235 4181
rect 3601 4176 13235 4178
rect 3601 4120 3606 4176
rect 3662 4120 13174 4176
rect 13230 4120 13235 4176
rect 3601 4118 13235 4120
rect 3601 4115 3667 4118
rect 13169 4115 13235 4118
rect 8201 4042 8267 4045
rect 3374 4040 8267 4042
rect 3374 3984 8206 4040
rect 8262 3984 8267 4040
rect 3374 3982 8267 3984
rect 8201 3979 8267 3982
rect 12157 4042 12223 4045
rect 13353 4042 13419 4045
rect 12157 4040 13419 4042
rect 12157 3984 12162 4040
rect 12218 3984 13358 4040
rect 13414 3984 13419 4040
rect 12157 3982 13419 3984
rect 12157 3979 12223 3982
rect 13353 3979 13419 3982
rect 14365 4042 14431 4045
rect 17125 4042 17191 4045
rect 14365 4040 17191 4042
rect 14365 3984 14370 4040
rect 14426 3984 17130 4040
rect 17186 3984 17191 4040
rect 14365 3982 17191 3984
rect 14365 3979 14431 3982
rect 17125 3979 17191 3982
rect 0 3906 480 3936
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 480 3846
rect 4061 3843 4127 3846
rect 18045 3906 18111 3909
rect 22320 3906 22800 3936
rect 18045 3904 22800 3906
rect 18045 3848 18050 3904
rect 18106 3848 22800 3904
rect 18045 3846 22800 3848
rect 18045 3843 18111 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 2221 3498 2287 3501
rect 0 3496 2287 3498
rect 0 3440 2226 3496
rect 2282 3440 2287 3496
rect 0 3438 2287 3440
rect 0 3408 480 3438
rect 2221 3435 2287 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 9673 3090 9739 3093
rect 11421 3090 11487 3093
rect 9673 3088 11487 3090
rect 9673 3032 9678 3088
rect 9734 3032 11426 3088
rect 11482 3032 11487 3088
rect 9673 3030 11487 3032
rect 9673 3027 9739 3030
rect 11421 3027 11487 3030
rect 0 2954 480 2984
rect 2405 2954 2471 2957
rect 0 2952 2471 2954
rect 0 2896 2410 2952
rect 2466 2896 2471 2952
rect 0 2894 2471 2896
rect 0 2864 480 2894
rect 2405 2891 2471 2894
rect 3325 2954 3391 2957
rect 20345 2954 20411 2957
rect 3325 2952 20411 2954
rect 3325 2896 3330 2952
rect 3386 2896 20350 2952
rect 20406 2896 20411 2952
rect 3325 2894 20411 2896
rect 3325 2891 3391 2894
rect 20345 2891 20411 2894
rect 2865 2818 2931 2821
rect 6269 2818 6335 2821
rect 2865 2816 6335 2818
rect 2865 2760 2870 2816
rect 2926 2760 6274 2816
rect 6330 2760 6335 2816
rect 2865 2758 6335 2760
rect 2865 2755 2931 2758
rect 6269 2755 6335 2758
rect 9857 2818 9923 2821
rect 12617 2818 12683 2821
rect 9857 2816 12683 2818
rect 9857 2760 9862 2816
rect 9918 2760 12622 2816
rect 12678 2760 12683 2816
rect 9857 2758 12683 2760
rect 9857 2755 9923 2758
rect 12617 2755 12683 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 2773 2682 2839 2685
rect 3141 2682 3207 2685
rect 2773 2680 3207 2682
rect 2773 2624 2778 2680
rect 2834 2624 3146 2680
rect 3202 2624 3207 2680
rect 2773 2622 3207 2624
rect 2773 2619 2839 2622
rect 3141 2619 3207 2622
rect 0 2546 480 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 480 2486
rect 1853 2483 1919 2486
rect 6729 2410 6795 2413
rect 7649 2410 7715 2413
rect 6729 2408 7715 2410
rect 6729 2352 6734 2408
rect 6790 2352 7654 2408
rect 7710 2352 7715 2408
rect 6729 2350 7715 2352
rect 6729 2347 6795 2350
rect 7649 2347 7715 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 1761 2002 1827 2005
rect 0 2000 1827 2002
rect 0 1944 1766 2000
rect 1822 1944 1827 2000
rect 0 1942 1827 1944
rect 0 1912 480 1942
rect 1761 1939 1827 1942
rect 0 1594 480 1624
rect 1945 1594 2011 1597
rect 0 1592 2011 1594
rect 0 1536 1950 1592
rect 2006 1536 2011 1592
rect 0 1534 2011 1536
rect 0 1504 480 1534
rect 1945 1531 2011 1534
rect 0 1050 480 1080
rect 1485 1050 1551 1053
rect 0 1048 1551 1050
rect 0 992 1490 1048
rect 1546 992 1551 1048
rect 0 990 1551 992
rect 0 960 480 990
rect 1485 987 1551 990
rect 0 642 480 672
rect 3049 642 3115 645
rect 0 640 3115 642
rect 0 584 3054 640
rect 3110 584 3115 640
rect 0 582 3115 584
rect 0 552 480 582
rect 3049 579 3115 582
rect 0 234 480 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 480 174
rect 3325 171 3391 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2024 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1605641404
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1932 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3772 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1605641404
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_26
timestamp 1605641404
transform 1 0 3496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1605641404
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46
timestamp 1605641404
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5428 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5612 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _069_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1605641404
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1605641404
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7360 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp 1605641404
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10028 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84
timestamp 1605641404
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1605641404
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1605641404
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_95
timestamp 1605641404
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1605641404
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1605641404
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11040 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1605641404
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1605641404
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1605641404
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1605641404
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 14444 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp 1605641404
transform 1 0 15088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1605641404
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15364 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1605641404
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1605641404
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1605641404
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16100 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_177
timestamp 1605641404
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1605641404
transform 1 0 16652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1605641404
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_184
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1605641404
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 18768 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1605641404
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1605641404
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1605641404
transform 1 0 20240 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1605641404
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1605641404
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1605641404
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1472 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1605641404
transform 1 0 2944 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4416 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1605641404
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6072 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1605641404
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7452 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1605641404
transform 1 0 6900 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1605641404
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10120 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1605641404
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_96
timestamp 1605641404
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11776 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_114
timestamp 1605641404
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13432 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1605641404
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16284 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1605641404
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1605641404
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 17940 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1605641404
transform 1 0 16836 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_187
timestamp 1605641404
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 20240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_199
timestamp 1605641404
transform 1 0 19412 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_207
timestamp 1605641404
transform 1 0 20148 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1605641404
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2668 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_33
timestamp 1605641404
transform 1 0 4140 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1605641404
transform 1 0 4876 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4968 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1605641404
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7820 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1605641404
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1605641404
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10028 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1605641404
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1605641404
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1605641404
transform 1 0 11500 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1605641404
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14444 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_136
timestamp 1605641404
transform 1 0 13616 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_144
timestamp 1605641404
transform 1 0 14352 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1605641404
transform 1 0 16100 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_161
timestamp 1605641404
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_166
timestamp 1605641404
transform 1 0 16376 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp 1605641404
transform 1 0 16928 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1605641404
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19596 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1605641404
transform 1 0 19136 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_200
timestamp 1605641404
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1605641404
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1656 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1605641404
transform 1 0 3312 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1605641404
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1605641404
transform 1 0 4876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5612 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_65
timestamp 1605641404
transform 1 0 7084 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1605641404
transform 1 0 7636 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1605641404
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1605641404
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 12420 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 1605641404
transform 1 0 11132 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1605641404
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13064 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13800 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_126
timestamp 1605641404
transform 1 0 12696 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1605641404
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_144
timestamp 1605641404
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1605641404
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_174
timestamp 1605641404
transform 1 0 17112 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_186
timestamp 1605641404
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_198
timestamp 1605641404
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1605641404
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1564 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_14
timestamp 1605641404
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_25
timestamp 1605641404
transform 1 0 3404 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1605641404
transform 1 0 4508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1605641404
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8740 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_76
timestamp 1605641404
transform 1 0 8096 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1605641404
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1605641404
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1605641404
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1605641404
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13892 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_132
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_138
timestamp 1605641404
transform 1 0 13800 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1605641404
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14904 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_149
timestamp 1605641404
transform 1 0 14812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1605641404
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1605641404
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1605641404
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1605641404
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1605641404
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1605641404
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_19
timestamp 1605641404
transform 1 0 2852 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3404 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1605641404
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1605641404
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1605641404
transform 1 0 4876 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_49
timestamp 1605641404
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5244 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1605641404
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1605641404
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6716 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1605641404
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8372 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7084 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1605641404
transform 1 0 6992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_81
timestamp 1605641404
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_71
timestamp 1605641404
transform 1 0 7636 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1605641404
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_99
timestamp 1605641404
transform 1 0 10212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1605641404
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11408 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_106
timestamp 1605641404
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_110
timestamp 1605641404
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1605641404
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1605641404
transform 1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 13064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1605641404
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp 1605641404
transform 1 0 13340 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1605641404
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1605641404
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1605641404
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15088 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1605641404
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1605641404
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15824 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 16284 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1605641404
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp 1605641404
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_169
timestamp 1605641404
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 16836 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1605641404
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1605641404
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_175
timestamp 1605641404
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1605641404
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_191
timestamp 1605641404
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_203
timestamp 1605641404
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1605641404
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1605641404
transform 1 0 20884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1605641404
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2208 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1605641404
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1605641404
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1605641404
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 1605641404
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1605641404
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1605641404
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10120 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1605641404
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1605641404
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1605641404
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_114
timestamp 1605641404
transform 1 0 11592 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13156 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1605641404
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17388 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_170
timestamp 1605641404
transform 1 0 16744 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_176
timestamp 1605641404
transform 1 0 17296 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_183
timestamp 1605641404
transform 1 0 17940 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_195
timestamp 1605641404
transform 1 0 19044 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1605641404
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1605641404
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 2944 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1605641404
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1605641404
transform 1 0 3220 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_36
timestamp 1605641404
transform 1 0 4416 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_42
timestamp 1605641404
transform 1 0 4968 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7360 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1605641404
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9568 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1605641404
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1605641404
transform 1 0 11224 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1605641404
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1605641404
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1605641404
transform 1 0 11500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1605641404
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_150
timestamp 1605641404
transform 1 0 14904 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_162
timestamp 1605641404
transform 1 0 16008 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1605641404
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1605641404
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1605641404
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1605641404
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1605641404
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_35
timestamp 1605641404
transform 1 0 4324 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4968 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp 1605641404
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_63
timestamp 1605641404
transform 1 0 6900 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1605641404
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1605641404
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1605641404
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1605641404
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12236 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 11684 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1605641404
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_118
timestamp 1605641404
transform 1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_137
timestamp 1605641404
transform 1 0 13708 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1605641404
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1605641404
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17940 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1605641404
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_182
timestamp 1605641404
transform 1 0 17848 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_189
timestamp 1605641404
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1605641404
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1605641404
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1605641404
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1605641404
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3036 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_37
timestamp 1605641404
transform 1 0 4508 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1605641404
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_82
timestamp 1605641404
transform 1 0 8648 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9752 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 9476 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_90
timestamp 1605641404
transform 1 0 9384 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1605641404
transform 1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1605641404
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_115
timestamp 1605641404
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1605641404
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1605641404
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1605641404
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1605641404
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1605641404
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1605641404
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1605641404
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1605641404
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5244 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1605641404
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1605641404
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6900 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1605641404
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1605641404
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1605641404
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_133
timestamp 1605641404
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1605641404
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1605641404
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1605641404
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1605641404
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1605641404
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1748 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1605641404
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3036 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3404 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1605641404
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_34
timestamp 1605641404
transform 1 0 4232 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5520 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1605641404
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1605641404
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1605641404
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_59
timestamp 1605641404
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8740 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_75
timestamp 1605641404
transform 1 0 8004 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_71
timestamp 1605641404
transform 1 0 7636 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1605641404
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10488 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_13_92
timestamp 1605641404
transform 1 0 9568 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_104
timestamp 1605641404
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1605641404
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_96
timestamp 1605641404
transform 1 0 9936 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1605641404
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_122
timestamp 1605641404
transform 1 0 12328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1605641404
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_134
timestamp 1605641404
transform 1 0 13432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1605641404
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1605641404
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1605641404
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1605641404
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1605641404
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1605641404
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1605641404
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1605641404
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1605641404
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1564 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4324 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1605641404
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_32
timestamp 1605641404
transform 1 0 4048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1605641404
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1605641404
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1605641404
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7452 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_67
timestamp 1605641404
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9108 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1605641404
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1605641404
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_108
timestamp 1605641404
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1605641404
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1605641404
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1605641404
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1605641404
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1605641404
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 19228 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1605641404
transform 1 0 19136 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_201
timestamp 1605641404
transform 1 0 19596 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_213
timestamp 1605641404
transform 1 0 20700 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1605641404
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 1840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2300 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1605641404
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1605641404
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_22
timestamp 1605641404
transform 1 0 3128 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1605641404
transform 1 0 4876 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6716 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5428 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1605641404
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8372 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_77
timestamp 1605641404
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1605641404
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1605641404
transform 1 0 11132 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1605641404
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_133
timestamp 1605641404
transform 1 0 13340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1605641404
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1605641404
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1605641404
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 19688 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1605641404
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1605641404
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2760 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1605641404
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 4416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1605641404
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_55
timestamp 1605641404
transform 1 0 6164 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1605641404
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1605641404
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9292 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1605641404
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1605641404
transform 1 0 10764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1605641404
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1605641404
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1605641404
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1605641404
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1605641404
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1605641404
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1605641404
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_212
timestamp 1605641404
transform 1 0 20608 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 4324 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4784 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1605641404
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1605641404
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1605641404
transform 1 0 8188 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_107
timestamp 1605641404
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_119
timestamp 1605641404
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1605641404
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_143
timestamp 1605641404
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1605641404
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1605641404
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1605641404
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1605641404
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_13
timestamp 1605641404
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_18
timestamp 1605641404
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1605641404
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1605641404
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1605641404
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1605641404
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_59
timestamp 1605641404
transform 1 0 6532 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8740 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7176 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_71
timestamp 1605641404
transform 1 0 7636 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1605641404
transform 1 0 7084 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_75
timestamp 1605641404
transform 1 0 8004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_99
timestamp 1605641404
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1605641404
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_111
timestamp 1605641404
transform 1 0 11316 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1605641404
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1605641404
transform 1 0 11132 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1605641404
transform 1 0 12236 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1605641404
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_133
timestamp 1605641404
transform 1 0 13340 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1605641404
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1605641404
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1605641404
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1605641404
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1605641404
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1605641404
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1605641404
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1605641404
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1605641404
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1605641404
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1605641404
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1605641404
transform 1 0 3864 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp 1605641404
transform 1 0 4232 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 6256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1605641404
transform 1 0 5796 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1605641404
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1605641404
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1605641404
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1605641404
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1605641404
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1605641404
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1605641404
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2300 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1605641404
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1605641404
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1605641404
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 5060 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6072 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_46
timestamp 1605641404
transform 1 0 5336 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 7636 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_70
timestamp 1605641404
transform 1 0 7544 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1605641404
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_96
timestamp 1605641404
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_101
timestamp 1605641404
transform 1 0 10396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_113
timestamp 1605641404
transform 1 0 11500 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1605641404
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1605641404
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1605641404
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1605641404
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1605641404
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1605641404
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2576 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1840 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1605641404
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1605641404
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 4784 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1605641404
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1605641404
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_43
timestamp 1605641404
transform 1 0 5060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_49
timestamp 1605641404
transform 1 0 5612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8740 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7728 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1605641404
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1605641404
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1605641404
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1605641404
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_112
timestamp 1605641404
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1605641404
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1605641404
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1605641404
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1605641404
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1605641404
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1605641404
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1605641404
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 2300 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2852 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1605641404
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1605641404
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4692 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1605641404
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1605641404
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1605641404
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5704 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_48
timestamp 1605641404
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7452 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1605641404
transform 1 0 7176 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1605641404
transform 1 0 8924 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1605641404
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_104
timestamp 1605641404
transform 1 0 10672 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1605641404
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1605641404
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_133
timestamp 1605641404
transform 1 0 13340 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1605641404
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1605641404
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1605641404
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1605641404
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1605641404
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1605641404
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1605641404
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3312 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1605641404
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_40
timestamp 1605641404
transform 1 0 4784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7728 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_65
timestamp 1605641404
transform 1 0 7084 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_71
timestamp 1605641404
transform 1 0 7636 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9752 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_88
timestamp 1605641404
transform 1 0 9200 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1605641404
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1605641404
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1605641404
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1605641404
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1605641404
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1605641404
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1605641404
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1605641404
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 1656 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1605641404
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2760 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_18
timestamp 1605641404
transform 1 0 2760 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 3496 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4232 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1605641404
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1605641404
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_30
timestamp 1605641404
transform 1 0 3864 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_50
timestamp 1605641404
transform 1 0 5704 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_45
timestamp 1605641404
transform 1 0 5244 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1605641404
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8648 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7728 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1605641404
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1605641404
transform 1 0 7636 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1605641404
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_74
timestamp 1605641404
transform 1 0 7912 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10580 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1605641404
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1605641404
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1605641404
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12236 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1605641404
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_109
timestamp 1605641404
transform 1 0 11132 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1605641404
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_137
timestamp 1605641404
transform 1 0 13708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1605641404
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1605641404
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1605641404
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1605641404
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1605641404
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1605641404
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1605641404
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1605641404
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1605641404
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1605641404
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_19
timestamp 1605641404
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3036 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1605641404
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_56
timestamp 1605641404
transform 1 0 6256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7084 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 1605641404
transform 1 0 6992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_71
timestamp 1605641404
transform 1 0 7636 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1605641404
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1605641404
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_99
timestamp 1605641404
transform 1 0 10212 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 12052 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11040 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_107
timestamp 1605641404
transform 1 0 10948 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_117
timestamp 1605641404
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_122
timestamp 1605641404
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_134
timestamp 1605641404
transform 1 0 13432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1605641404
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1605641404
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1605641404
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1605641404
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1605641404
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1605641404
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2300 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1605641404
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1605641404
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 3036 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_25
timestamp 1605641404
transform 1 0 3404 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_37
timestamp 1605641404
transform 1 0 4508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_49
timestamp 1605641404
transform 1 0 5612 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1605641404
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10396 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1605641404
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_98
timestamp 1605641404
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_107
timestamp 1605641404
transform 1 0 10948 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1605641404
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1605641404
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1605641404
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1605641404
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1605641404
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1605641404
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 1656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2944 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1605641404
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1605641404
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_26
timestamp 1605641404
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1605641404
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1605641404
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1605641404
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1605641404
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1605641404
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1605641404
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1605641404
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1605641404
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1605641404
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1605641404
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1605641404
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1605641404
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1605641404
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 2852 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1605641404
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1605641404
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1605641404
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_47
timestamp 1605641404
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1605641404
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1605641404
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1605641404
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1605641404
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1605641404
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1605641404
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1605641404
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1605641404
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1605641404
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_17
timestamp 1605641404
transform 1 0 2668 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1605641404
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1605641404
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1605641404
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1605641404
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1605641404
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1605641404
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1605641404
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2962 0 3018 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 22466 0 22522 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 22320 11432 22800 11552 6 ccff_head
port 9 nsew default input
rlabel metal3 s 22320 19048 22800 19168 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 91 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 92 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 93 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 94 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 95 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 96 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 97 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 98 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 99 nsew default input
rlabel metal3 s 22320 3816 22800 3936 6 prog_clk
port 100 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 101 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22568
<< end >>
