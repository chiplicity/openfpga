VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__3_
  CLASS BLOCK ;
  FOREIGN cbx_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 4.120 110.000 4.720 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 12.280 110.000 12.880 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 107.600 5.430 110.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END address[6]
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 107.600 16.010 110.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 107.600 27.050 110.000 ;
    END
  END bottom_grid_pin_8_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 20.440 110.000 21.040 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 107.600 38.090 110.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 29.280 110.000 29.880 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 37.440 110.000 38.040 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 46.280 110.000 46.880 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 2.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 54.440 110.000 55.040 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 107.600 49.130 110.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 63.280 110.000 63.880 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 71.440 110.000 72.040 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.400 55.040 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 80.280 110.000 80.880 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 107.600 60.170 110.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.400 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 2.400 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 107.600 71.210 110.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 107.600 82.250 110.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 107.600 93.290 110.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 88.440 110.000 89.040 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.400 86.320 ;
    END
  END chanx_right_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END enable
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 97.280 110.000 97.880 ;
    END
  END top_grid_pin_0_
  PIN top_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END top_grid_pin_10_
  PIN top_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END top_grid_pin_12_
  PIN top_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 2.400 107.400 ;
    END
  END top_grid_pin_14_
  PIN top_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END top_grid_pin_2_
  PIN top_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 107.600 104.330 110.000 ;
    END
  END top_grid_pin_4_
  PIN top_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 105.440 110.000 106.040 ;
    END
  END top_grid_pin_6_
  PIN top_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END top_grid_pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 23.055 10.640 24.655 98.160 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 41.385 10.640 42.985 98.160 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 0.070 9.560 108.030 98.160 ;
      LAYER met2 ;
        RECT 0.090 107.320 4.870 107.850 ;
        RECT 5.710 107.320 15.450 107.850 ;
        RECT 16.290 107.320 26.490 107.850 ;
        RECT 27.330 107.320 37.530 107.850 ;
        RECT 38.370 107.320 48.570 107.850 ;
        RECT 49.410 107.320 59.610 107.850 ;
        RECT 60.450 107.320 70.650 107.850 ;
        RECT 71.490 107.320 81.690 107.850 ;
        RECT 82.530 107.320 92.730 107.850 ;
        RECT 93.570 107.320 103.770 107.850 ;
        RECT 104.610 107.320 108.470 107.850 ;
        RECT 0.090 2.680 108.470 107.320 ;
        RECT 0.090 0.270 3.950 2.680 ;
        RECT 4.790 0.270 12.690 2.680 ;
        RECT 13.530 0.270 21.890 2.680 ;
        RECT 22.730 0.270 31.090 2.680 ;
        RECT 31.930 0.270 40.290 2.680 ;
        RECT 41.130 0.270 49.490 2.680 ;
        RECT 50.330 0.270 58.690 2.680 ;
        RECT 59.530 0.270 67.890 2.680 ;
        RECT 68.730 0.270 77.090 2.680 ;
        RECT 77.930 0.270 86.290 2.680 ;
        RECT 87.130 0.270 95.490 2.680 ;
        RECT 96.330 0.270 104.690 2.680 ;
        RECT 105.530 0.270 108.470 2.680 ;
      LAYER met3 ;
        RECT 0.270 107.800 108.290 107.945 ;
        RECT 2.800 106.440 108.290 107.800 ;
        RECT 2.800 106.400 107.200 106.440 ;
        RECT 0.270 105.040 107.200 106.400 ;
        RECT 0.270 102.360 108.290 105.040 ;
        RECT 2.800 100.960 108.290 102.360 ;
        RECT 0.270 98.280 108.290 100.960 ;
        RECT 0.270 96.920 107.200 98.280 ;
        RECT 2.800 96.880 107.200 96.920 ;
        RECT 2.800 95.520 108.290 96.880 ;
        RECT 0.270 92.160 108.290 95.520 ;
        RECT 2.800 90.760 108.290 92.160 ;
        RECT 0.270 89.440 108.290 90.760 ;
        RECT 0.270 88.040 107.200 89.440 ;
        RECT 0.270 86.720 108.290 88.040 ;
        RECT 2.800 85.320 108.290 86.720 ;
        RECT 0.270 81.280 108.290 85.320 ;
        RECT 2.800 79.880 107.200 81.280 ;
        RECT 0.270 76.520 108.290 79.880 ;
        RECT 2.800 75.120 108.290 76.520 ;
        RECT 0.270 72.440 108.290 75.120 ;
        RECT 0.270 71.080 107.200 72.440 ;
        RECT 2.800 71.040 107.200 71.080 ;
        RECT 2.800 69.680 108.290 71.040 ;
        RECT 0.270 65.640 108.290 69.680 ;
        RECT 2.800 64.280 108.290 65.640 ;
        RECT 2.800 64.240 107.200 64.280 ;
        RECT 0.270 62.880 107.200 64.240 ;
        RECT 0.270 60.200 108.290 62.880 ;
        RECT 2.800 58.800 108.290 60.200 ;
        RECT 0.270 55.440 108.290 58.800 ;
        RECT 2.800 54.040 107.200 55.440 ;
        RECT 0.270 50.000 108.290 54.040 ;
        RECT 2.800 48.600 108.290 50.000 ;
        RECT 0.270 47.280 108.290 48.600 ;
        RECT 0.270 45.880 107.200 47.280 ;
        RECT 0.270 44.560 108.290 45.880 ;
        RECT 2.800 43.160 108.290 44.560 ;
        RECT 0.270 39.800 108.290 43.160 ;
        RECT 2.800 38.440 108.290 39.800 ;
        RECT 2.800 38.400 107.200 38.440 ;
        RECT 0.270 37.040 107.200 38.400 ;
        RECT 0.270 34.360 108.290 37.040 ;
        RECT 2.800 32.960 108.290 34.360 ;
        RECT 0.270 30.280 108.290 32.960 ;
        RECT 0.270 28.920 107.200 30.280 ;
        RECT 2.800 28.880 107.200 28.920 ;
        RECT 2.800 27.520 108.290 28.880 ;
        RECT 0.270 23.480 108.290 27.520 ;
        RECT 2.800 22.080 108.290 23.480 ;
        RECT 0.270 21.440 108.290 22.080 ;
        RECT 0.270 20.040 107.200 21.440 ;
        RECT 0.270 18.720 108.290 20.040 ;
        RECT 2.800 17.320 108.290 18.720 ;
        RECT 0.270 13.280 108.290 17.320 ;
        RECT 2.800 11.880 107.200 13.280 ;
        RECT 0.270 7.840 108.290 11.880 ;
        RECT 2.800 6.440 108.290 7.840 ;
        RECT 0.270 5.120 108.290 6.440 ;
        RECT 0.270 3.720 107.200 5.120 ;
        RECT 0.270 3.080 108.290 3.720 ;
        RECT 2.800 1.680 108.290 3.080 ;
        RECT 0.270 0.175 108.290 1.680 ;
      LAYER met4 ;
        RECT 0.295 98.560 108.265 107.945 ;
        RECT 0.295 10.240 22.655 98.560 ;
        RECT 25.055 10.240 40.985 98.560 ;
        RECT 43.385 10.240 108.265 98.560 ;
        RECT 0.295 0.175 108.265 10.240 ;
      LAYER met5 ;
        RECT 8.860 7.700 94.180 56.900 ;
  END
END cbx_1__3_
END LIBRARY

