VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__3_
  CLASS BLOCK ;
  FOREIGN sb_1__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 112.730 BY 123.450 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 2.080 112.730 2.680 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 121.050 4.050 123.450 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 121.050 11.410 123.450 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 6.840 112.730 7.440 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 12.280 112.730 12.880 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 17.040 112.730 17.640 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 121.050 18.770 123.450 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 121.050 26.590 123.450 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 22.480 112.730 23.080 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 27.240 112.730 27.840 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 2.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 32.680 112.730 33.280 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 121.050 33.950 123.450 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 2.400 27.840 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 121.050 41.310 123.450 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 2.400 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.400 40.080 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 38.120 112.730 38.720 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 42.880 112.730 43.480 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 48.320 112.730 48.920 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.400 71.360 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 53.080 112.730 53.680 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 58.520 112.730 59.120 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 63.960 112.730 64.560 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 68.720 112.730 69.320 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 74.160 112.730 74.760 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 121.050 49.130 123.450 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 78.920 112.730 79.520 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 121.050 56.490 123.450 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 121.050 63.850 123.450 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 121.050 71.670 123.450 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 84.360 112.730 84.960 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 121.050 79.030 123.450 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.110 121.050 86.390 123.450 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 89.120 112.730 89.720 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 121.050 94.210 123.450 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 100.000 112.730 100.600 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 121.050 101.570 123.450 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 2.400 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 2.400 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 94.560 112.730 95.160 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.400 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.400 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END left_top_grid_pin_9_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 2.400 114.200 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 121.050 108.930 123.450 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 114.960 112.730 115.560 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 120.400 112.730 121.000 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 104.760 112.730 105.360 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 2.400 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 110.200 112.730 110.800 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 2.400 120.320 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 23.510 10.640 25.110 111.760 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 42.295 10.640 43.895 111.760 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 107.180 111.605 ;
      LAYER met1 ;
        RECT 0.530 0.380 110.790 121.340 ;
      LAYER met2 ;
        RECT 0.550 120.770 3.490 121.450 ;
        RECT 4.330 120.770 10.850 121.450 ;
        RECT 11.690 120.770 18.210 121.450 ;
        RECT 19.050 120.770 26.030 121.450 ;
        RECT 26.870 120.770 33.390 121.450 ;
        RECT 34.230 120.770 40.750 121.450 ;
        RECT 41.590 120.770 48.570 121.450 ;
        RECT 49.410 120.770 55.930 121.450 ;
        RECT 56.770 120.770 63.290 121.450 ;
        RECT 64.130 120.770 71.110 121.450 ;
        RECT 71.950 120.770 78.470 121.450 ;
        RECT 79.310 120.770 85.830 121.450 ;
        RECT 86.670 120.770 93.650 121.450 ;
        RECT 94.490 120.770 101.010 121.450 ;
        RECT 101.850 120.770 108.370 121.450 ;
        RECT 109.210 120.770 110.770 121.450 ;
        RECT 0.550 2.680 110.770 120.770 ;
        RECT 0.550 0.270 2.110 2.680 ;
        RECT 2.950 0.270 6.710 2.680 ;
        RECT 7.550 0.270 11.310 2.680 ;
        RECT 12.150 0.270 15.910 2.680 ;
        RECT 16.750 0.270 20.510 2.680 ;
        RECT 21.350 0.270 25.570 2.680 ;
        RECT 26.410 0.270 30.170 2.680 ;
        RECT 31.010 0.270 34.770 2.680 ;
        RECT 35.610 0.270 39.370 2.680 ;
        RECT 40.210 0.270 43.970 2.680 ;
        RECT 44.810 0.270 49.030 2.680 ;
        RECT 49.870 0.270 53.630 2.680 ;
        RECT 54.470 0.270 58.230 2.680 ;
        RECT 59.070 0.270 62.830 2.680 ;
        RECT 63.670 0.270 67.430 2.680 ;
        RECT 68.270 0.270 72.490 2.680 ;
        RECT 73.330 0.270 77.090 2.680 ;
        RECT 77.930 0.270 81.690 2.680 ;
        RECT 82.530 0.270 86.290 2.680 ;
        RECT 87.130 0.270 90.890 2.680 ;
        RECT 91.730 0.270 95.950 2.680 ;
        RECT 96.790 0.270 100.550 2.680 ;
        RECT 101.390 0.270 105.150 2.680 ;
        RECT 105.990 0.270 109.750 2.680 ;
        RECT 110.590 0.270 110.770 2.680 ;
      LAYER met3 ;
        RECT 2.800 120.000 109.930 120.400 ;
        RECT 2.800 119.320 111.050 120.000 ;
        RECT 0.270 115.960 111.050 119.320 ;
        RECT 0.270 114.600 109.930 115.960 ;
        RECT 2.800 114.560 109.930 114.600 ;
        RECT 2.800 113.200 111.050 114.560 ;
        RECT 0.270 111.200 111.050 113.200 ;
        RECT 0.270 109.800 109.930 111.200 ;
        RECT 0.270 108.480 111.050 109.800 ;
        RECT 2.800 107.080 111.050 108.480 ;
        RECT 0.270 105.760 111.050 107.080 ;
        RECT 0.270 104.360 109.930 105.760 ;
        RECT 0.270 102.360 111.050 104.360 ;
        RECT 2.800 101.000 111.050 102.360 ;
        RECT 2.800 100.960 109.930 101.000 ;
        RECT 0.270 99.600 109.930 100.960 ;
        RECT 0.270 96.240 111.050 99.600 ;
        RECT 2.800 95.560 111.050 96.240 ;
        RECT 2.800 94.840 109.930 95.560 ;
        RECT 0.270 94.160 109.930 94.840 ;
        RECT 0.270 90.120 111.050 94.160 ;
        RECT 2.800 88.720 109.930 90.120 ;
        RECT 0.270 85.360 111.050 88.720 ;
        RECT 0.270 84.000 109.930 85.360 ;
        RECT 2.800 83.960 109.930 84.000 ;
        RECT 2.800 82.600 111.050 83.960 ;
        RECT 0.270 79.920 111.050 82.600 ;
        RECT 0.270 78.520 109.930 79.920 ;
        RECT 0.270 77.880 111.050 78.520 ;
        RECT 2.800 76.480 111.050 77.880 ;
        RECT 0.270 75.160 111.050 76.480 ;
        RECT 0.270 73.760 109.930 75.160 ;
        RECT 0.270 71.760 111.050 73.760 ;
        RECT 2.800 70.360 111.050 71.760 ;
        RECT 0.270 69.720 111.050 70.360 ;
        RECT 0.270 68.320 109.930 69.720 ;
        RECT 0.270 65.640 111.050 68.320 ;
        RECT 2.800 64.960 111.050 65.640 ;
        RECT 2.800 64.240 109.930 64.960 ;
        RECT 0.270 63.560 109.930 64.240 ;
        RECT 0.270 59.520 111.050 63.560 ;
        RECT 0.270 58.840 109.930 59.520 ;
        RECT 2.800 58.120 109.930 58.840 ;
        RECT 2.800 57.440 111.050 58.120 ;
        RECT 0.270 54.080 111.050 57.440 ;
        RECT 0.270 52.720 109.930 54.080 ;
        RECT 2.800 52.680 109.930 52.720 ;
        RECT 2.800 51.320 111.050 52.680 ;
        RECT 0.270 49.320 111.050 51.320 ;
        RECT 0.270 47.920 109.930 49.320 ;
        RECT 0.270 46.600 111.050 47.920 ;
        RECT 2.800 45.200 111.050 46.600 ;
        RECT 0.270 43.880 111.050 45.200 ;
        RECT 0.270 42.480 109.930 43.880 ;
        RECT 0.270 40.480 111.050 42.480 ;
        RECT 2.800 39.120 111.050 40.480 ;
        RECT 2.800 39.080 109.930 39.120 ;
        RECT 0.270 37.720 109.930 39.080 ;
        RECT 0.270 34.360 111.050 37.720 ;
        RECT 2.800 33.680 111.050 34.360 ;
        RECT 2.800 32.960 109.930 33.680 ;
        RECT 0.270 32.280 109.930 32.960 ;
        RECT 0.270 28.240 111.050 32.280 ;
        RECT 2.800 26.840 109.930 28.240 ;
        RECT 0.270 23.480 111.050 26.840 ;
        RECT 0.270 22.120 109.930 23.480 ;
        RECT 2.800 22.080 109.930 22.120 ;
        RECT 2.800 20.720 111.050 22.080 ;
        RECT 0.270 18.040 111.050 20.720 ;
        RECT 0.270 16.640 109.930 18.040 ;
        RECT 0.270 16.000 111.050 16.640 ;
        RECT 2.800 14.600 111.050 16.000 ;
        RECT 0.270 13.280 111.050 14.600 ;
        RECT 0.270 11.880 109.930 13.280 ;
        RECT 0.270 9.880 111.050 11.880 ;
        RECT 2.800 8.480 111.050 9.880 ;
        RECT 0.270 7.840 111.050 8.480 ;
        RECT 0.270 6.975 109.930 7.840 ;
      LAYER met4 ;
        RECT 0.295 10.640 23.110 111.760 ;
        RECT 25.510 10.640 41.895 111.760 ;
        RECT 44.295 10.640 111.025 111.760 ;
  END
END sb_1__3_
END LIBRARY

