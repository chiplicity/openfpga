magic
tech sky130A
magscale 1 2
timestamp 1609016933
<< obsli1 >>
rect 1104 2015 22051 20545
<< obsm1 >>
rect 290 1156 22710 20576
<< metal2 >>
rect 294 22056 350 22856
rect 846 22056 902 22856
rect 1398 22056 1454 22856
rect 1950 22056 2006 22856
rect 2502 22056 2558 22856
rect 3054 22056 3110 22856
rect 3606 22056 3662 22856
rect 4158 22056 4214 22856
rect 4710 22056 4766 22856
rect 5262 22056 5318 22856
rect 5814 22056 5870 22856
rect 6458 22056 6514 22856
rect 7010 22056 7066 22856
rect 7562 22056 7618 22856
rect 8114 22056 8170 22856
rect 8666 22056 8722 22856
rect 9218 22056 9274 22856
rect 9770 22056 9826 22856
rect 10322 22056 10378 22856
rect 10874 22056 10930 22856
rect 11426 22056 11482 22856
rect 12070 22056 12126 22856
rect 12622 22056 12678 22856
rect 13174 22056 13230 22856
rect 13726 22056 13782 22856
rect 14278 22056 14334 22856
rect 14830 22056 14886 22856
rect 15382 22056 15438 22856
rect 15934 22056 15990 22856
rect 16486 22056 16542 22856
rect 17038 22056 17094 22856
rect 17682 22056 17738 22856
rect 18234 22056 18290 22856
rect 18786 22056 18842 22856
rect 19338 22056 19394 22856
rect 19890 22056 19946 22856
rect 20442 22056 20498 22856
rect 20994 22056 21050 22856
rect 21546 22056 21602 22856
rect 22098 22056 22154 22856
rect 22650 22056 22706 22856
<< obsm2 >>
rect 406 22000 790 22537
rect 958 22000 1342 22537
rect 1510 22000 1894 22537
rect 2062 22000 2446 22537
rect 2614 22000 2998 22537
rect 3166 22000 3550 22537
rect 3718 22000 4102 22537
rect 4270 22000 4654 22537
rect 4822 22000 5206 22537
rect 5374 22000 5758 22537
rect 5926 22000 6402 22537
rect 6570 22000 6954 22537
rect 7122 22000 7506 22537
rect 7674 22000 8058 22537
rect 8226 22000 8610 22537
rect 8778 22000 9162 22537
rect 9330 22000 9714 22537
rect 9882 22000 10266 22537
rect 10434 22000 10818 22537
rect 10986 22000 11370 22537
rect 11538 22000 12014 22537
rect 12182 22000 12566 22537
rect 12734 22000 13118 22537
rect 13286 22000 13670 22537
rect 13838 22000 14222 22537
rect 14390 22000 14774 22537
rect 14942 22000 15326 22537
rect 15494 22000 15878 22537
rect 16046 22000 16430 22537
rect 16598 22000 16982 22537
rect 17150 22000 17626 22537
rect 17794 22000 18178 22537
rect 18346 22000 18730 22537
rect 18898 22000 19282 22537
rect 19450 22000 19834 22537
rect 20002 22000 20386 22537
rect 20554 22000 20938 22537
rect 21106 22000 21490 22537
rect 21658 22000 22042 22537
rect 22210 22000 22594 22537
rect 296 23 22704 22000
<< metal3 >>
rect 22200 22440 23000 22560
rect 22200 22032 23000 22152
rect 22200 21488 23000 21608
rect 22200 21080 23000 21200
rect 22200 20672 23000 20792
rect 22200 20128 23000 20248
rect 22200 19720 23000 19840
rect 22200 19176 23000 19296
rect 22200 18768 23000 18888
rect 22200 18360 23000 18480
rect 22200 17816 23000 17936
rect 22200 17408 23000 17528
rect 0 17000 800 17120
rect 22200 17000 23000 17120
rect 22200 16456 23000 16576
rect 22200 16048 23000 16168
rect 22200 15504 23000 15624
rect 22200 15096 23000 15216
rect 22200 14688 23000 14808
rect 22200 14144 23000 14264
rect 22200 13736 23000 13856
rect 22200 13328 23000 13448
rect 22200 12784 23000 12904
rect 22200 12376 23000 12496
rect 22200 11832 23000 11952
rect 22200 11424 23000 11544
rect 22200 11016 23000 11136
rect 22200 10472 23000 10592
rect 22200 10064 23000 10184
rect 22200 9520 23000 9640
rect 22200 9112 23000 9232
rect 22200 8704 23000 8824
rect 22200 8160 23000 8280
rect 22200 7752 23000 7872
rect 22200 7344 23000 7464
rect 22200 6800 23000 6920
rect 22200 6392 23000 6512
rect 22200 5848 23000 5968
rect 0 5576 800 5696
rect 22200 5440 23000 5560
rect 22200 5032 23000 5152
rect 22200 4488 23000 4608
rect 22200 4080 23000 4200
rect 22200 3672 23000 3792
rect 22200 3128 23000 3248
rect 22200 2720 23000 2840
rect 22200 2176 23000 2296
rect 22200 1768 23000 1888
rect 22200 1360 23000 1480
rect 22200 816 23000 936
rect 22200 408 23000 528
rect 22200 0 23000 120
<< obsm3 >>
rect 800 22360 22120 22533
rect 800 22232 22200 22360
rect 800 21952 22120 22232
rect 800 21688 22200 21952
rect 800 21408 22120 21688
rect 800 21280 22200 21408
rect 800 21000 22120 21280
rect 800 20872 22200 21000
rect 800 20592 22120 20872
rect 800 20328 22200 20592
rect 800 20048 22120 20328
rect 800 19920 22200 20048
rect 800 19640 22120 19920
rect 800 19376 22200 19640
rect 800 19096 22120 19376
rect 800 18968 22200 19096
rect 800 18688 22120 18968
rect 800 18560 22200 18688
rect 800 18280 22120 18560
rect 800 18016 22200 18280
rect 800 17736 22120 18016
rect 800 17608 22200 17736
rect 800 17328 22120 17608
rect 800 17200 22200 17328
rect 880 16920 22120 17200
rect 800 16656 22200 16920
rect 800 16376 22120 16656
rect 800 16248 22200 16376
rect 800 15968 22120 16248
rect 800 15704 22200 15968
rect 800 15424 22120 15704
rect 800 15296 22200 15424
rect 800 15016 22120 15296
rect 800 14888 22200 15016
rect 800 14608 22120 14888
rect 800 14344 22200 14608
rect 800 14064 22120 14344
rect 800 13936 22200 14064
rect 800 13656 22120 13936
rect 800 13528 22200 13656
rect 800 13248 22120 13528
rect 800 12984 22200 13248
rect 800 12704 22120 12984
rect 800 12576 22200 12704
rect 800 12296 22120 12576
rect 800 12032 22200 12296
rect 800 11752 22120 12032
rect 800 11624 22200 11752
rect 800 11344 22120 11624
rect 800 11216 22200 11344
rect 800 10936 22120 11216
rect 800 10672 22200 10936
rect 800 10392 22120 10672
rect 800 10264 22200 10392
rect 800 9984 22120 10264
rect 800 9720 22200 9984
rect 800 9440 22120 9720
rect 800 9312 22200 9440
rect 800 9032 22120 9312
rect 800 8904 22200 9032
rect 800 8624 22120 8904
rect 800 8360 22200 8624
rect 800 8080 22120 8360
rect 800 7952 22200 8080
rect 800 7672 22120 7952
rect 800 7544 22200 7672
rect 800 7264 22120 7544
rect 800 7000 22200 7264
rect 800 6720 22120 7000
rect 800 6592 22200 6720
rect 800 6312 22120 6592
rect 800 6048 22200 6312
rect 800 5776 22120 6048
rect 880 5768 22120 5776
rect 880 5640 22200 5768
rect 880 5496 22120 5640
rect 800 5360 22120 5496
rect 800 5232 22200 5360
rect 800 4952 22120 5232
rect 800 4688 22200 4952
rect 800 4408 22120 4688
rect 800 4280 22200 4408
rect 800 4000 22120 4280
rect 800 3872 22200 4000
rect 800 3592 22120 3872
rect 800 3328 22200 3592
rect 800 3048 22120 3328
rect 800 2920 22200 3048
rect 800 2640 22120 2920
rect 800 2376 22200 2640
rect 800 2096 22120 2376
rect 800 1968 22200 2096
rect 800 1688 22120 1968
rect 800 1560 22200 1688
rect 800 1280 22120 1560
rect 800 1016 22200 1280
rect 800 736 22120 1016
rect 800 608 22200 736
rect 800 328 22120 608
rect 800 200 22200 328
rect 800 27 22120 200
<< metal4 >>
rect 4409 1984 4729 20576
rect 7875 1984 8195 20576
rect 11340 1984 11660 20576
rect 14805 1984 15125 20576
rect 18271 1984 18591 20576
<< obsm4 >>
rect 8275 1984 11260 20576
rect 11740 1984 14725 20576
rect 15205 1984 18191 20576
<< labels >>
rlabel metal3 s 0 5576 800 5696 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 0 17000 800 17120 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 22200 4080 23000 4200 6 chanx_right_in[0]
port 3 nsew signal input
rlabel metal3 s 22200 8704 23000 8824 6 chanx_right_in[10]
port 4 nsew signal input
rlabel metal3 s 22200 9112 23000 9232 6 chanx_right_in[11]
port 5 nsew signal input
rlabel metal3 s 22200 9520 23000 9640 6 chanx_right_in[12]
port 6 nsew signal input
rlabel metal3 s 22200 10064 23000 10184 6 chanx_right_in[13]
port 7 nsew signal input
rlabel metal3 s 22200 10472 23000 10592 6 chanx_right_in[14]
port 8 nsew signal input
rlabel metal3 s 22200 11016 23000 11136 6 chanx_right_in[15]
port 9 nsew signal input
rlabel metal3 s 22200 11424 23000 11544 6 chanx_right_in[16]
port 10 nsew signal input
rlabel metal3 s 22200 11832 23000 11952 6 chanx_right_in[17]
port 11 nsew signal input
rlabel metal3 s 22200 12376 23000 12496 6 chanx_right_in[18]
port 12 nsew signal input
rlabel metal3 s 22200 12784 23000 12904 6 chanx_right_in[19]
port 13 nsew signal input
rlabel metal3 s 22200 4488 23000 4608 6 chanx_right_in[1]
port 14 nsew signal input
rlabel metal3 s 22200 5032 23000 5152 6 chanx_right_in[2]
port 15 nsew signal input
rlabel metal3 s 22200 5440 23000 5560 6 chanx_right_in[3]
port 16 nsew signal input
rlabel metal3 s 22200 5848 23000 5968 6 chanx_right_in[4]
port 17 nsew signal input
rlabel metal3 s 22200 6392 23000 6512 6 chanx_right_in[5]
port 18 nsew signal input
rlabel metal3 s 22200 6800 23000 6920 6 chanx_right_in[6]
port 19 nsew signal input
rlabel metal3 s 22200 7344 23000 7464 6 chanx_right_in[7]
port 20 nsew signal input
rlabel metal3 s 22200 7752 23000 7872 6 chanx_right_in[8]
port 21 nsew signal input
rlabel metal3 s 22200 8160 23000 8280 6 chanx_right_in[9]
port 22 nsew signal input
rlabel metal3 s 22200 13328 23000 13448 6 chanx_right_out[0]
port 23 nsew signal output
rlabel metal3 s 22200 17816 23000 17936 6 chanx_right_out[10]
port 24 nsew signal output
rlabel metal3 s 22200 18360 23000 18480 6 chanx_right_out[11]
port 25 nsew signal output
rlabel metal3 s 22200 18768 23000 18888 6 chanx_right_out[12]
port 26 nsew signal output
rlabel metal3 s 22200 19176 23000 19296 6 chanx_right_out[13]
port 27 nsew signal output
rlabel metal3 s 22200 19720 23000 19840 6 chanx_right_out[14]
port 28 nsew signal output
rlabel metal3 s 22200 20128 23000 20248 6 chanx_right_out[15]
port 29 nsew signal output
rlabel metal3 s 22200 20672 23000 20792 6 chanx_right_out[16]
port 30 nsew signal output
rlabel metal3 s 22200 21080 23000 21200 6 chanx_right_out[17]
port 31 nsew signal output
rlabel metal3 s 22200 21488 23000 21608 6 chanx_right_out[18]
port 32 nsew signal output
rlabel metal3 s 22200 22032 23000 22152 6 chanx_right_out[19]
port 33 nsew signal output
rlabel metal3 s 22200 13736 23000 13856 6 chanx_right_out[1]
port 34 nsew signal output
rlabel metal3 s 22200 14144 23000 14264 6 chanx_right_out[2]
port 35 nsew signal output
rlabel metal3 s 22200 14688 23000 14808 6 chanx_right_out[3]
port 36 nsew signal output
rlabel metal3 s 22200 15096 23000 15216 6 chanx_right_out[4]
port 37 nsew signal output
rlabel metal3 s 22200 15504 23000 15624 6 chanx_right_out[5]
port 38 nsew signal output
rlabel metal3 s 22200 16048 23000 16168 6 chanx_right_out[6]
port 39 nsew signal output
rlabel metal3 s 22200 16456 23000 16576 6 chanx_right_out[7]
port 40 nsew signal output
rlabel metal3 s 22200 17000 23000 17120 6 chanx_right_out[8]
port 41 nsew signal output
rlabel metal3 s 22200 17408 23000 17528 6 chanx_right_out[9]
port 42 nsew signal output
rlabel metal2 s 846 22056 902 22856 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 6458 22056 6514 22856 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 7010 22056 7066 22856 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 7562 22056 7618 22856 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 8114 22056 8170 22856 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 8666 22056 8722 22856 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 9218 22056 9274 22856 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 9770 22056 9826 22856 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 10322 22056 10378 22856 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 10874 22056 10930 22856 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 11426 22056 11482 22856 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 1398 22056 1454 22856 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 1950 22056 2006 22856 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 2502 22056 2558 22856 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 3054 22056 3110 22856 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 3606 22056 3662 22856 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 4158 22056 4214 22856 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 4710 22056 4766 22856 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 5262 22056 5318 22856 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 5814 22056 5870 22856 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 12070 22056 12126 22856 6 chany_top_out[0]
port 63 nsew signal output
rlabel metal2 s 17682 22056 17738 22856 6 chany_top_out[10]
port 64 nsew signal output
rlabel metal2 s 18234 22056 18290 22856 6 chany_top_out[11]
port 65 nsew signal output
rlabel metal2 s 18786 22056 18842 22856 6 chany_top_out[12]
port 66 nsew signal output
rlabel metal2 s 19338 22056 19394 22856 6 chany_top_out[13]
port 67 nsew signal output
rlabel metal2 s 19890 22056 19946 22856 6 chany_top_out[14]
port 68 nsew signal output
rlabel metal2 s 20442 22056 20498 22856 6 chany_top_out[15]
port 69 nsew signal output
rlabel metal2 s 20994 22056 21050 22856 6 chany_top_out[16]
port 70 nsew signal output
rlabel metal2 s 21546 22056 21602 22856 6 chany_top_out[17]
port 71 nsew signal output
rlabel metal2 s 22098 22056 22154 22856 6 chany_top_out[18]
port 72 nsew signal output
rlabel metal2 s 22650 22056 22706 22856 6 chany_top_out[19]
port 73 nsew signal output
rlabel metal2 s 12622 22056 12678 22856 6 chany_top_out[1]
port 74 nsew signal output
rlabel metal2 s 13174 22056 13230 22856 6 chany_top_out[2]
port 75 nsew signal output
rlabel metal2 s 13726 22056 13782 22856 6 chany_top_out[3]
port 76 nsew signal output
rlabel metal2 s 14278 22056 14334 22856 6 chany_top_out[4]
port 77 nsew signal output
rlabel metal2 s 14830 22056 14886 22856 6 chany_top_out[5]
port 78 nsew signal output
rlabel metal2 s 15382 22056 15438 22856 6 chany_top_out[6]
port 79 nsew signal output
rlabel metal2 s 15934 22056 15990 22856 6 chany_top_out[7]
port 80 nsew signal output
rlabel metal2 s 16486 22056 16542 22856 6 chany_top_out[8]
port 81 nsew signal output
rlabel metal2 s 17038 22056 17094 22856 6 chany_top_out[9]
port 82 nsew signal output
rlabel metal3 s 22200 22440 23000 22560 6 prog_clk_0_E_in
port 83 nsew signal input
rlabel metal3 s 22200 2176 23000 2296 6 right_bottom_grid_pin_11_
port 84 nsew signal input
rlabel metal3 s 22200 2720 23000 2840 6 right_bottom_grid_pin_13_
port 85 nsew signal input
rlabel metal3 s 22200 3128 23000 3248 6 right_bottom_grid_pin_15_
port 86 nsew signal input
rlabel metal3 s 22200 3672 23000 3792 6 right_bottom_grid_pin_17_
port 87 nsew signal input
rlabel metal3 s 22200 0 23000 120 6 right_bottom_grid_pin_1_
port 88 nsew signal input
rlabel metal3 s 22200 408 23000 528 6 right_bottom_grid_pin_3_
port 89 nsew signal input
rlabel metal3 s 22200 816 23000 936 6 right_bottom_grid_pin_5_
port 90 nsew signal input
rlabel metal3 s 22200 1360 23000 1480 6 right_bottom_grid_pin_7_
port 91 nsew signal input
rlabel metal3 s 22200 1768 23000 1888 6 right_bottom_grid_pin_9_
port 92 nsew signal input
rlabel metal2 s 294 22056 350 22856 6 top_left_grid_pin_1_
port 93 nsew signal input
rlabel metal4 s 18271 1984 18591 20576 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 11340 1984 11660 20576 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 4409 1984 4729 20576 6 VPWR
port 96 nsew power bidirectional
rlabel metal4 s 14805 1984 15125 20576 6 VGND
port 97 nsew ground bidirectional
rlabel metal4 s 7875 1984 8195 20576 6 VGND
port 98 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 23000 22856
string LEFview TRUE
<< end >>
