* NGSPICE file created from cby_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt cby_2__1_ IO_ISOL_N ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ left_grid_pin_16_ left_grid_pin_17_ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_
+ left_grid_pin_21_ left_grid_pin_22_ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_
+ left_grid_pin_26_ left_grid_pin_27_ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_
+ left_grid_pin_31_ left_width_0_height_0__pin_0_ left_width_0_height_0__pin_1_lower
+ left_width_0_height_0__pin_1_upper prog_clk_0_N_out prog_clk_0_S_out prog_clk_0_W_in
+ right_grid_pin_0_ VPWR VGND
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.mux_l2_in_0_ mux_right_ipin_11.mux_l1_in_1_/X mux_right_ipin_11.mux_l1_in_0_/X
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_66_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_15.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_11.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_11.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_49_ chany_top_in[15] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_65_ chany_bottom_in[11] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_24_ sky130_fd_sc_hd__buf_4
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_11.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_11.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_48_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_64_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.mux_l2_in_3_ _32_/HI chany_top_in[14] mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_47_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_3.mux_l4_in_0_ mux_right_ipin_3.mux_l3_in_1_/X mux_right_ipin_3.mux_l3_in_0_/X
+ mux_right_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l2_in_3_ _20_/HI chany_top_in[19] mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l3_in_1_ mux_right_ipin_3.mux_l2_in_3_/X mux_right_ipin_3.mux_l2_in_2_/X
+ mux_right_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_63_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[8] mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmux_right_ipin_8.mux_l4_in_0_ mux_right_ipin_8.mux_l3_in_1_/X mux_right_ipin_8.mux_l3_in_0_/X
+ mux_right_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_46_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_17_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_8.mux_l3_in_1_ mux_right_ipin_8.mux_l2_in_3_/X mux_right_ipin_8.mux_l2_in_2_/X
+ mux_right_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[13] mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_3.mux_l3_in_0_ mux_right_ipin_3.mux_l2_in_1_/X mux_right_ipin_3.mux_l2_in_0_/X
+ mux_right_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_1_ chany_bottom_in[8] mux_right_ipin_3.mux_l1_in_2_/X
+ mux_right_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_45_ chany_top_in[11] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_3_ _27_/HI chany_top_in[17] mux_right_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_8.mux_l3_in_0_ mux_right_ipin_8.mux_l2_in_1_/X mux_right_ipin_8.mux_l2_in_0_/X
+ mux_right_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_8.mux_l1_in_2_/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.mux_l4_in_0_ mux_right_ipin_12.mux_l3_in_1_/X mux_right_ipin_12.mux_l3_in_0_/X
+ mux_right_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l1_in_2_ chany_top_in[9] chany_bottom_in[9] mux_right_ipin_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ chany_bottom_in[7] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l3_in_1_ mux_right_ipin_12.mux_l2_in_3_/X mux_right_ipin_12.mux_l2_in_2_/X
+ mux_right_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l2_in_0_ mux_right_ipin_3.mux_l1_in_1_/X mux_right_ipin_3.mux_l1_in_0_/X
+ mux_right_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[13] mux_right_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_3.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_8.mux_l2_in_0_ mux_right_ipin_8.mux_l1_in_1_/X mux_right_ipin_8.mux_l1_in_0_/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_8.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_60_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l3_in_0_ mux_right_ipin_12.mux_l2_in_1_/X mux_right_ipin_12.mux_l2_in_0_/X
+ mux_right_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_12.mux_l1_in_2_/X
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_12.mux_l1_in_2_ chany_top_in[7] chany_bottom_in[7] mux_right_ipin_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_8.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_42_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_0_ mux_right_ipin_12.mux_l1_in_1_/X mux_right_ipin_12.mux_l1_in_0_/X
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_12.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_28_ sky130_fd_sc_hd__buf_4
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_12.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_20_ sky130_fd_sc_hd__buf_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_41_ chany_top_in[7] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_12.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_40_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_6.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_4.mux_l2_in_3_ _33_/HI chany_top_in[15] mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_23_ VGND VGND VPWR VPWR _23_/HI _23_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_3.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_left_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_4.mux_l4_in_0_ mux_right_ipin_4.mux_l3_in_1_/X mux_right_ipin_4.mux_l3_in_0_/X
+ mux_right_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_9.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_9.mux_l2_in_3_ _21_/HI chany_top_in[14] mux_right_ipin_9.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l3_in_1_ mux_right_ipin_4.mux_l2_in_3_/X mux_right_ipin_4.mux_l2_in_2_/X
+ mux_right_ipin_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[9] mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_22_ VGND VGND VPWR VPWR _22_/HI _22_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_9.mux_l4_in_0_ mux_right_ipin_9.mux_l3_in_1_/X mux_right_ipin_9.mux_l3_in_0_/X
+ mux_right_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR left_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_4
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_9.mux_l3_in_1_ mux_right_ipin_9.mux_l2_in_3_/X mux_right_ipin_9.mux_l2_in_2_/X
+ mux_right_ipin_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_14.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_9.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_4.mux_l3_in_0_ mux_right_ipin_4.mux_l2_in_1_/X mux_right_ipin_4.mux_l2_in_0_/X
+ mux_right_ipin_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_11.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_21_ VGND VGND VPWR VPWR _21_/HI _21_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_4.mux_l2_in_1_ chany_bottom_in[9] mux_right_ipin_4.mux_l1_in_2_/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_15.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_31_ sky130_fd_sc_hd__buf_4
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_13.mux_l2_in_3_ _28_/HI chany_top_in[18] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_23_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_4.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.mux_l3_in_0_ mux_right_ipin_9.mux_l2_in_1_/X mux_right_ipin_9.mux_l2_in_0_/X
+ mux_right_ipin_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_9.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_13.mux_l4_in_0_ mux_right_ipin_13.mux_l3_in_1_/X mux_right_ipin_13.mux_l3_in_0_/X
+ mux_right_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_13.mux_l3_in_1_ mux_right_ipin_13.mux_l2_in_3_/X mux_right_ipin_13.mux_l2_in_2_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l2_in_0_ mux_right_ipin_4.mux_l1_in_1_/X mux_right_ipin_4.mux_l1_in_0_/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20_ VGND VGND VPWR VPWR _20_/HI _20_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_4.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_9.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_9.mux_l1_in_0_/X
+ mux_right_ipin_9.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l3_in_0_ mux_right_ipin_13.mux_l2_in_1_/X mux_right_ipin_13.mux_l2_in_0_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_16_ sky130_fd_sc_hd__buf_4
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_9.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_13.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_13.mux_l1_in_0_/X
+ mux_right_ipin_13.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_13.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_0.mux_l2_in_3_ _23_/HI chany_top_in[17] mux_right_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_59_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_5.mux_l2_in_3_ _17_/HI chany_top_in[18] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[11] mux_right_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_5.mux_l4_in_0_ mux_right_ipin_5.mux_l3_in_1_/X mux_right_ipin_5.mux_l3_in_0_/X
+ mux_right_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l3_in_1_ mux_right_ipin_5.mux_l2_in_3_/X mux_right_ipin_5.mux_l2_in_2_/X
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_58_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_5.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_11.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_27_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_19_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_5.mux_l3_in_0_ mux_right_ipin_5.mux_l2_in_1_/X mux_right_ipin_5.mux_l2_in_0_/X
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_74_ left_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR left_width_0_height_0__pin_1_upper
+ sky130_fd_sc_hd__buf_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ chany_bottom_in[3] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_5.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE left_width_0_height_0__pin_0_
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ sky130_fd_sc_hd__ebufn_4
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_14.mux_l2_in_3_ _29_/HI chany_top_in[19] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l4_in_0_ mux_right_ipin_14.mux_l3_in_1_/X mux_right_ipin_14.mux_l3_in_0_/X
+ mux_right_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_73_ chany_bottom_in[19] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_14.mux_l3_in_1_ mux_right_ipin_14.mux_l2_in_3_/X mux_right_ipin_14.mux_l2_in_2_/X
+ mux_right_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_56_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_5.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_5.mux_l1_in_0_/X
+ mux_right_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_39_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_14.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_72_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ chany_bottom_in[1] VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l3_in_0_ mux_right_ipin_14.mux_l2_in_1_/X mux_right_ipin_14.mux_l2_in_0_/X
+ mux_right_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_38_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_5.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_71_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_54_ chany_bottom_in[0] VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_37_ chany_top_in[3] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_10.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_14.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_14.mux_l1_in_0_/X
+ mux_right_ipin_14.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_14.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_30_ sky130_fd_sc_hd__buf_4
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_22_ sky130_fd_sc_hd__buf_4
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_13.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_53_ chany_top_in[19] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_8.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19_ VGND VGND VPWR VPWR _19_/HI _19_/LO sky130_fd_sc_hd__conb_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_1.mux_l2_in_3_ _24_/HI chany_top_in[14] mux_right_ipin_1.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35_ chany_top_in[1] VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_1.mux_l4_in_0_ mux_right_ipin_1.mux_l3_in_1_/X mux_right_ipin_1.mux_l3_in_0_/X
+ mux_right_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK mux_right_ipin_15.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18_ VGND VGND VPWR VPWR _18_/HI _18_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_6.mux_l2_in_3_ _18_/HI chany_top_in[19] mux_right_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_1.mux_l3_in_1_ mux_right_ipin_1.mux_l2_in_3_/X mux_right_ipin_1.mux_l2_in_2_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_left_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_1.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_1.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l4_in_0_ mux_right_ipin_6.mux_l3_in_1_/X mux_right_ipin_6.mux_l3_in_0_/X
+ mux_right_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_51_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xprog_clk_0_S_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_S_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_6.mux_l3_in_1_ mux_right_ipin_6.mux_l2_in_3_/X mux_right_ipin_6.mux_l2_in_2_/X
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
X_34_ chany_top_in[0] VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_6.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_1.mux_l3_in_0_ mux_right_ipin_1.mux_l2_in_1_/X mux_right_ipin_1.mux_l2_in_0_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_left_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_1.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_1.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_10.mux_l2_in_3_ _25_/HI chany_top_in[15] mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_6.mux_l3_in_0_ mux_right_ipin_6.mux_l2_in_1_/X mux_right_ipin_6.mux_l2_in_0_/X
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33_ VGND VGND VPWR VPWR _33_/HI _33_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_6.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_10.mux_l4_in_0_ mux_right_ipin_10.mux_l3_in_1_/X mux_right_ipin_10.mux_l3_in_0_/X
+ mux_right_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_15.mux_l2_in_3_ _30_/HI chany_top_in[16] mux_right_ipin_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_left_ipin_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_10.mux_l3_in_1_ mux_right_ipin_10.mux_l2_in_3_/X mux_right_ipin_10.mux_l2_in_2_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_25_ sky130_fd_sc_hd__buf_4
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_1.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_1.mux_l1_in_0_/X
+ mux_right_ipin_1.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_10.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_15.mux_l4_in_0_ mux_right_ipin_15.mux_l3_in_1_/X mux_right_ipin_15.mux_l3_in_0_/X
+ mux_right_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32_ VGND VGND VPWR VPWR _32_/HI _32_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_15.mux_l3_in_1_ mux_right_ipin_15.mux_l2_in_3_/X mux_right_ipin_15.mux_l2_in_2_/X
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_6.mux_l1_in_0_/X
+ mux_right_ipin_6.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_right_ipin_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ ccff_head VGND VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_10.mux_l3_in_0_ mux_right_ipin_10.mux_l2_in_1_/X mux_right_ipin_10.mux_l2_in_0_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l3_in_0_ mux_right_ipin_15.mux_l2_in_1_/X mux_right_ipin_15.mux_l2_in_0_/X
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_15.mux_l1_in_2_/X
+ mux_right_ipin_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l2_in_3_ _22_/HI chany_top_in[16] mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_15.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_10.mux_l1_in_0_/X
+ mux_right_ipin_10.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_10.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_26_ sky130_fd_sc_hd__buf_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_18_ sky130_fd_sc_hd__buf_4
Xmux_left_ipin_0.mux_l4_in_0_ mux_left_ipin_0.mux_l3_in_1_/X mux_left_ipin_0.mux_l3_in_0_/X
+ mux_left_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.mux_l3_in_1_ mux_left_ipin_0.mux_l2_in_3_/X mux_left_ipin_0.mux_l2_in_2_/X
+ mux_left_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_15.mux_l2_in_0_ mux_right_ipin_15.mux_l1_in_1_/X mux_right_ipin_15.mux_l1_in_0_/X
+ mux_right_ipin_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_10.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.mux_l3_in_0_ mux_left_ipin_0.mux_l2_in_1_/X mux_left_ipin_0.mux_l2_in_0_/X
+ mux_left_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_left_ipin_0.mux_l1_in_2_/X mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_left_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l2_in_3_ _31_/HI chany_top_in[15] mux_right_ipin_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_N_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_N_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_2.mux_l4_in_0_ mux_right_ipin_2.mux_l3_in_1_/X mux_right_ipin_2.mux_l3_in_0_/X
+ mux_right_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_7.mux_l2_in_3_ _19_/HI chany_top_in[18] mux_right_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l2_in_0_ mux_left_ipin_0.mux_l1_in_1_/X mux_left_ipin_0.mux_l1_in_0_/X
+ mux_left_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_2.mux_l3_in_1_ mux_right_ipin_2.mux_l2_in_3_/X mux_right_ipin_2.mux_l2_in_2_/X
+ mux_right_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_left_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l4_in_0_ mux_right_ipin_7.mux_l3_in_1_/X mux_right_ipin_7.mux_l3_in_0_/X
+ mux_right_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_2.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR sky130_fd_sc_hd__or2b_4
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l3_in_1_ mux_right_ipin_7.mux_l2_in_3_/X mux_right_ipin_7.mux_l2_in_2_/X
+ mux_right_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_1.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_7.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[12] mux_right_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_2.mux_l3_in_0_ mux_right_ipin_2.mux_l2_in_1_/X mux_right_ipin_2.mux_l2_in_0_/X
+ mux_right_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_left_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_2.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_13.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_29_ sky130_fd_sc_hd__buf_4
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_21_ sky130_fd_sc_hd__buf_4
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.mux_l2_in_3_ _26_/HI chany_top_in[16] mux_right_ipin_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_69_ chany_bottom_in[15] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_7.mux_l3_in_0_ mux_right_ipin_7.mux_l2_in_1_/X mux_right_ipin_7.mux_l2_in_0_/X
+ mux_right_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_7.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_7.mux_l1_in_2_/X
+ mux_right_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.mux_l4_in_0_ mux_right_ipin_11.mux_l3_in_1_/X mux_right_ipin_11.mux_l3_in_0_/X
+ mux_right_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_7.mux_l1_in_2_ chany_top_in[8] chany_bottom_in[8] mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.mux_l3_in_1_ mux_right_ipin_11.mux_l2_in_3_/X mux_right_ipin_11.mux_l2_in_2_/X
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_2.mux_l1_in_0_/X
+ mux_right_ipin_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_left_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR right_grid_pin_0_ sky130_fd_sc_hd__buf_4
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_11.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[12] mux_right_ipin_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_68_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l2_in_0_ mux_right_ipin_7.mux_l1_in_1_/X mux_right_ipin_7.mux_l1_in_0_/X
+ mux_right_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_7.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_7.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.mux_l3_in_0_ mux_right_ipin_11.mux_l2_in_1_/X mux_right_ipin_11.mux_l2_in_0_/X
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_right_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_11.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_11.mux_l1_in_2_/X
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_67_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_11.mux_l1_in_2_ chany_top_in[6] chany_bottom_in[6] mux_right_ipin_11.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_right_ipin_12.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_right_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
.ends

