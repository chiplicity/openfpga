magic
tech sky130A
magscale 1 2
timestamp 1605122828
<< locali >>
rect 4261 14807 4295 14977
rect 10517 14875 10551 15113
rect 11621 14943 11655 15045
rect 23121 14331 23155 14433
rect 3341 13719 3375 14025
rect 12909 13175 12943 13277
rect 6837 12699 6871 12801
rect 12081 10591 12115 10761
rect 12081 9979 12115 10217
rect 14105 9979 14139 10217
rect 13001 9367 13035 9673
rect 3249 8823 3283 8925
rect 12817 7735 12851 8041
rect 22845 7327 22879 7497
rect 6377 2839 6411 3077
<< viali >>
rect 5825 23817 5859 23851
rect 24777 23817 24811 23851
rect 5641 23613 5675 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 6285 23477 6319 23511
rect 24777 23273 24811 23307
rect 24593 23137 24627 23171
rect 1593 22729 1627 22763
rect 24685 22729 24719 22763
rect 25145 22729 25179 22763
rect 23949 22593 23983 22627
rect 1409 22525 1443 22559
rect 23673 22525 23707 22559
rect 24961 22525 24995 22559
rect 25513 22525 25547 22559
rect 2053 22389 2087 22423
rect 23489 22389 23523 22423
rect 1593 21641 1627 21675
rect 1409 21437 1443 21471
rect 2053 21301 2087 21335
rect 21741 21097 21775 21131
rect 2053 21029 2087 21063
rect 1777 20961 1811 20995
rect 21557 20961 21591 20995
rect 1593 20553 1627 20587
rect 21557 20553 21591 20587
rect 20821 20417 20855 20451
rect 1409 20349 1443 20383
rect 20545 20349 20579 20383
rect 2053 20213 2087 20247
rect 2329 20213 2363 20247
rect 20361 20213 20395 20247
rect 1593 20009 1627 20043
rect 24777 20009 24811 20043
rect 1409 19873 1443 19907
rect 24593 19873 24627 19907
rect 1409 19261 1443 19295
rect 1961 19261 1995 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 1593 19125 1627 19159
rect 2421 19125 2455 19159
rect 24409 19125 24443 19159
rect 24777 19125 24811 19159
rect 2697 18921 2731 18955
rect 18245 18921 18279 18955
rect 4353 18853 4387 18887
rect 1409 18785 1443 18819
rect 2513 18785 2547 18819
rect 4077 18785 4111 18819
rect 18061 18785 18095 18819
rect 23489 18785 23523 18819
rect 24593 18785 24627 18819
rect 22477 18717 22511 18751
rect 1593 18581 1627 18615
rect 1961 18581 1995 18615
rect 2421 18581 2455 18615
rect 23673 18581 23707 18615
rect 24777 18581 24811 18615
rect 1593 18377 1627 18411
rect 24777 18377 24811 18411
rect 1409 18173 1443 18207
rect 2513 18173 2547 18207
rect 22477 18173 22511 18207
rect 24593 18173 24627 18207
rect 25145 18173 25179 18207
rect 1961 18037 1995 18071
rect 2329 18037 2363 18071
rect 2697 18037 2731 18071
rect 3157 18037 3191 18071
rect 4169 18037 4203 18071
rect 18245 18037 18279 18071
rect 22661 18037 22695 18071
rect 23121 18037 23155 18071
rect 23857 18037 23891 18071
rect 24409 18037 24443 18071
rect 2881 17833 2915 17867
rect 4261 17833 4295 17867
rect 24777 17833 24811 17867
rect 1685 17765 1719 17799
rect 17417 17765 17451 17799
rect 1409 17697 1443 17731
rect 2697 17697 2731 17731
rect 4077 17697 4111 17731
rect 17141 17697 17175 17731
rect 21097 17697 21131 17731
rect 22385 17697 22419 17731
rect 23489 17697 23523 17731
rect 24593 17697 24627 17731
rect 2513 17629 2547 17663
rect 21281 17629 21315 17663
rect 2145 17493 2179 17527
rect 3341 17493 3375 17527
rect 3617 17493 3651 17527
rect 13093 17493 13127 17527
rect 22569 17493 22603 17527
rect 23673 17493 23707 17527
rect 24777 17289 24811 17323
rect 24501 17221 24535 17255
rect 2053 17153 2087 17187
rect 2145 17153 2179 17187
rect 3341 17153 3375 17187
rect 13553 17153 13587 17187
rect 21557 17153 21591 17187
rect 3157 17085 3191 17119
rect 4445 17085 4479 17119
rect 4997 17085 5031 17119
rect 13461 17085 13495 17119
rect 21373 17085 21407 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 2789 17017 2823 17051
rect 12817 17017 12851 17051
rect 13369 17017 13403 17051
rect 20085 17017 20119 17051
rect 20545 17017 20579 17051
rect 21465 17017 21499 17051
rect 22477 17017 22511 17051
rect 23949 17017 23983 17051
rect 1593 16949 1627 16983
rect 1961 16949 1995 16983
rect 4169 16949 4203 16983
rect 4629 16949 4663 16983
rect 12173 16949 12207 16983
rect 13001 16949 13035 16983
rect 17141 16949 17175 16983
rect 18797 16949 18831 16983
rect 20821 16949 20855 16983
rect 21005 16949 21039 16983
rect 22017 16949 22051 16983
rect 22569 16949 22603 16983
rect 3617 16745 3651 16779
rect 5365 16745 5399 16779
rect 13093 16745 13127 16779
rect 18337 16745 18371 16779
rect 19901 16745 19935 16779
rect 20913 16745 20947 16779
rect 23765 16745 23799 16779
rect 25513 16745 25547 16779
rect 1869 16677 1903 16711
rect 21373 16677 21407 16711
rect 22845 16677 22879 16711
rect 24317 16677 24351 16711
rect 1961 16609 1995 16643
rect 4077 16609 4111 16643
rect 4629 16609 4663 16643
rect 5181 16609 5215 16643
rect 13185 16609 13219 16643
rect 14473 16609 14507 16643
rect 14933 16609 14967 16643
rect 16957 16609 16991 16643
rect 17213 16609 17247 16643
rect 19533 16609 19567 16643
rect 19717 16609 19751 16643
rect 21281 16609 21315 16643
rect 22293 16609 22327 16643
rect 22937 16609 22971 16643
rect 24041 16609 24075 16643
rect 25329 16609 25363 16643
rect 2053 16541 2087 16575
rect 13369 16541 13403 16575
rect 21465 16541 21499 16575
rect 23029 16541 23063 16575
rect 2513 16473 2547 16507
rect 2881 16473 2915 16507
rect 3249 16473 3283 16507
rect 4261 16473 4295 16507
rect 1501 16405 1535 16439
rect 5089 16405 5123 16439
rect 12081 16405 12115 16439
rect 12541 16405 12575 16439
rect 12725 16405 12759 16439
rect 14105 16405 14139 16439
rect 20361 16405 20395 16439
rect 20637 16405 20671 16439
rect 22017 16405 22051 16439
rect 22477 16405 22511 16439
rect 2513 16201 2547 16235
rect 5733 16201 5767 16235
rect 6101 16201 6135 16235
rect 17049 16201 17083 16235
rect 20085 16201 20119 16235
rect 22661 16201 22695 16235
rect 25421 16201 25455 16235
rect 2973 16133 3007 16167
rect 1961 16065 1995 16099
rect 2145 16065 2179 16099
rect 3617 16065 3651 16099
rect 4813 16065 4847 16099
rect 13001 16065 13035 16099
rect 14565 16065 14599 16099
rect 20637 16065 20671 16099
rect 22201 16065 22235 16099
rect 24133 16065 24167 16099
rect 24225 16065 24259 16099
rect 24685 16065 24719 16099
rect 3433 15997 3467 16031
rect 4169 15997 4203 16031
rect 4629 15997 4663 16031
rect 12817 15997 12851 16031
rect 14473 15997 14507 16031
rect 20453 15997 20487 16031
rect 21189 15997 21223 16031
rect 22017 15997 22051 16031
rect 23121 15997 23155 16031
rect 25237 15997 25271 16031
rect 1869 15929 1903 15963
rect 14381 15929 14415 15963
rect 15577 15929 15611 15963
rect 19717 15929 19751 15963
rect 21557 15929 21591 15963
rect 22109 15929 22143 15963
rect 23489 15929 23523 15963
rect 24041 15929 24075 15963
rect 1501 15861 1535 15895
rect 3065 15861 3099 15895
rect 3525 15861 3559 15895
rect 4537 15861 4571 15895
rect 5457 15861 5491 15895
rect 9413 15861 9447 15895
rect 11805 15861 11839 15895
rect 12265 15861 12299 15895
rect 12449 15861 12483 15895
rect 12909 15861 12943 15895
rect 13461 15861 13495 15895
rect 13921 15861 13955 15895
rect 14013 15861 14047 15895
rect 15393 15861 15427 15895
rect 16589 15861 16623 15895
rect 17417 15861 17451 15895
rect 18061 15861 18095 15895
rect 18613 15861 18647 15895
rect 19073 15861 19107 15895
rect 20545 15861 20579 15895
rect 21649 15861 21683 15895
rect 23673 15861 23707 15895
rect 25053 15861 25087 15895
rect 25789 15861 25823 15895
rect 2789 15657 2823 15691
rect 3801 15657 3835 15691
rect 6377 15657 6411 15691
rect 6745 15657 6779 15691
rect 7113 15657 7147 15691
rect 14197 15657 14231 15691
rect 18797 15657 18831 15691
rect 19257 15657 19291 15691
rect 23121 15657 23155 15691
rect 23673 15657 23707 15691
rect 2053 15589 2087 15623
rect 5917 15589 5951 15623
rect 11437 15589 11471 15623
rect 13737 15589 13771 15623
rect 18061 15589 18095 15623
rect 22109 15589 22143 15623
rect 22753 15589 22787 15623
rect 24685 15589 24719 15623
rect 25145 15589 25179 15623
rect 2145 15521 2179 15555
rect 4445 15521 4479 15555
rect 5641 15521 5675 15555
rect 6929 15521 6963 15555
rect 11796 15521 11830 15555
rect 15669 15521 15703 15555
rect 19625 15521 19659 15555
rect 24409 15521 24443 15555
rect 24869 15521 24903 15555
rect 2237 15453 2271 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 10517 15453 10551 15487
rect 11529 15453 11563 15487
rect 15025 15453 15059 15487
rect 15761 15453 15795 15487
rect 15945 15453 15979 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 19717 15453 19751 15487
rect 19901 15453 19935 15487
rect 22201 15453 22235 15487
rect 22385 15453 22419 15487
rect 23765 15453 23799 15487
rect 23857 15453 23891 15487
rect 1685 15385 1719 15419
rect 3433 15385 3467 15419
rect 5549 15385 5583 15419
rect 13277 15385 13311 15419
rect 17693 15385 17727 15419
rect 20637 15385 20671 15419
rect 3065 15317 3099 15351
rect 4077 15317 4111 15351
rect 5089 15317 5123 15351
rect 7573 15317 7607 15351
rect 11069 15317 11103 15351
rect 12909 15317 12943 15351
rect 13645 15317 13679 15351
rect 14657 15317 14691 15351
rect 15301 15317 15335 15351
rect 16405 15317 16439 15351
rect 16773 15317 16807 15351
rect 17141 15317 17175 15351
rect 19073 15317 19107 15351
rect 20361 15317 20395 15351
rect 21189 15317 21223 15351
rect 21465 15317 21499 15351
rect 21741 15317 21775 15351
rect 23305 15317 23339 15351
rect 7941 15113 7975 15147
rect 8309 15113 8343 15147
rect 10517 15113 10551 15147
rect 10609 15113 10643 15147
rect 10793 15113 10827 15147
rect 11805 15113 11839 15147
rect 14657 15113 14691 15147
rect 17785 15113 17819 15147
rect 21281 15113 21315 15147
rect 22201 15113 22235 15147
rect 23029 15113 23063 15147
rect 2881 15045 2915 15079
rect 1869 14977 1903 15011
rect 2053 14977 2087 15011
rect 3617 14977 3651 15011
rect 4261 14977 4295 15011
rect 5089 14977 5123 15011
rect 7021 14977 7055 15011
rect 1777 14909 1811 14943
rect 3433 14909 3467 14943
rect 3341 14841 3375 14875
rect 4997 14909 5031 14943
rect 5733 14909 5767 14943
rect 6653 14909 6687 14943
rect 6837 14909 6871 14943
rect 8125 14909 8159 14943
rect 8677 14909 8711 14943
rect 10333 14909 10367 14943
rect 11621 15045 11655 15079
rect 14197 15045 14231 15079
rect 18337 15045 18371 15079
rect 11345 14977 11379 15011
rect 12173 14977 12207 15011
rect 15209 14977 15243 15011
rect 16773 14977 16807 15011
rect 18889 14977 18923 15011
rect 22569 14977 22603 15011
rect 24225 14977 24259 15011
rect 24685 14977 24719 15011
rect 25053 14977 25087 15011
rect 25421 14977 25455 15011
rect 11161 14909 11195 14943
rect 11621 14909 11655 14943
rect 12449 14909 12483 14943
rect 12716 14909 12750 14943
rect 16129 14909 16163 14943
rect 16589 14909 16623 14943
rect 18705 14909 18739 14943
rect 19901 14909 19935 14943
rect 22293 14909 22327 14943
rect 24133 14909 24167 14943
rect 25237 14909 25271 14943
rect 25973 14909 26007 14943
rect 6101 14841 6135 14875
rect 10517 14841 10551 14875
rect 11253 14841 11287 14875
rect 15117 14841 15151 14875
rect 16681 14841 16715 14875
rect 20146 14841 20180 14875
rect 21741 14841 21775 14875
rect 24041 14841 24075 14875
rect 1409 14773 1443 14807
rect 2421 14773 2455 14807
rect 2973 14773 3007 14807
rect 3985 14773 4019 14807
rect 4261 14773 4295 14807
rect 4353 14773 4387 14807
rect 4537 14773 4571 14807
rect 4905 14773 4939 14807
rect 7665 14773 7699 14807
rect 9229 14773 9263 14807
rect 13829 14773 13863 14807
rect 14565 14773 14599 14807
rect 15025 14773 15059 14807
rect 15669 14773 15703 14807
rect 16221 14773 16255 14807
rect 17417 14773 17451 14807
rect 18797 14773 18831 14807
rect 19441 14773 19475 14807
rect 19809 14773 19843 14807
rect 23489 14773 23523 14807
rect 23673 14773 23707 14807
rect 2421 14569 2455 14603
rect 2881 14569 2915 14603
rect 5457 14569 5491 14603
rect 7849 14569 7883 14603
rect 8217 14569 8251 14603
rect 11713 14569 11747 14603
rect 14749 14569 14783 14603
rect 17969 14569 18003 14603
rect 20637 14569 20671 14603
rect 22845 14569 22879 14603
rect 23305 14569 23339 14603
rect 4905 14501 4939 14535
rect 5825 14501 5859 14535
rect 6561 14501 6595 14535
rect 13246 14501 13280 14535
rect 21434 14501 21468 14535
rect 2789 14433 2823 14467
rect 4813 14433 4847 14467
rect 6469 14433 6503 14467
rect 7665 14433 7699 14467
rect 10600 14433 10634 14467
rect 15669 14433 15703 14467
rect 17233 14433 17267 14467
rect 18880 14433 18914 14467
rect 23121 14433 23155 14467
rect 23653 14433 23687 14467
rect 1409 14365 1443 14399
rect 3065 14365 3099 14399
rect 5089 14365 5123 14399
rect 6653 14365 6687 14399
rect 10333 14365 10367 14399
rect 13001 14365 13035 14399
rect 15761 14365 15795 14399
rect 15945 14365 15979 14399
rect 17325 14365 17359 14399
rect 17417 14365 17451 14399
rect 18613 14365 18647 14399
rect 21189 14365 21223 14399
rect 23397 14365 23431 14399
rect 4445 14297 4479 14331
rect 12817 14297 12851 14331
rect 15025 14297 15059 14331
rect 18337 14297 18371 14331
rect 22569 14297 22603 14331
rect 23121 14297 23155 14331
rect 1961 14229 1995 14263
rect 2237 14229 2271 14263
rect 3525 14229 3559 14263
rect 3801 14229 3835 14263
rect 4261 14229 4295 14263
rect 6101 14229 6135 14263
rect 7297 14229 7331 14263
rect 8585 14229 8619 14263
rect 8953 14229 8987 14263
rect 9413 14229 9447 14263
rect 10241 14229 10275 14263
rect 11989 14229 12023 14263
rect 12541 14229 12575 14263
rect 14381 14229 14415 14263
rect 15301 14229 15335 14263
rect 16313 14229 16347 14263
rect 16681 14229 16715 14263
rect 16865 14229 16899 14263
rect 19993 14229 20027 14263
rect 20269 14229 20303 14263
rect 24777 14229 24811 14263
rect 25053 14229 25087 14263
rect 1777 14025 1811 14059
rect 3341 14025 3375 14059
rect 3617 14025 3651 14059
rect 5825 14025 5859 14059
rect 7205 14025 7239 14059
rect 8953 14025 8987 14059
rect 11805 14025 11839 14059
rect 12449 14025 12483 14059
rect 13461 14025 13495 14059
rect 15025 14025 15059 14059
rect 15485 14025 15519 14059
rect 21373 14025 21407 14059
rect 21833 14025 21867 14059
rect 23397 14025 23431 14059
rect 3249 13957 3283 13991
rect 1869 13821 1903 13855
rect 2114 13753 2148 13787
rect 19441 13957 19475 13991
rect 24409 13957 24443 13991
rect 3985 13889 4019 13923
rect 7113 13889 7147 13923
rect 7757 13889 7791 13923
rect 9413 13889 9447 13923
rect 13001 13889 13035 13923
rect 13921 13889 13955 13923
rect 14565 13889 14599 13923
rect 16037 13889 16071 13923
rect 16221 13889 16255 13923
rect 19809 13889 19843 13923
rect 20821 13889 20855 13923
rect 21741 13889 21775 13923
rect 22477 13889 22511 13923
rect 25053 13889 25087 13923
rect 25421 13889 25455 13923
rect 4077 13821 4111 13855
rect 4333 13821 4367 13855
rect 6193 13821 6227 13855
rect 6561 13821 6595 13855
rect 7665 13821 7699 13855
rect 8217 13821 8251 13855
rect 8585 13821 8619 13855
rect 9505 13821 9539 13855
rect 9761 13821 9795 13855
rect 11161 13821 11195 13855
rect 12909 13821 12943 13855
rect 16865 13821 16899 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 22293 13821 22327 13855
rect 22845 13821 22879 13855
rect 7573 13753 7607 13787
rect 14381 13753 14415 13787
rect 18306 13753 18340 13787
rect 20177 13753 20211 13787
rect 20637 13753 20671 13787
rect 24317 13753 24351 13787
rect 3341 13685 3375 13719
rect 5457 13685 5491 13719
rect 10885 13685 10919 13719
rect 12265 13685 12299 13719
rect 12817 13685 12851 13719
rect 14013 13685 14047 13719
rect 14473 13685 14507 13719
rect 15577 13685 15611 13719
rect 15945 13685 15979 13719
rect 17877 13685 17911 13719
rect 20269 13685 20303 13719
rect 20729 13685 20763 13719
rect 22201 13685 22235 13719
rect 23857 13685 23891 13719
rect 24777 13685 24811 13719
rect 24869 13685 24903 13719
rect 1685 13481 1719 13515
rect 3433 13481 3467 13515
rect 3893 13481 3927 13515
rect 4537 13481 4571 13515
rect 6285 13481 6319 13515
rect 8769 13481 8803 13515
rect 9045 13481 9079 13515
rect 12081 13481 12115 13515
rect 13553 13481 13587 13515
rect 13645 13481 13679 13515
rect 18705 13481 18739 13515
rect 19441 13481 19475 13515
rect 21373 13481 21407 13515
rect 21833 13481 21867 13515
rect 22477 13481 22511 13515
rect 25513 13481 25547 13515
rect 2044 13413 2078 13447
rect 7297 13413 7331 13447
rect 7634 13413 7668 13447
rect 12449 13413 12483 13447
rect 14657 13413 14691 13447
rect 19349 13413 19383 13447
rect 23388 13413 23422 13447
rect 1777 13345 1811 13379
rect 4905 13345 4939 13379
rect 5172 13345 5206 13379
rect 7389 13345 7423 13379
rect 10241 13345 10275 13379
rect 12541 13345 12575 13379
rect 14013 13345 14047 13379
rect 14105 13345 14139 13379
rect 15301 13345 15335 13379
rect 17029 13345 17063 13379
rect 21741 13345 21775 13379
rect 25329 13345 25363 13379
rect 9505 13277 9539 13311
rect 10333 13277 10367 13311
rect 10425 13277 10459 13311
rect 12725 13277 12759 13311
rect 12909 13277 12943 13311
rect 13185 13277 13219 13311
rect 14289 13277 14323 13311
rect 15485 13277 15519 13311
rect 16037 13277 16071 13311
rect 16773 13277 16807 13311
rect 19625 13277 19659 13311
rect 21925 13277 21959 13311
rect 23121 13277 23155 13311
rect 11989 13209 12023 13243
rect 20729 13209 20763 13243
rect 22753 13209 22787 13243
rect 3157 13141 3191 13175
rect 6561 13141 6595 13175
rect 9873 13141 9907 13175
rect 10885 13141 10919 13175
rect 11253 13141 11287 13175
rect 12909 13141 12943 13175
rect 15117 13141 15151 13175
rect 16405 13141 16439 13175
rect 18153 13141 18187 13175
rect 18981 13141 19015 13175
rect 20269 13141 20303 13175
rect 21281 13141 21315 13175
rect 24501 13141 24535 13175
rect 24777 13141 24811 13175
rect 25145 13141 25179 13175
rect 1869 12937 1903 12971
rect 3617 12937 3651 12971
rect 4721 12937 4755 12971
rect 7205 12937 7239 12971
rect 8769 12937 8803 12971
rect 9965 12937 9999 12971
rect 12633 12937 12667 12971
rect 15945 12937 15979 12971
rect 17785 12937 17819 12971
rect 20637 12937 20671 12971
rect 21097 12937 21131 12971
rect 21465 12937 21499 12971
rect 23121 12937 23155 12971
rect 25329 12937 25363 12971
rect 1777 12869 1811 12903
rect 19625 12869 19659 12903
rect 2421 12801 2455 12835
rect 4077 12801 4111 12835
rect 4169 12801 4203 12835
rect 5733 12801 5767 12835
rect 6193 12801 6227 12835
rect 6837 12801 6871 12835
rect 7757 12801 7791 12835
rect 8217 12801 8251 12835
rect 12909 12801 12943 12835
rect 16313 12801 16347 12835
rect 16957 12801 16991 12835
rect 18613 12801 18647 12835
rect 20177 12801 20211 12835
rect 22661 12801 22695 12835
rect 24593 12801 24627 12835
rect 25605 12801 25639 12835
rect 2973 12733 3007 12767
rect 3525 12733 3559 12767
rect 6561 12733 6595 12767
rect 7665 12733 7699 12767
rect 8861 12733 8895 12767
rect 10149 12733 10183 12767
rect 13921 12733 13955 12767
rect 14188 12733 14222 12767
rect 17509 12733 17543 12767
rect 18429 12733 18463 12767
rect 21925 12733 21959 12767
rect 22477 12733 22511 12767
rect 23489 12733 23523 12767
rect 24501 12733 24535 12767
rect 5089 12665 5123 12699
rect 5549 12665 5583 12699
rect 6837 12665 6871 12699
rect 7573 12665 7607 12699
rect 9137 12665 9171 12699
rect 10416 12665 10450 12699
rect 18521 12665 18555 12699
rect 19165 12665 19199 12699
rect 19993 12665 20027 12699
rect 24409 12665 24443 12699
rect 2237 12597 2271 12631
rect 2329 12597 2363 12631
rect 3985 12597 4019 12631
rect 5181 12597 5215 12631
rect 5641 12597 5675 12631
rect 7021 12597 7055 12631
rect 11529 12597 11563 12631
rect 12081 12597 12115 12631
rect 13737 12597 13771 12631
rect 15301 12597 15335 12631
rect 16405 12597 16439 12631
rect 16773 12597 16807 12631
rect 16865 12597 16899 12631
rect 18061 12597 18095 12631
rect 19533 12597 19567 12631
rect 20085 12597 20119 12631
rect 22017 12597 22051 12631
rect 22385 12597 22419 12631
rect 23857 12597 23891 12631
rect 24041 12597 24075 12631
rect 1593 12393 1627 12427
rect 2145 12393 2179 12427
rect 6469 12393 6503 12427
rect 8401 12393 8435 12427
rect 8953 12393 8987 12427
rect 9689 12393 9723 12427
rect 11713 12393 11747 12427
rect 15117 12393 15151 12427
rect 15577 12393 15611 12427
rect 15853 12393 15887 12427
rect 16497 12393 16531 12427
rect 18889 12393 18923 12427
rect 20085 12393 20119 12427
rect 21649 12393 21683 12427
rect 22109 12393 22143 12427
rect 23305 12393 23339 12427
rect 23673 12393 23707 12427
rect 2789 12325 2823 12359
rect 11621 12325 11655 12359
rect 17040 12325 17074 12359
rect 20361 12325 20395 12359
rect 2237 12257 2271 12291
rect 4077 12257 4111 12291
rect 4344 12257 4378 12291
rect 6101 12257 6135 12291
rect 7021 12257 7055 12291
rect 7288 12257 7322 12291
rect 10057 12257 10091 12291
rect 12909 12257 12943 12291
rect 13176 12257 13210 12291
rect 15669 12257 15703 12291
rect 19349 12257 19383 12291
rect 20729 12257 20763 12291
rect 20913 12257 20947 12291
rect 22661 12257 22695 12291
rect 23857 12257 23891 12291
rect 24124 12257 24158 12291
rect 2329 12189 2363 12223
rect 6929 12189 6963 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 10793 12189 10827 12223
rect 11161 12189 11195 12223
rect 11897 12189 11931 12223
rect 16773 12189 16807 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 21097 12189 21131 12223
rect 22753 12189 22787 12223
rect 22937 12189 22971 12223
rect 1777 12121 1811 12155
rect 3801 12121 3835 12155
rect 18981 12121 19015 12155
rect 3525 12053 3559 12087
rect 5457 12053 5491 12087
rect 5733 12053 5767 12087
rect 9505 12053 9539 12087
rect 11253 12053 11287 12087
rect 12541 12053 12575 12087
rect 14289 12053 14323 12087
rect 14657 12053 14691 12087
rect 18153 12053 18187 12087
rect 18429 12053 18463 12087
rect 20545 12053 20579 12087
rect 22293 12053 22327 12087
rect 25237 12053 25271 12087
rect 1777 11849 1811 11883
rect 3433 11849 3467 11883
rect 7849 11849 7883 11883
rect 9321 11849 9355 11883
rect 9965 11849 9999 11883
rect 10241 11849 10275 11883
rect 11345 11849 11379 11883
rect 11713 11849 11747 11883
rect 12265 11849 12299 11883
rect 13461 11849 13495 11883
rect 13921 11849 13955 11883
rect 14749 11849 14783 11883
rect 16313 11849 16347 11883
rect 16773 11849 16807 11883
rect 17141 11849 17175 11883
rect 17785 11849 17819 11883
rect 18429 11849 18463 11883
rect 20177 11849 20211 11883
rect 22477 11849 22511 11883
rect 4445 11781 4479 11815
rect 6009 11781 6043 11815
rect 7757 11781 7791 11815
rect 12449 11781 12483 11815
rect 19901 11781 19935 11815
rect 25329 11781 25363 11815
rect 2237 11713 2271 11747
rect 2329 11713 2363 11747
rect 3985 11713 4019 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 6837 11713 6871 11747
rect 8401 11713 8435 11747
rect 10701 11713 10735 11747
rect 10885 11713 10919 11747
rect 13001 11713 13035 11747
rect 18521 11713 18555 11747
rect 23949 11713 23983 11747
rect 3341 11645 3375 11679
rect 3801 11645 3835 11679
rect 4905 11645 4939 11679
rect 7389 11645 7423 11679
rect 8309 11645 8343 11679
rect 9597 11645 9631 11679
rect 12817 11645 12851 11679
rect 14933 11645 14967 11679
rect 17325 11645 17359 11679
rect 18777 11645 18811 11679
rect 20729 11645 20763 11679
rect 24216 11645 24250 11679
rect 6653 11577 6687 11611
rect 8217 11577 8251 11611
rect 8953 11577 8987 11611
rect 15200 11577 15234 11611
rect 20974 11577 21008 11611
rect 23489 11577 23523 11611
rect 1685 11509 1719 11543
rect 2145 11509 2179 11543
rect 2881 11509 2915 11543
rect 3893 11509 3927 11543
rect 4997 11509 5031 11543
rect 5365 11509 5399 11543
rect 9413 11509 9447 11543
rect 10609 11509 10643 11543
rect 12909 11509 12943 11543
rect 14197 11509 14231 11543
rect 20545 11509 20579 11543
rect 22109 11509 22143 11543
rect 22845 11509 22879 11543
rect 25697 11509 25731 11543
rect 25973 11509 26007 11543
rect 1777 11305 1811 11339
rect 2237 11305 2271 11339
rect 3525 11305 3559 11339
rect 4629 11305 4663 11339
rect 6193 11305 6227 11339
rect 8125 11305 8159 11339
rect 9689 11305 9723 11339
rect 12081 11305 12115 11339
rect 13277 11305 13311 11339
rect 13461 11305 13495 11339
rect 15025 11305 15059 11339
rect 16773 11305 16807 11339
rect 17233 11305 17267 11339
rect 18061 11305 18095 11339
rect 18337 11305 18371 11339
rect 19257 11305 19291 11339
rect 19625 11305 19659 11339
rect 21097 11305 21131 11339
rect 22845 11305 22879 11339
rect 23857 11305 23891 11339
rect 23949 11305 23983 11339
rect 24501 11305 24535 11339
rect 25237 11305 25271 11339
rect 1593 11237 1627 11271
rect 2789 11237 2823 11271
rect 5089 11237 5123 11271
rect 6561 11237 6595 11271
rect 7297 11237 7331 11271
rect 9505 11237 9539 11271
rect 12541 11237 12575 11271
rect 16313 11237 16347 11271
rect 20637 11237 20671 11271
rect 23397 11237 23431 11271
rect 24961 11237 24995 11271
rect 25697 11237 25731 11271
rect 2145 11169 2179 11203
rect 3893 11169 3927 11203
rect 4997 11169 5031 11203
rect 10708 11169 10742 11203
rect 10968 11169 11002 11203
rect 13829 11169 13863 11203
rect 15669 11169 15703 11203
rect 17141 11169 17175 11203
rect 18521 11169 18555 11203
rect 19073 11169 19107 11203
rect 19717 11169 19751 11203
rect 22201 11169 22235 11203
rect 22293 11169 22327 11203
rect 25053 11169 25087 11203
rect 2329 11101 2363 11135
rect 5181 11101 5215 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 12909 11101 12943 11135
rect 13921 11101 13955 11135
rect 14013 11101 14047 11135
rect 14473 11101 14507 11135
rect 17325 11101 17359 11135
rect 19809 11101 19843 11135
rect 21741 11101 21775 11135
rect 22477 11101 22511 11135
rect 24133 11101 24167 11135
rect 3709 11033 3743 11067
rect 4537 11033 4571 11067
rect 5641 11033 5675 11067
rect 6101 11033 6135 11067
rect 7757 11033 7791 11067
rect 10241 11033 10275 11067
rect 15853 11033 15887 11067
rect 21833 11033 21867 11067
rect 23489 11033 23523 11067
rect 7665 10965 7699 10999
rect 9045 10965 9079 10999
rect 15577 10965 15611 10999
rect 16681 10965 16715 10999
rect 1777 10761 1811 10795
rect 4077 10761 4111 10795
rect 4445 10761 4479 10795
rect 5917 10761 5951 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 9229 10761 9263 10795
rect 10057 10761 10091 10795
rect 10333 10761 10367 10795
rect 12081 10761 12115 10795
rect 12173 10761 12207 10795
rect 14841 10761 14875 10795
rect 15301 10761 15335 10795
rect 16405 10761 16439 10795
rect 16773 10761 16807 10795
rect 19257 10761 19291 10795
rect 21097 10761 21131 10795
rect 23489 10761 23523 10795
rect 3249 10693 3283 10727
rect 6653 10693 6687 10727
rect 1869 10625 1903 10659
rect 4537 10625 4571 10659
rect 9689 10625 9723 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 14289 10625 14323 10659
rect 15117 10625 15151 10659
rect 15853 10625 15887 10659
rect 17877 10625 17911 10659
rect 18705 10625 18739 10659
rect 22569 10625 22603 10659
rect 4804 10557 4838 10591
rect 6837 10557 6871 10591
rect 9045 10557 9079 10591
rect 10885 10557 10919 10591
rect 12081 10557 12115 10591
rect 12633 10557 12667 10591
rect 14105 10557 14139 10591
rect 15669 10557 15703 10591
rect 16865 10557 16899 10591
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 19717 10557 19751 10591
rect 21557 10557 21591 10591
rect 23949 10557 23983 10591
rect 25973 10557 26007 10591
rect 2136 10489 2170 10523
rect 3525 10489 3559 10523
rect 7082 10489 7116 10523
rect 19625 10489 19659 10523
rect 19984 10489 20018 10523
rect 22385 10489 22419 10523
rect 22477 10489 22511 10523
rect 24216 10489 24250 10523
rect 6285 10421 6319 10455
rect 8217 10421 8251 10455
rect 10517 10421 10551 10455
rect 11621 10421 11655 10455
rect 12817 10421 12851 10455
rect 13461 10421 13495 10455
rect 13737 10421 13771 10455
rect 14197 10421 14231 10455
rect 15761 10421 15795 10455
rect 17049 10421 17083 10455
rect 17509 10421 17543 10455
rect 18061 10421 18095 10455
rect 21833 10421 21867 10455
rect 22017 10421 22051 10455
rect 23029 10421 23063 10455
rect 25329 10421 25363 10455
rect 25605 10421 25639 10455
rect 3065 10217 3099 10251
rect 4629 10217 4663 10251
rect 6285 10217 6319 10251
rect 6837 10217 6871 10251
rect 7113 10217 7147 10251
rect 9045 10217 9079 10251
rect 10517 10217 10551 10251
rect 12081 10217 12115 10251
rect 3709 10149 3743 10183
rect 5172 10149 5206 10183
rect 1685 10081 1719 10115
rect 1952 10081 1986 10115
rect 3433 10081 3467 10115
rect 4905 10081 4939 10115
rect 7297 10081 7331 10115
rect 7656 10081 7690 10115
rect 10609 10081 10643 10115
rect 10876 10081 10910 10115
rect 7389 10013 7423 10047
rect 14105 10217 14139 10251
rect 14289 10217 14323 10251
rect 14749 10217 14783 10251
rect 15945 10217 15979 10251
rect 18153 10217 18187 10251
rect 18797 10217 18831 10251
rect 19717 10217 19751 10251
rect 20729 10217 20763 10251
rect 22293 10217 22327 10251
rect 23213 10217 23247 10251
rect 23949 10217 23983 10251
rect 24225 10217 24259 10251
rect 24869 10217 24903 10251
rect 25789 10217 25823 10251
rect 13185 10081 13219 10115
rect 13277 10013 13311 10047
rect 13369 10013 13403 10047
rect 16672 10149 16706 10183
rect 19073 10149 19107 10183
rect 15301 10081 15335 10115
rect 16405 10081 16439 10115
rect 19625 10081 19659 10115
rect 21649 10081 21683 10115
rect 22661 10081 22695 10115
rect 24777 10081 24811 10115
rect 15117 10013 15151 10047
rect 19809 10013 19843 10047
rect 21741 10013 21775 10047
rect 21925 10013 21959 10047
rect 23305 10013 23339 10047
rect 23397 10013 23431 10047
rect 24961 10013 24995 10047
rect 8769 9945 8803 9979
rect 12081 9945 12115 9979
rect 12817 9945 12851 9979
rect 14105 9945 14139 9979
rect 21189 9945 21223 9979
rect 9413 9877 9447 9911
rect 9965 9877 9999 9911
rect 11989 9877 12023 9911
rect 12265 9877 12299 9911
rect 12633 9877 12667 9911
rect 13921 9877 13955 9911
rect 15485 9877 15519 9911
rect 16221 9877 16255 9911
rect 17785 9877 17819 9911
rect 19257 9877 19291 9911
rect 20269 9877 20303 9911
rect 21281 9877 21315 9911
rect 22845 9877 22879 9911
rect 24409 9877 24443 9911
rect 25513 9877 25547 9911
rect 5733 9673 5767 9707
rect 13001 9673 13035 9707
rect 16957 9673 16991 9707
rect 17325 9673 17359 9707
rect 19809 9673 19843 9707
rect 26157 9673 26191 9707
rect 1593 9605 1627 9639
rect 4721 9605 4755 9639
rect 6653 9605 6687 9639
rect 10241 9605 10275 9639
rect 10609 9605 10643 9639
rect 2145 9537 2179 9571
rect 3801 9537 3835 9571
rect 4629 9537 4663 9571
rect 5365 9537 5399 9571
rect 7573 9537 7607 9571
rect 9873 9537 9907 9571
rect 11345 9537 11379 9571
rect 4169 9469 4203 9503
rect 11069 9469 11103 9503
rect 11161 9469 11195 9503
rect 1961 9401 1995 9435
rect 3065 9401 3099 9435
rect 5089 9401 5123 9435
rect 6101 9401 6135 9435
rect 7113 9401 7147 9435
rect 7840 9401 7874 9435
rect 12173 9401 12207 9435
rect 14473 9605 14507 9639
rect 20269 9605 20303 9639
rect 25145 9605 25179 9639
rect 25421 9605 25455 9639
rect 15485 9537 15519 9571
rect 18061 9537 18095 9571
rect 20913 9537 20947 9571
rect 22661 9537 22695 9571
rect 25789 9537 25823 9571
rect 13185 9469 13219 9503
rect 15577 9469 15611 9503
rect 15844 9469 15878 9503
rect 20637 9469 20671 9503
rect 22385 9469 22419 9503
rect 23765 9469 23799 9503
rect 18306 9401 18340 9435
rect 20729 9401 20763 9435
rect 23489 9401 23523 9435
rect 24010 9401 24044 9435
rect 2053 9333 2087 9367
rect 2697 9333 2731 9367
rect 3157 9333 3191 9367
rect 3525 9333 3559 9367
rect 3617 9333 3651 9367
rect 5181 9333 5215 9367
rect 7481 9333 7515 9367
rect 8953 9333 8987 9367
rect 9321 9333 9355 9367
rect 10701 9333 10735 9367
rect 11805 9333 11839 9367
rect 12909 9333 12943 9367
rect 13001 9333 13035 9367
rect 17785 9333 17819 9367
rect 19441 9333 19475 9367
rect 20177 9333 20211 9367
rect 21281 9333 21315 9367
rect 21649 9333 21683 9367
rect 22017 9333 22051 9367
rect 22477 9333 22511 9367
rect 23029 9333 23063 9367
rect 2237 9129 2271 9163
rect 2421 9129 2455 9163
rect 4169 9129 4203 9163
rect 6193 9129 6227 9163
rect 6837 9129 6871 9163
rect 9045 9129 9079 9163
rect 10609 9129 10643 9163
rect 12909 9129 12943 9163
rect 15025 9129 15059 9163
rect 15669 9129 15703 9163
rect 15761 9129 15795 9163
rect 16865 9129 16899 9163
rect 17325 9129 17359 9163
rect 18337 9129 18371 9163
rect 19257 9129 19291 9163
rect 20637 9129 20671 9163
rect 21097 9129 21131 9163
rect 22937 9129 22971 9163
rect 23949 9129 23983 9163
rect 24869 9129 24903 9163
rect 25237 9129 25271 9163
rect 25605 9129 25639 9163
rect 1409 9061 1443 9095
rect 4629 9061 4663 9095
rect 10946 9061 10980 9095
rect 16773 9061 16807 9095
rect 17233 9061 17267 9095
rect 20361 9061 20395 9095
rect 21741 9061 21775 9095
rect 1961 8993 1995 9027
rect 2789 8993 2823 9027
rect 4537 8993 4571 9027
rect 6101 8993 6135 9027
rect 7297 8993 7331 9027
rect 7564 8993 7598 9027
rect 9689 8993 9723 9027
rect 10701 8993 10735 9027
rect 13369 8993 13403 9027
rect 13625 8993 13659 9027
rect 19625 8993 19659 9027
rect 19717 8993 19751 9027
rect 23857 8993 23891 9027
rect 25053 8993 25087 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 4813 8925 4847 8959
rect 6377 8925 6411 8959
rect 12449 8925 12483 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 15853 8925 15887 8959
rect 17417 8925 17451 8959
rect 18797 8925 18831 8959
rect 19901 8925 19935 8959
rect 21833 8925 21867 8959
rect 21925 8925 21959 8959
rect 24041 8925 24075 8959
rect 3801 8857 3835 8891
rect 5733 8857 5767 8891
rect 7113 8857 7147 8891
rect 14749 8857 14783 8891
rect 23305 8857 23339 8891
rect 3249 8789 3283 8823
rect 3525 8789 3559 8823
rect 5273 8789 5307 8823
rect 5549 8789 5583 8823
rect 8677 8789 8711 8823
rect 9413 8789 9447 8823
rect 10241 8789 10275 8823
rect 12081 8789 12115 8823
rect 12541 8789 12575 8823
rect 15301 8789 15335 8823
rect 16405 8789 16439 8823
rect 17969 8789 18003 8823
rect 19073 8789 19107 8823
rect 21373 8789 21407 8823
rect 22477 8789 22511 8823
rect 23489 8789 23523 8823
rect 24501 8789 24535 8823
rect 1777 8585 1811 8619
rect 3249 8585 3283 8619
rect 4721 8585 4755 8619
rect 4905 8585 4939 8619
rect 7021 8585 7055 8619
rect 8769 8585 8803 8619
rect 10333 8585 10367 8619
rect 11897 8585 11931 8619
rect 12173 8585 12207 8619
rect 12633 8585 12667 8619
rect 13185 8585 13219 8619
rect 15393 8585 15427 8619
rect 17325 8585 17359 8619
rect 17693 8585 17727 8619
rect 18705 8585 18739 8619
rect 20177 8585 20211 8619
rect 20913 8585 20947 8619
rect 22385 8585 22419 8619
rect 25053 8585 25087 8619
rect 25697 8585 25731 8619
rect 5917 8517 5951 8551
rect 6653 8517 6687 8551
rect 10793 8517 10827 8551
rect 5457 8449 5491 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 9413 8449 9447 8483
rect 9505 8449 9539 8483
rect 10701 8449 10735 8483
rect 11345 8449 11379 8483
rect 16773 8449 16807 8483
rect 23673 8449 23707 8483
rect 25329 8449 25363 8483
rect 1869 8381 1903 8415
rect 2136 8381 2170 8415
rect 4261 8381 4295 8415
rect 9321 8381 9355 8415
rect 11161 8381 11195 8415
rect 11253 8381 11287 8415
rect 12449 8381 12483 8415
rect 13553 8381 13587 8415
rect 13820 8381 13854 8415
rect 15761 8381 15795 8415
rect 16681 8381 16715 8415
rect 18797 8381 18831 8415
rect 20453 8381 20487 8415
rect 21005 8381 21039 8415
rect 23489 8381 23523 8415
rect 3525 8313 3559 8347
rect 5365 8313 5399 8347
rect 8493 8313 8527 8347
rect 16129 8313 16163 8347
rect 18245 8313 18279 8347
rect 19042 8313 19076 8347
rect 21250 8313 21284 8347
rect 22753 8313 22787 8347
rect 23940 8313 23974 8347
rect 5273 8245 5307 8279
rect 7389 8245 7423 8279
rect 8033 8245 8067 8279
rect 8953 8245 8987 8279
rect 14933 8245 14967 8279
rect 16221 8245 16255 8279
rect 16589 8245 16623 8279
rect 23121 8245 23155 8279
rect 26065 8245 26099 8279
rect 1961 8041 1995 8075
rect 2237 8041 2271 8075
rect 3893 8041 3927 8075
rect 4169 8041 4203 8075
rect 4537 8041 4571 8075
rect 5549 8041 5583 8075
rect 7021 8041 7055 8075
rect 8401 8041 8435 8075
rect 9229 8041 9263 8075
rect 10517 8041 10551 8075
rect 12357 8041 12391 8075
rect 12817 8041 12851 8075
rect 13185 8041 13219 8075
rect 14289 8041 14323 8075
rect 16129 8041 16163 8075
rect 17693 8041 17727 8075
rect 19349 8041 19383 8075
rect 20085 8041 20119 8075
rect 20545 8041 20579 8075
rect 22293 8041 22327 8075
rect 23397 8041 23431 8075
rect 24685 8041 24719 8075
rect 25605 8041 25639 8075
rect 5273 7973 5307 8007
rect 7481 7973 7515 8007
rect 2789 7905 2823 7939
rect 3525 7905 3559 7939
rect 5917 7905 5951 7939
rect 7389 7905 7423 7939
rect 8033 7905 8067 7939
rect 9873 7905 9907 7939
rect 11244 7905 11278 7939
rect 1409 7837 1443 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 6561 7837 6595 7871
rect 7665 7837 7699 7871
rect 8585 7837 8619 7871
rect 10977 7837 11011 7871
rect 2421 7769 2455 7803
rect 13645 7973 13679 8007
rect 15761 7973 15795 8007
rect 16580 7973 16614 8007
rect 18613 7973 18647 8007
rect 22201 7973 22235 8007
rect 22937 7973 22971 8007
rect 13093 7905 13127 7939
rect 13553 7905 13587 7939
rect 18889 7905 18923 7939
rect 20729 7905 20763 7939
rect 23765 7905 23799 7939
rect 24961 7905 24995 7939
rect 13737 7837 13771 7871
rect 15301 7837 15335 7871
rect 16313 7837 16347 7871
rect 19441 7837 19475 7871
rect 19533 7837 19567 7871
rect 22477 7837 22511 7871
rect 23305 7837 23339 7871
rect 23857 7837 23891 7871
rect 23949 7837 23983 7871
rect 18981 7769 19015 7803
rect 20361 7769 20395 7803
rect 6101 7701 6135 7735
rect 6929 7701 6963 7735
rect 10057 7701 10091 7735
rect 10885 7701 10919 7735
rect 12633 7701 12667 7735
rect 12817 7701 12851 7735
rect 14657 7701 14691 7735
rect 14933 7701 14967 7735
rect 18153 7701 18187 7735
rect 18705 7701 18739 7735
rect 21465 7701 21499 7735
rect 21833 7701 21867 7735
rect 25145 7701 25179 7735
rect 2329 7497 2363 7531
rect 3985 7497 4019 7531
rect 4721 7497 4755 7531
rect 6929 7497 6963 7531
rect 8033 7497 8067 7531
rect 8677 7497 8711 7531
rect 10333 7497 10367 7531
rect 10793 7497 10827 7531
rect 12265 7497 12299 7531
rect 15669 7497 15703 7531
rect 17785 7497 17819 7531
rect 19073 7497 19107 7531
rect 19441 7497 19475 7531
rect 19901 7497 19935 7531
rect 21925 7497 21959 7531
rect 22845 7497 22879 7531
rect 23121 7497 23155 7531
rect 23489 7497 23523 7531
rect 24593 7497 24627 7531
rect 25973 7497 26007 7531
rect 1961 7429 1995 7463
rect 6561 7429 6595 7463
rect 16037 7429 16071 7463
rect 21557 7429 21591 7463
rect 3065 7361 3099 7395
rect 3433 7361 3467 7395
rect 4169 7361 4203 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 9137 7361 9171 7395
rect 9781 7361 9815 7395
rect 11437 7361 11471 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 18705 7361 18739 7395
rect 20453 7361 20487 7395
rect 22661 7361 22695 7395
rect 25053 7361 25087 7395
rect 25145 7361 25179 7395
rect 2789 7293 2823 7327
rect 7297 7293 7331 7327
rect 9597 7293 9631 7327
rect 12449 7293 12483 7327
rect 13553 7293 13587 7327
rect 13820 7293 13854 7327
rect 15301 7293 15335 7327
rect 16313 7293 16347 7327
rect 18521 7293 18555 7327
rect 20361 7293 20395 7327
rect 22385 7293 22419 7327
rect 22845 7293 22879 7327
rect 5089 7225 5123 7259
rect 5549 7225 5583 7259
rect 11253 7225 11287 7259
rect 16773 7225 16807 7259
rect 17417 7225 17451 7259
rect 18429 7225 18463 7259
rect 24041 7225 24075 7259
rect 1409 7157 1443 7191
rect 2421 7157 2455 7191
rect 2881 7157 2915 7191
rect 5181 7157 5215 7191
rect 6285 7157 6319 7191
rect 8309 7157 8343 7191
rect 9229 7157 9263 7191
rect 9689 7157 9723 7191
rect 10701 7157 10735 7191
rect 11161 7157 11195 7191
rect 11805 7157 11839 7191
rect 12633 7157 12667 7191
rect 13185 7157 13219 7191
rect 14933 7157 14967 7191
rect 16129 7157 16163 7191
rect 16405 7157 16439 7191
rect 18061 7157 18095 7191
rect 20269 7157 20303 7191
rect 20913 7157 20947 7191
rect 22017 7157 22051 7191
rect 22477 7157 22511 7191
rect 24501 7157 24535 7191
rect 24961 7157 24995 7191
rect 25605 7157 25639 7191
rect 2973 6953 3007 6987
rect 5089 6953 5123 6987
rect 6101 6953 6135 6987
rect 7021 6953 7055 6987
rect 11713 6953 11747 6987
rect 12541 6953 12575 6987
rect 13277 6953 13311 6987
rect 16681 6953 16715 6987
rect 17049 6953 17083 6987
rect 19625 6953 19659 6987
rect 20361 6953 20395 6987
rect 22569 6953 22603 6987
rect 2053 6885 2087 6919
rect 5457 6885 5491 6919
rect 4077 6817 4111 6851
rect 4629 6817 4663 6851
rect 8401 6817 8435 6851
rect 8493 6817 8527 6851
rect 9321 6817 9355 6851
rect 10221 6817 10255 6851
rect 12633 6817 12667 6851
rect 13921 6817 13955 6851
rect 15301 6817 15335 6851
rect 16405 6817 16439 6851
rect 17785 6817 17819 6851
rect 19073 6817 19107 6851
rect 19717 6817 19751 6851
rect 20913 6817 20947 6851
rect 21180 6817 21214 6851
rect 23029 6817 23063 6851
rect 23388 6817 23422 6851
rect 25329 6817 25363 6851
rect 2145 6749 2179 6783
rect 2329 6749 2363 6783
rect 4905 6749 4939 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 7113 6749 7147 6783
rect 7297 6749 7331 6783
rect 9965 6749 9999 6783
rect 12725 6749 12759 6783
rect 13645 6749 13679 6783
rect 14105 6749 14139 6783
rect 15485 6749 15519 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 18245 6749 18279 6783
rect 19901 6749 19935 6783
rect 23121 6749 23155 6783
rect 1685 6681 1719 6715
rect 11989 6681 12023 6715
rect 12173 6681 12207 6715
rect 19257 6681 19291 6715
rect 24777 6681 24811 6715
rect 3341 6613 3375 6647
rect 3893 6613 3927 6647
rect 6561 6613 6595 6647
rect 6653 6613 6687 6647
rect 7665 6613 7699 6647
rect 8033 6613 8067 6647
rect 8217 6613 8251 6647
rect 8677 6613 8711 6647
rect 11345 6613 11379 6647
rect 14749 6613 14783 6647
rect 15117 6613 15151 6647
rect 18061 6613 18095 6647
rect 20729 6613 20763 6647
rect 22293 6613 22327 6647
rect 24501 6613 24535 6647
rect 25145 6613 25179 6647
rect 25513 6613 25547 6647
rect 2053 6409 2087 6443
rect 5181 6409 5215 6443
rect 6285 6409 6319 6443
rect 6653 6409 6687 6443
rect 7941 6409 7975 6443
rect 8585 6409 8619 6443
rect 8861 6409 8895 6443
rect 10425 6409 10459 6443
rect 10701 6409 10735 6443
rect 11161 6409 11195 6443
rect 11897 6409 11931 6443
rect 17141 6409 17175 6443
rect 17785 6409 17819 6443
rect 18521 6409 18555 6443
rect 20269 6409 20303 6443
rect 20821 6409 20855 6443
rect 21833 6409 21867 6443
rect 23673 6409 23707 6443
rect 25053 6409 25087 6443
rect 26341 6409 26375 6443
rect 4077 6341 4111 6375
rect 13737 6341 13771 6375
rect 17509 6341 17543 6375
rect 20729 6341 20763 6375
rect 3433 6273 3467 6307
rect 4445 6273 4479 6307
rect 5641 6273 5675 6307
rect 5733 6273 5767 6307
rect 7389 6273 7423 6307
rect 13645 6273 13679 6307
rect 14381 6273 14415 6307
rect 21281 6273 21315 6307
rect 21373 6273 21407 6307
rect 22201 6273 22235 6307
rect 24133 6273 24167 6307
rect 24317 6273 24351 6307
rect 24685 6273 24719 6307
rect 25421 6273 25455 6307
rect 1409 6205 1443 6239
rect 3341 6205 3375 6239
rect 5089 6205 5123 6239
rect 5549 6205 5583 6239
rect 7297 6205 7331 6239
rect 9052 6205 9086 6239
rect 9301 6205 9335 6239
rect 11253 6205 11287 6239
rect 12449 6205 12483 6239
rect 13185 6205 13219 6239
rect 15761 6205 15795 6239
rect 18613 6205 18647 6239
rect 21189 6205 21223 6239
rect 22385 6205 22419 6239
rect 24041 6205 24075 6239
rect 25237 6205 25271 6239
rect 2789 6137 2823 6171
rect 4813 6137 4847 6171
rect 12725 6137 12759 6171
rect 14105 6137 14139 6171
rect 15117 6137 15151 6171
rect 15669 6137 15703 6171
rect 16006 6137 16040 6171
rect 18858 6137 18892 6171
rect 1593 6069 1627 6103
rect 2421 6069 2455 6103
rect 2881 6069 2915 6103
rect 3249 6069 3283 6103
rect 4905 6069 4939 6103
rect 6837 6069 6871 6103
rect 7205 6069 7239 6103
rect 11437 6069 11471 6103
rect 12173 6069 12207 6103
rect 14197 6069 14231 6103
rect 14749 6069 14783 6103
rect 19993 6069 20027 6103
rect 22569 6069 22603 6103
rect 23213 6069 23247 6103
rect 25973 6069 26007 6103
rect 3709 5865 3743 5899
rect 5457 5865 5491 5899
rect 6377 5865 6411 5899
rect 7849 5865 7883 5899
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 9137 5865 9171 5899
rect 10333 5865 10367 5899
rect 11989 5865 12023 5899
rect 13369 5865 13403 5899
rect 13645 5865 13679 5899
rect 14013 5865 14047 5899
rect 14105 5865 14139 5899
rect 15117 5865 15151 5899
rect 17049 5865 17083 5899
rect 20913 5865 20947 5899
rect 22385 5865 22419 5899
rect 24041 5865 24075 5899
rect 25053 5865 25087 5899
rect 25421 5865 25455 5899
rect 25789 5865 25823 5899
rect 3341 5797 3375 5831
rect 8309 5797 8343 5831
rect 15546 5797 15580 5831
rect 24409 5797 24443 5831
rect 1685 5729 1719 5763
rect 1952 5729 1986 5763
rect 4077 5729 4111 5763
rect 4333 5729 4367 5763
rect 6736 5729 6770 5763
rect 9321 5729 9355 5763
rect 11897 5729 11931 5763
rect 17417 5729 17451 5763
rect 17785 5729 17819 5763
rect 18337 5729 18371 5763
rect 18604 5729 18638 5763
rect 21281 5729 21315 5763
rect 21925 5729 21959 5763
rect 22845 5729 22879 5763
rect 22937 5729 22971 5763
rect 6469 5661 6503 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 12081 5661 12115 5695
rect 12541 5661 12575 5695
rect 14197 5661 14231 5695
rect 14657 5661 14691 5695
rect 15301 5661 15335 5695
rect 20729 5661 20763 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 23121 5661 23155 5695
rect 24501 5661 24535 5695
rect 24685 5661 24719 5695
rect 9965 5593 9999 5627
rect 11529 5593 11563 5627
rect 13093 5593 13127 5627
rect 3065 5525 3099 5559
rect 5825 5525 5859 5559
rect 10977 5525 11011 5559
rect 11437 5525 11471 5559
rect 16681 5525 16715 5559
rect 18245 5525 18279 5559
rect 19717 5525 19751 5559
rect 20085 5525 20119 5559
rect 22477 5525 22511 5559
rect 23673 5525 23707 5559
rect 3709 5321 3743 5355
rect 4353 5321 4387 5355
rect 5917 5321 5951 5355
rect 6285 5321 6319 5355
rect 7297 5321 7331 5355
rect 8309 5321 8343 5355
rect 9781 5321 9815 5355
rect 10793 5321 10827 5355
rect 12173 5321 12207 5355
rect 12909 5321 12943 5355
rect 13369 5321 13403 5355
rect 14933 5321 14967 5355
rect 15761 5321 15795 5355
rect 16865 5321 16899 5355
rect 18705 5321 18739 5355
rect 20637 5321 20671 5355
rect 21557 5321 21591 5355
rect 22937 5321 22971 5355
rect 23305 5321 23339 5355
rect 25053 5321 25087 5355
rect 25329 5321 25363 5355
rect 25697 5321 25731 5355
rect 26065 5321 26099 5355
rect 4077 5253 4111 5287
rect 9689 5253 9723 5287
rect 14473 5253 14507 5287
rect 18245 5253 18279 5287
rect 2329 5185 2363 5219
rect 6653 5185 6687 5219
rect 7757 5185 7791 5219
rect 7941 5185 7975 5219
rect 10333 5185 10367 5219
rect 11345 5185 11379 5219
rect 13829 5185 13863 5219
rect 14013 5185 14047 5219
rect 16313 5185 16347 5219
rect 16497 5185 16531 5219
rect 19165 5185 19199 5219
rect 22109 5185 22143 5219
rect 22661 5185 22695 5219
rect 4537 5117 4571 5151
rect 4793 5117 4827 5151
rect 9321 5117 9355 5151
rect 10241 5117 10275 5151
rect 15393 5117 15427 5151
rect 16221 5117 16255 5151
rect 18061 5117 18095 5151
rect 19257 5117 19291 5151
rect 19524 5117 19558 5151
rect 21097 5117 21131 5151
rect 21925 5117 21959 5151
rect 23673 5117 23707 5151
rect 2596 5049 2630 5083
rect 8953 5049 8987 5083
rect 10149 5049 10183 5083
rect 11805 5049 11839 5083
rect 13277 5049 13311 5083
rect 13737 5049 13771 5083
rect 17785 5049 17819 5083
rect 23918 5049 23952 5083
rect 1685 4981 1719 5015
rect 2053 4981 2087 5015
rect 7205 4981 7239 5015
rect 7665 4981 7699 5015
rect 11161 4981 11195 5015
rect 15853 4981 15887 5015
rect 17325 4981 17359 5015
rect 21465 4981 21499 5015
rect 22017 4981 22051 5015
rect 4997 4777 5031 4811
rect 5365 4777 5399 4811
rect 6009 4777 6043 4811
rect 7481 4777 7515 4811
rect 9505 4777 9539 4811
rect 11069 4777 11103 4811
rect 12173 4777 12207 4811
rect 14013 4777 14047 4811
rect 14289 4777 14323 4811
rect 17785 4777 17819 4811
rect 18245 4777 18279 4811
rect 20637 4777 20671 4811
rect 22017 4777 22051 4811
rect 22937 4777 22971 4811
rect 23673 4777 23707 4811
rect 25053 4777 25087 4811
rect 25513 4777 25547 4811
rect 12510 4709 12544 4743
rect 15844 4709 15878 4743
rect 19625 4709 19659 4743
rect 1961 4641 1995 4675
rect 2053 4641 2087 4675
rect 4445 4641 4479 4675
rect 5917 4641 5951 4675
rect 7573 4641 7607 4675
rect 9137 4641 9171 4675
rect 9689 4641 9723 4675
rect 9956 4641 9990 4675
rect 15577 4641 15611 4675
rect 18153 4641 18187 4675
rect 19349 4641 19383 4675
rect 20085 4641 20119 4675
rect 21281 4641 21315 4675
rect 22845 4641 22879 4675
rect 24409 4641 24443 4675
rect 2237 4573 2271 4607
rect 6193 4573 6227 4607
rect 7757 4573 7791 4607
rect 8125 4573 8159 4607
rect 12265 4573 12299 4607
rect 18429 4573 18463 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 23029 4573 23063 4607
rect 24501 4573 24535 4607
rect 24593 4573 24627 4607
rect 3617 4505 3651 4539
rect 22385 4505 22419 4539
rect 1593 4437 1627 4471
rect 2605 4437 2639 4471
rect 3341 4437 3375 4471
rect 4261 4437 4295 4471
rect 4629 4437 4663 4471
rect 5549 4437 5583 4471
rect 6929 4437 6963 4471
rect 7113 4437 7147 4471
rect 8677 4437 8711 4471
rect 11437 4437 11471 4471
rect 11805 4437 11839 4471
rect 13645 4437 13679 4471
rect 14749 4437 14783 4471
rect 15117 4437 15151 4471
rect 16957 4437 16991 4471
rect 17325 4437 17359 4471
rect 17693 4437 17727 4471
rect 18889 4437 18923 4471
rect 19165 4437 19199 4471
rect 20913 4437 20947 4471
rect 22477 4437 22511 4471
rect 24041 4437 24075 4471
rect 1501 4233 1535 4267
rect 2881 4233 2915 4267
rect 4629 4233 4663 4267
rect 4997 4233 5031 4267
rect 5365 4233 5399 4267
rect 6193 4233 6227 4267
rect 8217 4233 8251 4267
rect 9873 4233 9907 4267
rect 10885 4233 10919 4267
rect 11253 4233 11287 4267
rect 15393 4233 15427 4267
rect 15669 4233 15703 4267
rect 22753 4233 22787 4267
rect 23489 4233 23523 4267
rect 24685 4233 24719 4267
rect 6837 4165 6871 4199
rect 19165 4165 19199 4199
rect 1961 4097 1995 4131
rect 2145 4097 2179 4131
rect 5733 4097 5767 4131
rect 7389 4097 7423 4131
rect 10517 4097 10551 4131
rect 13001 4097 13035 4131
rect 13829 4097 13863 4131
rect 14565 4097 14599 4131
rect 16405 4097 16439 4131
rect 17417 4097 17451 4131
rect 18613 4097 18647 4131
rect 19901 4097 19935 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 24225 4097 24259 4131
rect 25053 4097 25087 4131
rect 25513 4097 25547 4131
rect 26341 4097 26375 4131
rect 1869 4029 1903 4063
rect 3249 4029 3283 4063
rect 5457 4029 5491 4063
rect 6561 4029 6595 4063
rect 7297 4029 7331 4063
rect 7941 4029 7975 4063
rect 8585 4029 8619 4063
rect 10241 4029 10275 4063
rect 12265 4029 12299 4063
rect 12817 4029 12851 4063
rect 14381 4029 14415 4063
rect 16313 4029 16347 4063
rect 17785 4029 17819 4063
rect 18521 4029 18555 4063
rect 19625 4029 19659 4063
rect 24041 4029 24075 4063
rect 25237 4029 25271 4063
rect 25973 4029 26007 4063
rect 3516 3961 3550 3995
rect 8861 3961 8895 3995
rect 10333 3961 10367 3995
rect 13461 3961 13495 3995
rect 14473 3961 14507 3995
rect 16221 3961 16255 3995
rect 17049 3961 17083 3995
rect 18429 3961 18463 3995
rect 20913 3961 20947 3995
rect 21272 3961 21306 3995
rect 2513 3893 2547 3927
rect 7205 3893 7239 3927
rect 9321 3893 9355 3927
rect 9781 3893 9815 3927
rect 11897 3893 11931 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 14013 3893 14047 3927
rect 15853 3893 15887 3927
rect 18061 3893 18095 3927
rect 19441 3893 19475 3927
rect 22385 3893 22419 3927
rect 23121 3893 23155 3927
rect 23673 3893 23707 3927
rect 24133 3893 24167 3927
rect 1501 3689 1535 3723
rect 2605 3689 2639 3723
rect 4537 3689 4571 3723
rect 5181 3689 5215 3723
rect 7113 3689 7147 3723
rect 7941 3689 7975 3723
rect 11069 3689 11103 3723
rect 11529 3689 11563 3723
rect 11989 3689 12023 3723
rect 12817 3689 12851 3723
rect 12909 3689 12943 3723
rect 15485 3689 15519 3723
rect 15853 3689 15887 3723
rect 16865 3689 16899 3723
rect 18153 3689 18187 3723
rect 18521 3689 18555 3723
rect 19717 3689 19751 3723
rect 21189 3689 21223 3723
rect 21465 3689 21499 3723
rect 24041 3689 24075 3723
rect 25513 3689 25547 3723
rect 1961 3621 1995 3655
rect 5457 3621 5491 3655
rect 6000 3621 6034 3655
rect 7389 3621 7423 3655
rect 8953 3621 8987 3655
rect 13461 3621 13495 3655
rect 15117 3621 15151 3655
rect 15945 3621 15979 3655
rect 17417 3621 17451 3655
rect 18889 3621 18923 3655
rect 22100 3621 22134 3655
rect 24501 3621 24535 3655
rect 1869 3553 1903 3587
rect 4445 3553 4479 3587
rect 5733 3553 5767 3587
rect 8309 3553 8343 3587
rect 9689 3553 9723 3587
rect 9956 3553 9990 3587
rect 14013 3553 14047 3587
rect 19625 3553 19659 3587
rect 21833 3553 21867 3587
rect 24409 3553 24443 3587
rect 2145 3485 2179 3519
rect 3433 3485 3467 3519
rect 3893 3485 3927 3519
rect 4721 3485 4755 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 13093 3485 13127 3519
rect 16037 3485 16071 3519
rect 17509 3485 17543 3519
rect 17693 3485 17727 3519
rect 19901 3485 19935 3519
rect 24593 3485 24627 3519
rect 2973 3417 3007 3451
rect 4077 3417 4111 3451
rect 7849 3417 7883 3451
rect 12449 3417 12483 3451
rect 14749 3417 14783 3451
rect 19257 3417 19291 3451
rect 23213 3417 23247 3451
rect 25053 3417 25087 3451
rect 9321 3349 9355 3383
rect 12357 3349 12391 3383
rect 13921 3349 13955 3383
rect 14197 3349 14231 3383
rect 16589 3349 16623 3383
rect 17049 3349 17083 3383
rect 20361 3349 20395 3383
rect 20729 3349 20763 3383
rect 23765 3349 23799 3383
rect 1685 3145 1719 3179
rect 2053 3145 2087 3179
rect 3065 3145 3099 3179
rect 5273 3145 5307 3179
rect 5825 3145 5859 3179
rect 6193 3145 6227 3179
rect 8309 3145 8343 3179
rect 10149 3145 10183 3179
rect 10425 3145 10459 3179
rect 10977 3145 11011 3179
rect 11897 3145 11931 3179
rect 13829 3145 13863 3179
rect 15761 3145 15795 3179
rect 16129 3145 16163 3179
rect 17325 3145 17359 3179
rect 18337 3145 18371 3179
rect 20177 3145 20211 3179
rect 22017 3145 22051 3179
rect 22293 3145 22327 3179
rect 22753 3145 22787 3179
rect 23121 3145 23155 3179
rect 25053 3145 25087 3179
rect 25329 3145 25363 3179
rect 25697 3145 25731 3179
rect 3433 3077 3467 3111
rect 6377 3077 6411 3111
rect 6653 3077 6687 3111
rect 8033 3077 8067 3111
rect 16221 3077 16255 3111
rect 19809 3077 19843 3111
rect 20453 3077 20487 3111
rect 26065 3077 26099 3111
rect 2605 3009 2639 3043
rect 3617 3009 3651 3043
rect 2421 2941 2455 2975
rect 3884 2873 3918 2907
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 8769 3009 8803 3043
rect 11345 3009 11379 3043
rect 14105 3009 14139 3043
rect 14565 3009 14599 3043
rect 15209 3009 15243 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 23397 3009 23431 3043
rect 7205 2941 7239 2975
rect 11069 2941 11103 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 15025 2941 15059 2975
rect 18429 2941 18463 2975
rect 20637 2941 20671 2975
rect 20893 2941 20927 2975
rect 23673 2941 23707 2975
rect 23929 2941 23963 2975
rect 9014 2873 9048 2907
rect 15117 2873 15151 2907
rect 16589 2873 16623 2907
rect 18696 2873 18730 2907
rect 2513 2805 2547 2839
rect 4997 2805 5031 2839
rect 6377 2805 6411 2839
rect 6837 2805 6871 2839
rect 12265 2805 12299 2839
rect 14657 2805 14691 2839
rect 17601 2805 17635 2839
rect 1409 2601 1443 2635
rect 1869 2601 1903 2635
rect 2237 2601 2271 2635
rect 2421 2601 2455 2635
rect 2789 2601 2823 2635
rect 5181 2601 5215 2635
rect 6377 2601 6411 2635
rect 6745 2601 6779 2635
rect 7757 2601 7791 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 11253 2601 11287 2635
rect 12081 2601 12115 2635
rect 14565 2601 14599 2635
rect 15945 2601 15979 2635
rect 16589 2601 16623 2635
rect 17785 2601 17819 2635
rect 18337 2601 18371 2635
rect 19809 2601 19843 2635
rect 21189 2601 21223 2635
rect 21557 2601 21591 2635
rect 22293 2601 22327 2635
rect 24041 2601 24075 2635
rect 25053 2601 25087 2635
rect 25605 2601 25639 2635
rect 3433 2533 3467 2567
rect 4445 2533 4479 2567
rect 9597 2533 9631 2567
rect 12449 2533 12483 2567
rect 12900 2533 12934 2567
rect 14841 2533 14875 2567
rect 15853 2533 15887 2567
rect 20913 2533 20947 2567
rect 25513 2533 25547 2567
rect 2881 2465 2915 2499
rect 5733 2465 5767 2499
rect 7665 2465 7699 2499
rect 8125 2465 8159 2499
rect 8217 2465 8251 2499
rect 11437 2465 11471 2499
rect 15209 2465 15243 2499
rect 17049 2465 17083 2499
rect 18061 2465 18095 2499
rect 18705 2465 18739 2499
rect 20545 2465 20579 2499
rect 24409 2465 24443 2499
rect 2973 2397 3007 2431
rect 4537 2397 4571 2431
rect 4721 2397 4755 2431
rect 7297 2397 7331 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 12633 2397 12667 2431
rect 16037 2397 16071 2431
rect 18797 2397 18831 2431
rect 18889 2397 18923 2431
rect 19349 2397 19383 2431
rect 21649 2397 21683 2431
rect 21741 2397 21775 2431
rect 24501 2397 24535 2431
rect 24685 2397 24719 2431
rect 4077 2329 4111 2363
rect 5549 2329 5583 2363
rect 10885 2329 10919 2363
rect 15485 2329 15519 2363
rect 17233 2329 17267 2363
rect 23489 2329 23523 2363
rect 3801 2261 3835 2295
rect 5917 2261 5951 2295
rect 8861 2261 8895 2295
rect 11621 2261 11655 2295
rect 14013 2261 14047 2295
rect 16865 2261 16899 2295
rect 20177 2261 20211 2295
rect 22569 2261 22603 2295
rect 23029 2261 23063 2295
rect 23765 2261 23799 2295
<< metal1 >>
rect 3694 25984 3700 26036
rect 3752 26024 3758 26036
rect 8294 26024 8300 26036
rect 3752 25996 8300 26024
rect 3752 25984 3758 25996
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 24118 25168 24124 25220
rect 24176 25208 24182 25220
rect 24486 25208 24492 25220
rect 24176 25180 24492 25208
rect 24176 25168 24182 25180
rect 24486 25168 24492 25180
rect 24544 25168 24550 25220
rect 4062 25100 4068 25152
rect 4120 25140 4126 25152
rect 5534 25140 5540 25152
rect 4120 25112 5540 25140
rect 4120 25100 4126 25112
rect 5534 25100 5540 25112
rect 5592 25100 5598 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5592 23820 5825 23848
rect 5592 23808 5598 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 24210 23808 24216 23860
rect 24268 23848 24274 23860
rect 24765 23851 24823 23857
rect 24765 23848 24777 23851
rect 24268 23820 24777 23848
rect 24268 23808 24274 23820
rect 24765 23817 24777 23820
rect 24811 23817 24823 23851
rect 24765 23811 24823 23817
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23644 5687 23647
rect 5675 23616 6316 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 6288 23517 6316 23616
rect 24118 23604 24124 23656
rect 24176 23644 24182 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24176 23616 24593 23644
rect 24176 23604 24182 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 6273 23511 6331 23517
rect 6273 23477 6285 23511
rect 6319 23508 6331 23511
rect 6822 23508 6828 23520
rect 6319 23480 6828 23508
rect 6319 23477 6331 23480
rect 6273 23471 6331 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 24854 23304 24860 23316
rect 24811 23276 24860 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 24670 22760 24676 22772
rect 23952 22732 24676 22760
rect 23952 22633 23980 22732
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 25133 22763 25191 22769
rect 25133 22760 25145 22763
rect 24912 22732 25145 22760
rect 24912 22720 24918 22732
rect 25133 22729 25145 22732
rect 25179 22729 25191 22763
rect 25133 22723 25191 22729
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 23661 22559 23719 22565
rect 23661 22556 23673 22559
rect 1443 22528 2084 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2056 22432 2084 22528
rect 23492 22528 23673 22556
rect 23492 22432 23520 22528
rect 23661 22525 23673 22528
rect 23707 22525 23719 22559
rect 24946 22556 24952 22568
rect 24907 22528 24952 22556
rect 23661 22519 23719 22525
rect 24946 22516 24952 22528
rect 25004 22556 25010 22568
rect 25501 22559 25559 22565
rect 25501 22556 25513 22559
rect 25004 22528 25513 22556
rect 25004 22516 25010 22528
rect 25501 22525 25513 22528
rect 25547 22525 25559 22559
rect 25501 22519 25559 22525
rect 2038 22420 2044 22432
rect 1999 22392 2044 22420
rect 2038 22380 2044 22392
rect 2096 22380 2102 22432
rect 23474 22420 23480 22432
rect 23435 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 2084 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2056 21344 2084 21440
rect 2038 21332 2044 21344
rect 1999 21304 2044 21332
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 21726 21128 21732 21140
rect 21687 21100 21732 21128
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 2038 21060 2044 21072
rect 1999 21032 2044 21060
rect 2038 21020 2044 21032
rect 2096 21020 2102 21072
rect 1765 20995 1823 21001
rect 1765 20961 1777 20995
rect 1811 20992 1823 20995
rect 2314 20992 2320 21004
rect 1811 20964 2320 20992
rect 1811 20961 1823 20964
rect 1765 20955 1823 20961
rect 2314 20952 2320 20964
rect 2372 20952 2378 21004
rect 21542 20992 21548 21004
rect 21503 20964 21548 20992
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1486 20544 1492 20596
rect 1544 20584 1550 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1544 20556 1593 20584
rect 1544 20544 1550 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 21542 20584 21548 20596
rect 1581 20547 1639 20553
rect 20824 20556 21548 20584
rect 20824 20457 20852 20556
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 20364 20352 20545 20380
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 2314 20244 2320 20256
rect 2275 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 20364 20253 20392 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20349 20247 20407 20253
rect 20349 20244 20361 20247
rect 19392 20216 20361 20244
rect 19392 20204 19398 20216
rect 20349 20213 20361 20216
rect 20395 20213 20407 20247
rect 20349 20207 20407 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 24762 20040 24768 20052
rect 24723 20012 24768 20040
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2406 19904 2412 19916
rect 1443 19876 2412 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 24210 19864 24216 19916
rect 24268 19904 24274 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24268 19876 24593 19904
rect 24268 19864 24274 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1578 19292 1584 19304
rect 1443 19264 1584 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1578 19252 1584 19264
rect 1636 19292 1642 19304
rect 1949 19295 2007 19301
rect 1949 19292 1961 19295
rect 1636 19264 1961 19292
rect 1636 19252 1642 19264
rect 1949 19261 1961 19264
rect 1995 19261 2007 19295
rect 24578 19292 24584 19304
rect 24539 19264 24584 19292
rect 1949 19255 2007 19261
rect 24578 19252 24584 19264
rect 24636 19292 24642 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24636 19264 25145 19292
rect 24636 19252 24642 19264
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 1486 19116 1492 19168
rect 1544 19156 1550 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 1544 19128 1593 19156
rect 1544 19116 1550 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 2406 19156 2412 19168
rect 2367 19128 2412 19156
rect 1581 19119 1639 19125
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 24394 19156 24400 19168
rect 24355 19128 24400 19156
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 24670 19116 24676 19168
rect 24728 19156 24734 19168
rect 24765 19159 24823 19165
rect 24765 19156 24777 19159
rect 24728 19128 24777 19156
rect 24728 19116 24734 19128
rect 24765 19125 24777 19128
rect 24811 19125 24823 19159
rect 24765 19119 24823 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2682 18952 2688 18964
rect 2643 18924 2688 18952
rect 2682 18912 2688 18924
rect 2740 18912 2746 18964
rect 18230 18952 18236 18964
rect 18191 18924 18236 18952
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 4338 18884 4344 18896
rect 4299 18856 4344 18884
rect 4338 18844 4344 18856
rect 4396 18844 4402 18896
rect 23934 18844 23940 18896
rect 23992 18884 23998 18896
rect 25314 18884 25320 18896
rect 23992 18856 25320 18884
rect 23992 18844 23998 18856
rect 25314 18844 25320 18856
rect 25372 18844 25378 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2501 18819 2559 18825
rect 1443 18788 2452 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 2424 18621 2452 18788
rect 2501 18785 2513 18819
rect 2547 18816 2559 18819
rect 3142 18816 3148 18828
rect 2547 18788 3148 18816
rect 2547 18785 2559 18788
rect 2501 18779 2559 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4430 18816 4436 18828
rect 4111 18788 4436 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4430 18776 4436 18788
rect 4488 18776 4494 18828
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 18012 18788 18061 18816
rect 18012 18776 18018 18788
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 23474 18816 23480 18828
rect 23435 18788 23480 18816
rect 18049 18779 18107 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24210 18776 24216 18828
rect 24268 18816 24274 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24268 18788 24593 18816
rect 24268 18776 24274 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 22465 18751 22523 18757
rect 22465 18717 22477 18751
rect 22511 18748 22523 18751
rect 23290 18748 23296 18760
rect 22511 18720 23296 18748
rect 22511 18717 22523 18720
rect 22465 18711 22523 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1820 18584 1961 18612
rect 1820 18572 1826 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 1949 18575 2007 18581
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2958 18612 2964 18624
rect 2455 18584 2964 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 23661 18615 23719 18621
rect 23661 18581 23673 18615
rect 23707 18612 23719 18615
rect 24026 18612 24032 18624
rect 23707 18584 24032 18612
rect 23707 18581 23719 18584
rect 23661 18575 23719 18581
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 24762 18612 24768 18624
rect 24723 18584 24768 18612
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1452 18380 1593 18408
rect 1452 18368 1458 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 1581 18371 1639 18377
rect 24118 18368 24124 18420
rect 24176 18408 24182 18420
rect 24765 18411 24823 18417
rect 24765 18408 24777 18411
rect 24176 18380 24777 18408
rect 24176 18368 24182 18380
rect 24765 18377 24777 18380
rect 24811 18377 24823 18411
rect 24765 18371 24823 18377
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2501 18207 2559 18213
rect 2501 18204 2513 18207
rect 1443 18176 1992 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1964 18080 1992 18176
rect 2332 18176 2513 18204
rect 2332 18080 2360 18176
rect 2501 18173 2513 18176
rect 2547 18173 2559 18207
rect 2501 18167 2559 18173
rect 22465 18207 22523 18213
rect 22465 18173 22477 18207
rect 22511 18204 22523 18207
rect 24578 18204 24584 18216
rect 22511 18176 23152 18204
rect 24539 18176 24584 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2314 18068 2320 18080
rect 2275 18040 2320 18068
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 2685 18071 2743 18077
rect 2685 18037 2697 18071
rect 2731 18068 2743 18071
rect 2774 18068 2780 18080
rect 2731 18040 2780 18068
rect 2731 18037 2743 18040
rect 2685 18031 2743 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 3142 18068 3148 18080
rect 3055 18040 3148 18068
rect 3142 18028 3148 18040
rect 3200 18068 3206 18080
rect 3878 18068 3884 18080
rect 3200 18040 3884 18068
rect 3200 18028 3206 18040
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18068 4215 18071
rect 4430 18068 4436 18080
rect 4203 18040 4436 18068
rect 4203 18037 4215 18040
rect 4157 18031 4215 18037
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 18012 18040 18245 18068
rect 18012 18028 18018 18040
rect 18233 18037 18245 18040
rect 18279 18037 18291 18071
rect 18233 18031 18291 18037
rect 22649 18071 22707 18077
rect 22649 18037 22661 18071
rect 22695 18068 22707 18071
rect 23014 18068 23020 18080
rect 22695 18040 23020 18068
rect 22695 18037 22707 18040
rect 22649 18031 22707 18037
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 23124 18077 23152 18176
rect 24578 18164 24584 18176
rect 24636 18204 24642 18216
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24636 18176 25145 18204
rect 24636 18164 24642 18176
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 23198 18068 23204 18080
rect 23155 18040 23204 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 23532 18040 23857 18068
rect 23532 18028 23538 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 24210 18028 24216 18080
rect 24268 18068 24274 18080
rect 24397 18071 24455 18077
rect 24397 18068 24409 18071
rect 24268 18040 24409 18068
rect 24268 18028 24274 18040
rect 24397 18037 24409 18040
rect 24443 18037 24455 18071
rect 24397 18031 24455 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 4212 17836 4261 17864
rect 4212 17824 4218 17836
rect 4249 17833 4261 17836
rect 4295 17833 4307 17867
rect 4249 17827 4307 17833
rect 24670 17824 24676 17876
rect 24728 17864 24734 17876
rect 24765 17867 24823 17873
rect 24765 17864 24777 17867
rect 24728 17836 24777 17864
rect 24728 17824 24734 17836
rect 24765 17833 24777 17836
rect 24811 17833 24823 17867
rect 24765 17827 24823 17833
rect 1673 17799 1731 17805
rect 1673 17765 1685 17799
rect 1719 17796 1731 17799
rect 2314 17796 2320 17808
rect 1719 17768 2320 17796
rect 1719 17765 1731 17768
rect 1673 17759 1731 17765
rect 2314 17756 2320 17768
rect 2372 17756 2378 17808
rect 17405 17799 17463 17805
rect 17405 17765 17417 17799
rect 17451 17796 17463 17799
rect 17862 17796 17868 17808
rect 17451 17768 17868 17796
rect 17451 17765 17463 17768
rect 17405 17759 17463 17765
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1486 17728 1492 17740
rect 1443 17700 1492 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1486 17688 1492 17700
rect 1544 17728 1550 17740
rect 1762 17728 1768 17740
rect 1544 17700 1768 17728
rect 1544 17688 1550 17700
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 2682 17728 2688 17740
rect 2643 17700 2688 17728
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4338 17728 4344 17740
rect 4111 17700 4344 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17129 17731 17187 17737
rect 17129 17728 17141 17731
rect 16908 17700 17141 17728
rect 16908 17688 16914 17700
rect 17129 17697 17141 17700
rect 17175 17697 17187 17731
rect 17129 17691 17187 17697
rect 21085 17731 21143 17737
rect 21085 17697 21097 17731
rect 21131 17728 21143 17731
rect 21818 17728 21824 17740
rect 21131 17700 21824 17728
rect 21131 17697 21143 17700
rect 21085 17691 21143 17697
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 22373 17731 22431 17737
rect 22373 17697 22385 17731
rect 22419 17728 22431 17731
rect 22462 17728 22468 17740
rect 22419 17700 22468 17728
rect 22419 17697 22431 17700
rect 22373 17691 22431 17697
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17728 23535 17731
rect 23566 17728 23572 17740
rect 23523 17700 23572 17728
rect 23523 17697 23535 17700
rect 23477 17691 23535 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 2130 17620 2136 17672
rect 2188 17660 2194 17672
rect 2501 17663 2559 17669
rect 2501 17660 2513 17663
rect 2188 17632 2513 17660
rect 2188 17620 2194 17632
rect 2501 17629 2513 17632
rect 2547 17629 2559 17663
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 2501 17623 2559 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2133 17527 2191 17533
rect 2133 17524 2145 17527
rect 2096 17496 2145 17524
rect 2096 17484 2102 17496
rect 2133 17493 2145 17496
rect 2179 17524 2191 17527
rect 2222 17524 2228 17536
rect 2179 17496 2228 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 3329 17527 3387 17533
rect 3329 17493 3341 17527
rect 3375 17524 3387 17527
rect 3418 17524 3424 17536
rect 3375 17496 3424 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 3602 17524 3608 17536
rect 3563 17496 3608 17524
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 22557 17527 22615 17533
rect 22557 17493 22569 17527
rect 22603 17524 22615 17527
rect 23474 17524 23480 17536
rect 22603 17496 23480 17524
rect 22603 17493 22615 17496
rect 22557 17487 22615 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 23658 17524 23664 17536
rect 23619 17496 23664 17524
rect 23658 17484 23664 17496
rect 23716 17484 23722 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 23808 17292 24777 17320
rect 23808 17280 23814 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 24765 17283 24823 17289
rect 23842 17212 23848 17264
rect 23900 17252 23906 17264
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 23900 17224 24501 17252
rect 23900 17212 23906 17224
rect 24489 17221 24501 17224
rect 24535 17252 24547 17255
rect 24670 17252 24676 17264
rect 24535 17224 24676 17252
rect 24535 17221 24547 17224
rect 24489 17215 24547 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 2038 17184 2044 17196
rect 1999 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2188 17156 2233 17184
rect 2188 17144 2194 17156
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3329 17187 3387 17193
rect 3329 17184 3341 17187
rect 3016 17156 3341 17184
rect 3016 17144 3022 17156
rect 3329 17153 3341 17156
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 13354 17144 13360 17196
rect 13412 17184 13418 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13412 17156 13553 17184
rect 13412 17144 13418 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 13541 17147 13599 17153
rect 20088 17156 21557 17184
rect 3142 17116 3148 17128
rect 3055 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17116 3206 17128
rect 3602 17116 3608 17128
rect 3200 17088 3608 17116
rect 3200 17076 3206 17088
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 4433 17119 4491 17125
rect 4433 17085 4445 17119
rect 4479 17116 4491 17119
rect 4798 17116 4804 17128
rect 4479 17088 4804 17116
rect 4479 17085 4491 17088
rect 4433 17079 4491 17085
rect 4798 17076 4804 17088
rect 4856 17116 4862 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4856 17088 4997 17116
rect 4856 17076 4862 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13136 17088 13461 17116
rect 13136 17076 13142 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 12805 17051 12863 17057
rect 2832 17020 2877 17048
rect 2832 17008 2838 17020
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13262 17048 13268 17060
rect 12851 17020 13268 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13262 17008 13268 17020
rect 13320 17048 13326 17060
rect 13357 17051 13415 17057
rect 13357 17048 13369 17051
rect 13320 17020 13369 17048
rect 13320 17008 13326 17020
rect 13357 17017 13369 17020
rect 13403 17017 13415 17051
rect 13357 17011 13415 17017
rect 18414 17008 18420 17060
rect 18472 17048 18478 17060
rect 20088 17057 20116 17156
rect 21545 17153 21557 17156
rect 21591 17184 21603 17187
rect 22002 17184 22008 17196
rect 21591 17156 22008 17184
rect 21591 17153 21603 17156
rect 21545 17147 21603 17153
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21361 17119 21419 17125
rect 21361 17116 21373 17119
rect 20772 17088 21373 17116
rect 20772 17076 20778 17088
rect 21361 17085 21373 17088
rect 21407 17085 21419 17119
rect 21361 17079 21419 17085
rect 24486 17076 24492 17128
rect 24544 17116 24550 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24544 17088 24593 17116
rect 24544 17076 24550 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 20073 17051 20131 17057
rect 20073 17048 20085 17051
rect 18472 17020 20085 17048
rect 18472 17008 18478 17020
rect 20073 17017 20085 17020
rect 20119 17017 20131 17051
rect 20073 17011 20131 17017
rect 20533 17051 20591 17057
rect 20533 17017 20545 17051
rect 20579 17048 20591 17051
rect 21453 17051 21511 17057
rect 21453 17048 21465 17051
rect 20579 17020 21465 17048
rect 20579 17017 20591 17020
rect 20533 17011 20591 17017
rect 21453 17017 21465 17020
rect 21499 17048 21511 17051
rect 22278 17048 22284 17060
rect 21499 17020 22284 17048
rect 21499 17017 21511 17020
rect 21453 17011 21511 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22462 17048 22468 17060
rect 22423 17020 22468 17048
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 23566 17008 23572 17060
rect 23624 17048 23630 17060
rect 23937 17051 23995 17057
rect 23937 17048 23949 17051
rect 23624 17020 23949 17048
rect 23624 17008 23630 17020
rect 23937 17017 23949 17020
rect 23983 17048 23995 17051
rect 24762 17048 24768 17060
rect 23983 17020 24768 17048
rect 23983 17017 23995 17020
rect 23937 17011 23995 17017
rect 24762 17008 24768 17020
rect 24820 17008 24826 17060
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1728 16952 1961 16980
rect 1728 16940 1734 16952
rect 1949 16949 1961 16952
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4338 16980 4344 16992
rect 4203 16952 4344 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4614 16980 4620 16992
rect 4575 16952 4620 16980
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 12158 16980 12164 16992
rect 12119 16952 12164 16980
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12952 16952 13001 16980
rect 12952 16940 12958 16952
rect 12989 16949 13001 16952
rect 13035 16949 13047 16983
rect 12989 16943 13047 16949
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 16908 16952 17141 16980
rect 16908 16940 16914 16952
rect 17129 16949 17141 16952
rect 17175 16949 17187 16983
rect 18782 16980 18788 16992
rect 18743 16952 18788 16980
rect 17129 16943 17187 16949
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 20809 16983 20867 16989
rect 20809 16980 20821 16983
rect 20772 16952 20821 16980
rect 20772 16940 20778 16952
rect 20809 16949 20821 16952
rect 20855 16949 20867 16983
rect 20990 16980 20996 16992
rect 20951 16952 20996 16980
rect 20809 16943 20867 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21876 16952 22017 16980
rect 21876 16940 21882 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 22554 16980 22560 16992
rect 22515 16952 22560 16980
rect 22005 16943 22063 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 1636 16748 3617 16776
rect 1636 16736 1642 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 3605 16739 3663 16745
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 5353 16779 5411 16785
rect 5353 16776 5365 16779
rect 4120 16748 5365 16776
rect 4120 16736 4126 16748
rect 5353 16745 5365 16748
rect 5399 16745 5411 16779
rect 5353 16739 5411 16745
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12308 16748 13093 16776
rect 12308 16736 12314 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 18414 16776 18420 16788
rect 18371 16748 18420 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16776 19947 16779
rect 19978 16776 19984 16788
rect 19935 16748 19984 16776
rect 19935 16745 19947 16748
rect 19889 16739 19947 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20901 16779 20959 16785
rect 20901 16745 20913 16779
rect 20947 16776 20959 16779
rect 21910 16776 21916 16788
rect 20947 16748 21916 16776
rect 20947 16745 20959 16748
rect 20901 16739 20959 16745
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 23934 16776 23940 16788
rect 23799 16748 23940 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 25498 16776 25504 16788
rect 25459 16748 25504 16776
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 1857 16711 1915 16717
rect 1857 16677 1869 16711
rect 1903 16708 1915 16711
rect 17402 16708 17408 16720
rect 1903 16680 2728 16708
rect 1903 16677 1915 16680
rect 1857 16671 1915 16677
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 1949 16643 2007 16649
rect 1728 16612 1900 16640
rect 1728 16600 1734 16612
rect 1872 16504 1900 16612
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2498 16640 2504 16652
rect 1995 16612 2504 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 2700 16640 2728 16680
rect 16960 16680 17408 16708
rect 2774 16640 2780 16652
rect 2700 16612 2780 16640
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 4080 16572 4108 16603
rect 4246 16600 4252 16652
rect 4304 16600 4310 16652
rect 4614 16640 4620 16652
rect 4575 16612 4620 16640
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16640 5227 16643
rect 5442 16640 5448 16652
rect 5215 16612 5448 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16640 13231 16643
rect 13446 16640 13452 16652
rect 13219 16612 13452 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 16960 16649 16988 16680
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 21361 16711 21419 16717
rect 21361 16677 21373 16711
rect 21407 16708 21419 16711
rect 21450 16708 21456 16720
rect 21407 16680 21456 16708
rect 21407 16677 21419 16680
rect 21361 16671 21419 16677
rect 21450 16668 21456 16680
rect 21508 16668 21514 16720
rect 22830 16708 22836 16720
rect 22791 16680 22836 16708
rect 22830 16668 22836 16680
rect 22888 16668 22894 16720
rect 24210 16668 24216 16720
rect 24268 16708 24274 16720
rect 24305 16711 24363 16717
rect 24305 16708 24317 16711
rect 24268 16680 24317 16708
rect 24268 16668 24274 16680
rect 24305 16677 24317 16680
rect 24351 16677 24363 16711
rect 24305 16671 24363 16677
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14240 16612 14473 16640
rect 14240 16600 14246 16612
rect 14461 16609 14473 16612
rect 14507 16640 14519 16643
rect 14921 16643 14979 16649
rect 14921 16640 14933 16643
rect 14507 16612 14933 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 14921 16609 14933 16612
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17201 16643 17259 16649
rect 17201 16640 17213 16643
rect 17092 16612 17213 16640
rect 17092 16600 17098 16612
rect 17201 16609 17213 16612
rect 17247 16609 17259 16643
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 17201 16603 17259 16609
rect 19260 16612 19533 16640
rect 4154 16572 4160 16584
rect 4080 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1872 16476 2513 16504
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2866 16504 2872 16516
rect 2827 16476 2872 16504
rect 2501 16467 2559 16473
rect 2866 16464 2872 16476
rect 2924 16504 2930 16516
rect 4264 16513 4292 16600
rect 13354 16572 13360 16584
rect 13315 16544 13360 16572
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 19260 16572 19288 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19702 16640 19708 16652
rect 19663 16612 19708 16640
rect 19521 16603 19579 16609
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20640 16612 21281 16640
rect 18656 16544 19288 16572
rect 18656 16532 18662 16544
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 20640 16572 20668 16612
rect 21269 16609 21281 16612
rect 21315 16640 21327 16643
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 21315 16612 22293 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 22922 16640 22928 16652
rect 22883 16612 22928 16640
rect 22281 16603 22339 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16640 24087 16643
rect 24670 16640 24676 16652
rect 24075 16612 24676 16640
rect 24075 16609 24087 16612
rect 24029 16603 24087 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25774 16640 25780 16652
rect 25363 16612 25780 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 20128 16544 20668 16572
rect 21453 16575 21511 16581
rect 20128 16532 20134 16544
rect 21453 16541 21465 16575
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 3237 16507 3295 16513
rect 3237 16504 3249 16507
rect 2924 16476 3249 16504
rect 2924 16464 2930 16476
rect 3237 16473 3249 16476
rect 3283 16473 3295 16507
rect 3237 16467 3295 16473
rect 4249 16507 4307 16513
rect 4249 16473 4261 16507
rect 4295 16473 4307 16507
rect 4249 16467 4307 16473
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21468 16504 21496 16535
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 22738 16572 22744 16584
rect 22060 16544 22744 16572
rect 22060 16532 22066 16544
rect 22738 16532 22744 16544
rect 22796 16572 22802 16584
rect 23017 16575 23075 16581
rect 23017 16572 23029 16575
rect 22796 16544 23029 16572
rect 22796 16532 22802 16544
rect 23017 16541 23029 16544
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 21324 16476 21496 16504
rect 21324 16464 21330 16476
rect 1489 16439 1547 16445
rect 1489 16405 1501 16439
rect 1535 16436 1547 16439
rect 2130 16436 2136 16448
rect 1535 16408 2136 16436
rect 1535 16405 1547 16408
rect 1489 16399 1547 16405
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 5077 16439 5135 16445
rect 5077 16405 5089 16439
rect 5123 16436 5135 16439
rect 5534 16436 5540 16448
rect 5123 16408 5540 16436
rect 5123 16405 5135 16408
rect 5077 16399 5135 16405
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 12066 16436 12072 16448
rect 10836 16408 12072 16436
rect 10836 16396 10842 16408
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12526 16436 12532 16448
rect 12487 16408 12532 16436
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 12710 16436 12716 16448
rect 12671 16408 12716 16436
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 14090 16436 14096 16448
rect 14051 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 20346 16436 20352 16448
rect 20307 16408 20352 16436
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20496 16408 20637 16436
rect 20496 16396 20502 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 22002 16436 22008 16448
rect 21963 16408 22008 16436
rect 20625 16399 20683 16405
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 22462 16436 22468 16448
rect 22423 16408 22468 16436
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 2498 16232 2504 16244
rect 1452 16204 2504 16232
rect 1452 16192 1458 16204
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5592 16204 5733 16232
rect 5592 16192 5598 16204
rect 5721 16201 5733 16204
rect 5767 16232 5779 16235
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 5767 16204 6101 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6089 16201 6101 16204
rect 6135 16232 6147 16235
rect 6362 16232 6368 16244
rect 6135 16204 6368 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 20070 16232 20076 16244
rect 20031 16204 20076 16232
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 22649 16235 22707 16241
rect 22649 16201 22661 16235
rect 22695 16232 22707 16235
rect 22922 16232 22928 16244
rect 22695 16204 22928 16232
rect 22695 16201 22707 16204
rect 22649 16195 22707 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 25406 16232 25412 16244
rect 25367 16204 25412 16232
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 2961 16167 3019 16173
rect 2961 16133 2973 16167
rect 3007 16164 3019 16167
rect 3234 16164 3240 16176
rect 3007 16136 3240 16164
rect 3007 16133 3019 16136
rect 2961 16127 3019 16133
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 22060 16136 22140 16164
rect 22060 16124 22066 16136
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 1949 16099 2007 16105
rect 1949 16096 1961 16099
rect 1636 16068 1961 16096
rect 1636 16056 1642 16068
rect 1949 16065 1961 16068
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2498 16096 2504 16108
rect 2179 16068 2504 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2866 16056 2872 16108
rect 2924 16096 2930 16108
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 2924 16068 3617 16096
rect 2924 16056 2930 16068
rect 3605 16065 3617 16068
rect 3651 16065 3663 16099
rect 4798 16096 4804 16108
rect 4759 16068 4804 16096
rect 3605 16059 3663 16065
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 12986 16096 12992 16108
rect 12584 16068 12992 16096
rect 12584 16056 12590 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 20346 16056 20352 16108
rect 20404 16096 20410 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20404 16068 20637 16096
rect 20404 16056 20410 16068
rect 20625 16065 20637 16068
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 21358 16056 21364 16108
rect 21416 16096 21422 16108
rect 22112 16096 22140 16136
rect 22738 16124 22744 16176
rect 22796 16164 22802 16176
rect 22796 16136 24256 16164
rect 22796 16124 22802 16136
rect 22189 16099 22247 16105
rect 22189 16096 22201 16099
rect 21416 16068 22201 16096
rect 21416 16056 21422 16068
rect 22189 16065 22201 16068
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 23934 16056 23940 16108
rect 23992 16096 23998 16108
rect 24118 16096 24124 16108
rect 23992 16068 24124 16096
rect 23992 16056 23998 16068
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 24228 16105 24256 16136
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16096 24271 16099
rect 24673 16099 24731 16105
rect 24673 16096 24685 16099
rect 24259 16068 24685 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 24673 16065 24685 16068
rect 24719 16065 24731 16099
rect 24673 16059 24731 16065
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3016 16000 3433 16028
rect 3016 15988 3022 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 4154 16028 4160 16040
rect 4115 16000 4160 16028
rect 3421 15991 3479 15997
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4540 16000 4629 16028
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15960 1915 15963
rect 1903 15932 3096 15960
rect 1903 15929 1915 15932
rect 1857 15923 1915 15929
rect 3068 15904 3096 15932
rect 4540 15904 4568 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 12805 16031 12863 16037
rect 12805 16028 12817 16031
rect 12124 16000 12817 16028
rect 12124 15988 12130 16000
rect 12805 15997 12817 16000
rect 12851 15997 12863 16031
rect 14461 16031 14519 16037
rect 14461 16028 14473 16031
rect 12805 15991 12863 15997
rect 13924 16000 14473 16028
rect 12158 15960 12164 15972
rect 11808 15932 12164 15960
rect 1489 15895 1547 15901
rect 1489 15861 1501 15895
rect 1535 15892 1547 15895
rect 1762 15892 1768 15904
rect 1535 15864 1768 15892
rect 1535 15861 1547 15864
rect 1489 15855 1547 15861
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 3050 15892 3056 15904
rect 3011 15864 3056 15892
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 3326 15852 3332 15904
rect 3384 15892 3390 15904
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 3384 15864 3525 15892
rect 3384 15852 3390 15864
rect 3513 15861 3525 15864
rect 3559 15861 3571 15895
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 3513 15855 3571 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5442 15892 5448 15904
rect 5403 15864 5448 15892
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 11808 15901 11836 15932
rect 12158 15920 12164 15932
rect 12216 15960 12222 15972
rect 13354 15960 13360 15972
rect 12216 15932 13360 15960
rect 12216 15920 12222 15932
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 13924 15904 13952 16000
rect 14461 15997 14473 16000
rect 14507 15997 14519 16031
rect 20438 16028 20444 16040
rect 20399 16000 20444 16028
rect 14461 15991 14519 15997
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 16028 21235 16031
rect 22002 16028 22008 16040
rect 21223 16000 22008 16028
rect 21223 15997 21235 16000
rect 21177 15991 21235 15997
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 22888 16000 23121 16028
rect 22888 15988 22894 16000
rect 23109 15997 23121 16000
rect 23155 16028 23167 16031
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 23155 16000 24164 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 24136 15972 24164 16000
rect 25056 16000 25237 16028
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14369 15963 14427 15969
rect 14369 15960 14381 15963
rect 14148 15932 14381 15960
rect 14148 15920 14154 15932
rect 14369 15929 14381 15932
rect 14415 15929 14427 15963
rect 14369 15923 14427 15929
rect 14826 15920 14832 15972
rect 14884 15960 14890 15972
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 14884 15932 15577 15960
rect 14884 15920 14890 15932
rect 15565 15929 15577 15932
rect 15611 15929 15623 15963
rect 15565 15923 15623 15929
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 19702 15960 19708 15972
rect 18012 15932 19708 15960
rect 18012 15920 18018 15932
rect 19702 15920 19708 15932
rect 19760 15920 19766 15972
rect 21545 15963 21603 15969
rect 21545 15929 21557 15963
rect 21591 15960 21603 15963
rect 21726 15960 21732 15972
rect 21591 15932 21732 15960
rect 21591 15929 21603 15932
rect 21545 15923 21603 15929
rect 21726 15920 21732 15932
rect 21784 15960 21790 15972
rect 22097 15963 22155 15969
rect 22097 15960 22109 15963
rect 21784 15932 22109 15960
rect 21784 15920 21790 15932
rect 22097 15929 22109 15932
rect 22143 15929 22155 15963
rect 23474 15960 23480 15972
rect 23387 15932 23480 15960
rect 22097 15923 22155 15929
rect 23474 15920 23480 15932
rect 23532 15960 23538 15972
rect 24029 15963 24087 15969
rect 24029 15960 24041 15963
rect 23532 15932 24041 15960
rect 23532 15920 23538 15932
rect 24029 15929 24041 15932
rect 24075 15929 24087 15963
rect 24029 15923 24087 15929
rect 24118 15920 24124 15972
rect 24176 15920 24182 15972
rect 25056 15904 25084 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11756 15864 11805 15892
rect 11756 15852 11762 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 12250 15892 12256 15904
rect 12211 15864 12256 15892
rect 11793 15855 11851 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12492 15864 12537 15892
rect 12492 15852 12498 15864
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12860 15864 12909 15892
rect 12860 15852 12866 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 13446 15892 13452 15904
rect 13407 15864 13452 15892
rect 12897 15855 12955 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 13906 15892 13912 15904
rect 13867 15864 13912 15892
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14274 15892 14280 15904
rect 14047 15864 14280 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15930 15892 15936 15904
rect 15427 15864 15936 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 16577 15895 16635 15901
rect 16577 15892 16589 15895
rect 16356 15864 16589 15892
rect 16356 15852 16362 15864
rect 16577 15861 16589 15864
rect 16623 15861 16635 15895
rect 17402 15892 17408 15904
rect 17363 15864 17408 15892
rect 16577 15855 16635 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 18046 15892 18052 15904
rect 18007 15864 18052 15892
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 19061 15895 19119 15901
rect 19061 15892 19073 15895
rect 18748 15864 19073 15892
rect 18748 15852 18754 15864
rect 19061 15861 19073 15864
rect 19107 15861 19119 15895
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 19061 15855 19119 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 21634 15892 21640 15904
rect 21595 15864 21640 15892
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 23566 15852 23572 15904
rect 23624 15892 23630 15904
rect 23661 15895 23719 15901
rect 23661 15892 23673 15895
rect 23624 15864 23673 15892
rect 23624 15852 23630 15864
rect 23661 15861 23673 15864
rect 23707 15861 23719 15895
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 23661 15855 23719 15861
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 25774 15892 25780 15904
rect 25735 15864 25780 15892
rect 25774 15852 25780 15864
rect 25832 15852 25838 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 2832 15660 2877 15688
rect 2832 15648 2838 15660
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3108 15660 3801 15688
rect 3108 15648 3114 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 3878 15648 3884 15700
rect 3936 15688 3942 15700
rect 5166 15688 5172 15700
rect 3936 15660 5172 15688
rect 3936 15648 3942 15660
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 6362 15688 6368 15700
rect 6323 15660 6368 15688
rect 6362 15648 6368 15660
rect 6420 15688 6426 15700
rect 6733 15691 6791 15697
rect 6733 15688 6745 15691
rect 6420 15660 6745 15688
rect 6420 15648 6426 15660
rect 6733 15657 6745 15660
rect 6779 15688 6791 15691
rect 6822 15688 6828 15700
rect 6779 15660 6828 15688
rect 6779 15657 6791 15660
rect 6733 15651 6791 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7098 15688 7104 15700
rect 7059 15660 7104 15688
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13412 15660 14197 15688
rect 13412 15648 13418 15660
rect 14185 15657 14197 15660
rect 14231 15688 14243 15691
rect 14550 15688 14556 15700
rect 14231 15660 14556 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 20438 15688 20444 15700
rect 19291 15660 20444 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 22462 15648 22468 15700
rect 22520 15688 22526 15700
rect 23109 15691 23167 15697
rect 23109 15688 23121 15691
rect 22520 15660 23121 15688
rect 22520 15648 22526 15660
rect 23109 15657 23121 15660
rect 23155 15688 23167 15691
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 23155 15660 23673 15688
rect 23155 15657 23167 15660
rect 23109 15651 23167 15657
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 2041 15623 2099 15629
rect 2041 15589 2053 15623
rect 2087 15620 2099 15623
rect 2314 15620 2320 15632
rect 2087 15592 2320 15620
rect 2087 15589 2099 15592
rect 2041 15583 2099 15589
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 5905 15623 5963 15629
rect 5905 15620 5917 15623
rect 5500 15592 5917 15620
rect 5500 15580 5506 15592
rect 5905 15589 5917 15592
rect 5951 15589 5963 15623
rect 5905 15583 5963 15589
rect 11425 15623 11483 15629
rect 11425 15589 11437 15623
rect 11471 15620 11483 15623
rect 11471 15592 11928 15620
rect 11471 15589 11483 15592
rect 11425 15583 11483 15589
rect 2130 15512 2136 15564
rect 2188 15552 2194 15564
rect 3142 15552 3148 15564
rect 2188 15524 3148 15552
rect 2188 15512 2194 15524
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 3752 15524 4445 15552
rect 3752 15512 3758 15524
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 5994 15552 6000 15564
rect 5675 15524 6000 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15552 6975 15555
rect 7650 15552 7656 15564
rect 6963 15524 7656 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 11790 15561 11796 15564
rect 11784 15552 11796 15561
rect 11751 15524 11796 15552
rect 11784 15515 11796 15524
rect 11790 15512 11796 15515
rect 11848 15512 11854 15564
rect 11900 15552 11928 15592
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13725 15623 13783 15629
rect 13725 15620 13737 15623
rect 12492 15592 13737 15620
rect 12492 15580 12498 15592
rect 13725 15589 13737 15592
rect 13771 15589 13783 15623
rect 13725 15583 13783 15589
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 18012 15592 18061 15620
rect 18012 15580 18018 15592
rect 18049 15589 18061 15592
rect 18095 15589 18107 15623
rect 22097 15623 22155 15629
rect 18049 15583 18107 15589
rect 19444 15592 19932 15620
rect 13630 15552 13636 15564
rect 11900 15524 13636 15552
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2225 15487 2283 15493
rect 2225 15484 2237 15487
rect 2004 15456 2237 15484
rect 2004 15444 2010 15456
rect 2225 15453 2237 15456
rect 2271 15484 2283 15487
rect 2498 15484 2504 15496
rect 2271 15456 2504 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4304 15456 4537 15484
rect 4304 15444 4310 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 4798 15484 4804 15496
rect 4755 15456 4804 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 10042 15444 10048 15496
rect 10100 15484 10106 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 10100 15456 10517 15484
rect 10100 15444 10106 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 11514 15484 11520 15496
rect 11475 15456 11520 15484
rect 10505 15447 10563 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 15010 15484 15016 15496
rect 14971 15456 15016 15484
rect 15010 15444 15016 15456
rect 15068 15484 15074 15496
rect 15672 15484 15700 15515
rect 15068 15456 15700 15484
rect 15068 15444 15074 15456
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 15804 15456 15849 15484
rect 15804 15444 15810 15456
rect 15930 15444 15936 15496
rect 15988 15484 15994 15496
rect 15988 15456 16436 15484
rect 15988 15444 15994 15456
rect 1673 15419 1731 15425
rect 1673 15385 1685 15419
rect 1719 15416 1731 15419
rect 1762 15416 1768 15428
rect 1719 15388 1768 15416
rect 1719 15385 1731 15388
rect 1673 15379 1731 15385
rect 1762 15376 1768 15388
rect 1820 15416 1826 15428
rect 3421 15419 3479 15425
rect 3421 15416 3433 15419
rect 1820 15388 3433 15416
rect 1820 15376 1826 15388
rect 3421 15385 3433 15388
rect 3467 15385 3479 15419
rect 5534 15416 5540 15428
rect 5495 15388 5540 15416
rect 3421 15379 3479 15385
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13265 15419 13323 15425
rect 13265 15416 13277 15419
rect 12860 15388 13277 15416
rect 12860 15376 12866 15388
rect 13265 15385 13277 15388
rect 13311 15416 13323 15419
rect 13722 15416 13728 15428
rect 13311 15388 13728 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13722 15376 13728 15388
rect 13780 15376 13786 15428
rect 16408 15360 16436 15456
rect 17494 15444 17500 15496
rect 17552 15484 17558 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 17552 15456 18153 15484
rect 17552 15444 17558 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18288 15456 18337 15484
rect 18288 15444 18294 15456
rect 18325 15453 18337 15456
rect 18371 15484 18383 15487
rect 19444 15484 19472 15592
rect 19610 15552 19616 15564
rect 19571 15524 19616 15552
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 18371 15456 19472 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19904 15493 19932 15592
rect 22097 15589 22109 15623
rect 22143 15620 22155 15623
rect 22186 15620 22192 15632
rect 22143 15592 22192 15620
rect 22143 15589 22155 15592
rect 22097 15583 22155 15589
rect 22186 15580 22192 15592
rect 22244 15620 22250 15632
rect 22554 15620 22560 15632
rect 22244 15592 22560 15620
rect 22244 15580 22250 15592
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 22738 15620 22744 15632
rect 22699 15592 22744 15620
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 24670 15620 24676 15632
rect 24631 15592 24676 15620
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 24946 15580 24952 15632
rect 25004 15620 25010 15632
rect 25133 15623 25191 15629
rect 25133 15620 25145 15623
rect 25004 15592 25145 15620
rect 25004 15580 25010 15592
rect 25133 15589 25145 15592
rect 25179 15589 25191 15623
rect 25133 15583 25191 15589
rect 23658 15512 23664 15564
rect 23716 15552 23722 15564
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 23716 15524 24409 15552
rect 23716 15512 23722 15524
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 24857 15555 24915 15561
rect 24857 15521 24869 15555
rect 24903 15552 24915 15555
rect 25038 15552 25044 15564
rect 24903 15524 25044 15552
rect 24903 15521 24915 15524
rect 24857 15515 24915 15521
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19576 15456 19717 15484
rect 19576 15444 19582 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20438 15484 20444 15496
rect 19935 15456 20444 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 22152 15456 22201 15484
rect 22152 15444 22158 15456
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 22370 15484 22376 15496
rect 22331 15456 22376 15484
rect 22189 15447 22247 15453
rect 22370 15444 22376 15456
rect 22428 15444 22434 15496
rect 23566 15444 23572 15496
rect 23624 15484 23630 15496
rect 23753 15487 23811 15493
rect 23753 15484 23765 15487
rect 23624 15456 23765 15484
rect 23624 15444 23630 15456
rect 23753 15453 23765 15456
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 23842 15444 23848 15496
rect 23900 15484 23906 15496
rect 23900 15456 23945 15484
rect 23900 15444 23906 15456
rect 17681 15419 17739 15425
rect 17681 15385 17693 15419
rect 17727 15416 17739 15419
rect 20530 15416 20536 15428
rect 17727 15388 20536 15416
rect 17727 15385 17739 15388
rect 17681 15379 17739 15385
rect 20530 15376 20536 15388
rect 20588 15416 20594 15428
rect 20625 15419 20683 15425
rect 20625 15416 20637 15419
rect 20588 15388 20637 15416
rect 20588 15376 20594 15388
rect 20625 15385 20637 15388
rect 20671 15385 20683 15419
rect 20625 15379 20683 15385
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 2314 15348 2320 15360
rect 1360 15320 2320 15348
rect 1360 15308 1366 15320
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 2498 15308 2504 15360
rect 2556 15348 2562 15360
rect 2774 15348 2780 15360
rect 2556 15320 2780 15348
rect 2556 15308 2562 15320
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 2958 15308 2964 15360
rect 3016 15348 3022 15360
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 3016 15320 3065 15348
rect 3016 15308 3022 15320
rect 3053 15317 3065 15320
rect 3099 15317 3111 15351
rect 4062 15348 4068 15360
rect 4023 15320 4068 15348
rect 3053 15311 3111 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 5040 15320 5089 15348
rect 5040 15308 5046 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 7561 15351 7619 15357
rect 7561 15317 7573 15351
rect 7607 15348 7619 15351
rect 8110 15348 8116 15360
rect 7607 15320 8116 15348
rect 7607 15317 7619 15320
rect 7561 15311 7619 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12897 15351 12955 15357
rect 12897 15317 12909 15351
rect 12943 15348 12955 15351
rect 13170 15348 13176 15360
rect 12943 15320 13176 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 14642 15348 14648 15360
rect 14603 15320 14648 15348
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 15286 15348 15292 15360
rect 15247 15320 15292 15348
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 16390 15348 16396 15360
rect 16351 15320 16396 15348
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 16761 15351 16819 15357
rect 16761 15348 16773 15351
rect 16632 15320 16773 15348
rect 16632 15308 16638 15320
rect 16761 15317 16773 15320
rect 16807 15348 16819 15351
rect 17129 15351 17187 15357
rect 17129 15348 17141 15351
rect 16807 15320 17141 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 17129 15317 17141 15320
rect 17175 15348 17187 15351
rect 17402 15348 17408 15360
rect 17175 15320 17408 15348
rect 17175 15317 17187 15320
rect 17129 15311 17187 15317
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 19061 15351 19119 15357
rect 19061 15348 19073 15351
rect 18932 15320 19073 15348
rect 18932 15308 18938 15320
rect 19061 15317 19073 15320
rect 19107 15317 19119 15351
rect 19061 15311 19119 15317
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15348 20407 15351
rect 20438 15348 20444 15360
rect 20395 15320 20444 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 21177 15351 21235 15357
rect 21177 15317 21189 15351
rect 21223 15348 21235 15351
rect 21266 15348 21272 15360
rect 21223 15320 21272 15348
rect 21223 15317 21235 15320
rect 21177 15311 21235 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 21726 15348 21732 15360
rect 21687 15320 21732 15348
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 23293 15351 23351 15357
rect 23293 15348 23305 15351
rect 22520 15320 23305 15348
rect 22520 15308 22526 15320
rect 23293 15317 23305 15320
rect 23339 15317 23351 15351
rect 23293 15311 23351 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2047 15116 2912 15144
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 2047 15017 2075 15116
rect 2884 15085 2912 15116
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 7926 15144 7932 15156
rect 6880 15116 7932 15144
rect 6880 15104 6886 15116
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 10192 15116 10517 15144
rect 10192 15104 10198 15116
rect 10505 15113 10517 15116
rect 10551 15144 10563 15147
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 10551 15116 10609 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10597 15107 10655 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 13872 15116 14657 15144
rect 13872 15104 13878 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 17773 15147 17831 15153
rect 17773 15113 17785 15147
rect 17819 15144 17831 15147
rect 17862 15144 17868 15156
rect 17819 15116 17868 15144
rect 17819 15113 17831 15116
rect 17773 15107 17831 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 21269 15147 21327 15153
rect 21269 15113 21281 15147
rect 21315 15144 21327 15147
rect 21358 15144 21364 15156
rect 21315 15116 21364 15144
rect 21315 15113 21327 15116
rect 21269 15107 21327 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 22186 15144 22192 15156
rect 22147 15116 22192 15144
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22428 15116 23029 15144
rect 22428 15104 22434 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 2869 15079 2927 15085
rect 2869 15045 2881 15079
rect 2915 15076 2927 15079
rect 11609 15079 11667 15085
rect 2915 15048 3648 15076
rect 2915 15045 2927 15048
rect 2869 15039 2927 15045
rect 3620 15020 3648 15048
rect 11609 15045 11621 15079
rect 11655 15076 11667 15079
rect 12434 15076 12440 15088
rect 11655 15048 12440 15076
rect 11655 15045 11667 15048
rect 11609 15039 11667 15045
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 13630 15036 13636 15088
rect 13688 15076 13694 15088
rect 14182 15076 14188 15088
rect 13688 15048 14188 15076
rect 13688 15036 13694 15048
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 18325 15079 18383 15085
rect 18325 15045 18337 15079
rect 18371 15076 18383 15079
rect 19334 15076 19340 15088
rect 18371 15048 19340 15076
rect 18371 15045 18383 15048
rect 18325 15039 18383 15045
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 24762 15036 24768 15088
rect 24820 15076 24826 15088
rect 24820 15048 25452 15076
rect 24820 15036 24826 15048
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 3602 15008 3608 15020
rect 3563 14980 3608 15008
rect 2041 14971 2099 14977
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 4798 15008 4804 15020
rect 4295 14980 4804 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4798 14968 4804 14980
rect 4856 15008 4862 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4856 14980 5089 15008
rect 4856 14968 4862 14980
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 6972 14980 7021 15008
rect 6972 14968 6978 14980
rect 7009 14977 7021 14980
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 11112 14980 11345 15008
rect 11112 14968 11118 14980
rect 11333 14977 11345 14980
rect 11379 15008 11391 15011
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11379 14980 12173 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 12161 14977 12173 14980
rect 12207 15008 12219 15011
rect 12207 14980 12572 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 4062 14940 4068 14952
rect 3467 14912 4068 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4982 14940 4988 14952
rect 4396 14912 4988 14940
rect 4396 14900 4402 14912
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 5994 14940 6000 14952
rect 5767 14912 6000 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 6822 14940 6828 14952
rect 6687 14912 6828 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 8018 14900 8024 14952
rect 8076 14940 8082 14952
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 8076 14912 8125 14940
rect 8076 14900 8082 14912
rect 8113 14909 8125 14912
rect 8159 14940 8171 14943
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8159 14912 8677 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10367 14912 11161 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 11149 14909 11161 14912
rect 11195 14940 11207 14943
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11195 14912 11621 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 12434 14940 12440 14952
rect 12395 14912 12440 14940
rect 11609 14903 11667 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12544 14940 12572 14980
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14792 14980 15209 15008
rect 14792 14968 14798 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 16758 15008 16764 15020
rect 16719 14980 16764 15008
rect 15197 14971 15255 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 18874 15008 18880 15020
rect 18835 14980 18880 15008
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 15008 22615 15011
rect 23382 15008 23388 15020
rect 22603 14980 23388 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 23842 14968 23848 15020
rect 23900 15008 23906 15020
rect 25424 15017 25452 15048
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23900 14980 24225 15008
rect 23900 14968 23906 14980
rect 24213 14977 24225 14980
rect 24259 15008 24271 15011
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24259 14980 24685 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24673 14977 24685 14980
rect 24719 15008 24731 15011
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24719 14980 25053 15008
rect 24719 14977 24731 14980
rect 24673 14971 24731 14977
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 25409 15011 25467 15017
rect 25409 14977 25421 15011
rect 25455 14977 25467 15011
rect 25409 14971 25467 14977
rect 12704 14943 12762 14949
rect 12704 14940 12716 14943
rect 12544 14912 12716 14940
rect 12704 14909 12716 14912
rect 12750 14940 12762 14943
rect 13170 14940 13176 14952
rect 12750 14912 13176 14940
rect 12750 14909 12762 14912
rect 12704 14903 12762 14909
rect 13170 14900 13176 14912
rect 13228 14940 13234 14952
rect 14752 14940 14780 14968
rect 13228 14912 14780 14940
rect 13228 14900 13234 14912
rect 15838 14900 15844 14952
rect 15896 14940 15902 14952
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 15896 14912 16129 14940
rect 15896 14900 15902 14912
rect 16117 14909 16129 14912
rect 16163 14940 16175 14943
rect 16577 14943 16635 14949
rect 16577 14940 16589 14943
rect 16163 14912 16589 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16577 14909 16589 14912
rect 16623 14940 16635 14943
rect 16942 14940 16948 14952
rect 16623 14912 16948 14940
rect 16623 14909 16635 14912
rect 16577 14903 16635 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 18782 14940 18788 14952
rect 18739 14912 18788 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19536 14912 19901 14940
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 3375 14844 4568 14872
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 4540 14816 4568 14844
rect 4908 14844 6101 14872
rect 1397 14807 1455 14813
rect 1397 14773 1409 14807
rect 1443 14804 1455 14807
rect 2130 14804 2136 14816
rect 1443 14776 2136 14804
rect 1443 14773 1455 14776
rect 1397 14767 1455 14773
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 2406 14804 2412 14816
rect 2367 14776 2412 14804
rect 2406 14764 2412 14776
rect 2464 14764 2470 14816
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 2961 14807 3019 14813
rect 2961 14804 2973 14807
rect 2924 14776 2973 14804
rect 2924 14764 2930 14776
rect 2961 14773 2973 14776
rect 3007 14773 3019 14807
rect 2961 14767 3019 14773
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3936 14776 3985 14804
rect 3936 14764 3942 14776
rect 3973 14773 3985 14776
rect 4019 14804 4031 14807
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 4019 14776 4261 14804
rect 4019 14773 4031 14776
rect 3973 14767 4031 14773
rect 4249 14773 4261 14776
rect 4295 14804 4307 14807
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4295 14776 4353 14804
rect 4295 14773 4307 14776
rect 4249 14767 4307 14773
rect 4341 14773 4353 14776
rect 4387 14773 4399 14807
rect 4522 14804 4528 14816
rect 4483 14776 4528 14804
rect 4341 14767 4399 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 4908 14813 4936 14844
rect 6089 14841 6101 14844
rect 6135 14841 6147 14875
rect 6089 14835 6147 14841
rect 10505 14875 10563 14881
rect 10505 14841 10517 14875
rect 10551 14872 10563 14875
rect 11241 14875 11299 14881
rect 11241 14872 11253 14875
rect 10551 14844 11253 14872
rect 10551 14841 10563 14844
rect 10505 14835 10563 14841
rect 11241 14841 11253 14844
rect 11287 14841 11299 14875
rect 11241 14835 11299 14841
rect 12802 14832 12808 14884
rect 12860 14872 12866 14884
rect 14642 14872 14648 14884
rect 12860 14844 14648 14872
rect 12860 14832 12866 14844
rect 14642 14832 14648 14844
rect 14700 14872 14706 14884
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14700 14844 15117 14872
rect 14700 14832 14706 14844
rect 15105 14841 15117 14844
rect 15151 14841 15163 14875
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 15105 14835 15163 14841
rect 15672 14844 16681 14872
rect 15672 14816 15700 14844
rect 16669 14841 16681 14844
rect 16715 14841 16727 14875
rect 16669 14835 16727 14841
rect 18598 14832 18604 14884
rect 18656 14872 18662 14884
rect 19536 14872 19564 14912
rect 19889 14909 19901 14912
rect 19935 14940 19947 14943
rect 20530 14940 20536 14952
rect 19935 14912 20536 14940
rect 19935 14909 19947 14912
rect 19889 14903 19947 14909
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22278 14940 22284 14952
rect 21968 14912 22284 14940
rect 21968 14900 21974 14912
rect 22278 14900 22284 14912
rect 22336 14900 22342 14952
rect 23658 14900 23664 14952
rect 23716 14940 23722 14952
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23716 14912 24133 14940
rect 23716 14900 23722 14912
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 25222 14940 25228 14952
rect 25183 14912 25228 14940
rect 24121 14903 24179 14909
rect 25222 14900 25228 14912
rect 25280 14940 25286 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25280 14912 25973 14940
rect 25280 14900 25286 14912
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 18656 14844 19564 14872
rect 18656 14832 18662 14844
rect 19610 14832 19616 14884
rect 19668 14832 19674 14884
rect 20070 14832 20076 14884
rect 20128 14881 20134 14884
rect 20128 14875 20192 14881
rect 20128 14841 20146 14875
rect 20180 14841 20192 14875
rect 20128 14835 20192 14841
rect 20128 14832 20134 14835
rect 21542 14832 21548 14884
rect 21600 14872 21606 14884
rect 21729 14875 21787 14881
rect 21729 14872 21741 14875
rect 21600 14844 21741 14872
rect 21600 14832 21606 14844
rect 21729 14841 21741 14844
rect 21775 14872 21787 14875
rect 22094 14872 22100 14884
rect 21775 14844 22100 14872
rect 21775 14841 21787 14844
rect 21729 14835 21787 14841
rect 22094 14832 22100 14844
rect 22152 14832 22158 14884
rect 24029 14875 24087 14881
rect 24029 14872 24041 14875
rect 23492 14844 24041 14872
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4856 14776 4905 14804
rect 4856 14764 4862 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 7650 14804 7656 14816
rect 7611 14776 7656 14804
rect 4893 14767 4951 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 9214 14804 9220 14816
rect 9175 14776 9220 14804
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 13044 14776 13829 14804
rect 13044 14764 13050 14776
rect 13817 14773 13829 14776
rect 13863 14773 13875 14807
rect 13817 14767 13875 14773
rect 14553 14807 14611 14813
rect 14553 14773 14565 14807
rect 14599 14804 14611 14807
rect 15010 14804 15016 14816
rect 14599 14776 15016 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 18785 14807 18843 14813
rect 18785 14804 18797 14807
rect 18380 14776 18797 14804
rect 18380 14764 18386 14776
rect 18785 14773 18797 14776
rect 18831 14804 18843 14807
rect 18966 14804 18972 14816
rect 18831 14776 18972 14804
rect 18831 14773 18843 14776
rect 18785 14767 18843 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19426 14804 19432 14816
rect 19387 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19628 14804 19656 14832
rect 23492 14816 23520 14844
rect 24029 14841 24041 14844
rect 24075 14841 24087 14875
rect 24029 14835 24087 14841
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19628 14776 19809 14804
rect 19797 14773 19809 14776
rect 19843 14804 19855 14807
rect 20438 14804 20444 14816
rect 19843 14776 20444 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 23474 14804 23480 14816
rect 23435 14776 23480 14804
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 23658 14804 23664 14816
rect 23619 14776 23664 14804
rect 23658 14764 23664 14776
rect 23716 14764 23722 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2682 14600 2688 14612
rect 2455 14572 2688 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 3418 14600 3424 14612
rect 2915 14572 3424 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 4580 14572 5457 14600
rect 4580 14560 4586 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 7834 14600 7840 14612
rect 7795 14572 7840 14600
rect 5445 14563 5503 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7984 14572 8217 14600
rect 7984 14560 7990 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 11701 14603 11759 14609
rect 11701 14569 11713 14603
rect 11747 14600 11759 14603
rect 11790 14600 11796 14612
rect 11747 14572 11796 14600
rect 11747 14569 11759 14572
rect 11701 14563 11759 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 14734 14600 14740 14612
rect 14695 14572 14740 14600
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 17957 14603 18015 14609
rect 17957 14569 17969 14603
rect 18003 14600 18015 14603
rect 18230 14600 18236 14612
rect 18003 14572 18236 14600
rect 18003 14569 18015 14572
rect 17957 14563 18015 14569
rect 18230 14560 18236 14572
rect 18288 14560 18294 14612
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 20588 14572 20637 14600
rect 20588 14560 20594 14572
rect 20625 14569 20637 14572
rect 20671 14600 20683 14603
rect 20714 14600 20720 14612
rect 20671 14572 20720 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 22278 14560 22284 14612
rect 22336 14600 22342 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22336 14572 22845 14600
rect 22336 14560 22342 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 23293 14603 23351 14609
rect 23293 14569 23305 14603
rect 23339 14600 23351 14603
rect 23566 14600 23572 14612
rect 23339 14572 23572 14600
rect 23339 14569 23351 14572
rect 23293 14563 23351 14569
rect 23566 14560 23572 14572
rect 23624 14560 23630 14612
rect 4893 14535 4951 14541
rect 4893 14532 4905 14535
rect 4724 14504 4905 14532
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 2740 14436 2789 14464
rect 2740 14424 2746 14436
rect 2777 14433 2789 14436
rect 2823 14464 2835 14467
rect 4614 14464 4620 14476
rect 2823 14436 4620 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4724 14396 4752 14504
rect 4893 14501 4905 14504
rect 4939 14532 4951 14535
rect 5813 14535 5871 14541
rect 5813 14532 5825 14535
rect 4939 14504 5825 14532
rect 4939 14501 4951 14504
rect 4893 14495 4951 14501
rect 5813 14501 5825 14504
rect 5859 14501 5871 14535
rect 5813 14495 5871 14501
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14532 6607 14535
rect 6638 14532 6644 14544
rect 6595 14504 6644 14532
rect 6595 14501 6607 14504
rect 6549 14495 6607 14501
rect 6638 14492 6644 14504
rect 6696 14492 6702 14544
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 13234 14535 13292 14541
rect 13234 14532 13246 14535
rect 13044 14504 13246 14532
rect 13044 14492 13050 14504
rect 13234 14501 13246 14504
rect 13280 14501 13292 14535
rect 16758 14532 16764 14544
rect 16671 14504 16764 14532
rect 13234 14495 13292 14501
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 5442 14464 5448 14476
rect 4847 14436 5448 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6236 14436 6469 14464
rect 6236 14424 6242 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 7653 14467 7711 14473
rect 7653 14433 7665 14467
rect 7699 14464 7711 14467
rect 8202 14464 8208 14476
rect 7699 14436 8208 14464
rect 7699 14433 7711 14436
rect 7653 14427 7711 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 10588 14467 10646 14473
rect 10588 14433 10600 14467
rect 10634 14464 10646 14467
rect 10870 14464 10876 14476
rect 10634 14436 10876 14464
rect 10634 14433 10646 14436
rect 10588 14427 10646 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 13630 14464 13636 14476
rect 13004 14436 13636 14464
rect 4580 14368 4752 14396
rect 5077 14399 5135 14405
rect 4580 14356 4586 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 6086 14396 6092 14408
rect 5123 14368 6092 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 6086 14356 6092 14368
rect 6144 14396 6150 14408
rect 13004 14405 13032 14436
rect 13630 14424 13636 14436
rect 13688 14464 13694 14476
rect 13998 14464 14004 14476
rect 13688 14436 14004 14464
rect 13688 14424 13694 14436
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14464 15715 14467
rect 16022 14464 16028 14476
rect 15703 14436 16028 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 6144 14368 6653 14396
rect 6144 14356 6150 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4433 14331 4491 14337
rect 4433 14328 4445 14331
rect 4212 14300 4445 14328
rect 4212 14288 4218 14300
rect 4433 14297 4445 14300
rect 4479 14297 4491 14331
rect 4433 14291 4491 14297
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14260 2010 14272
rect 2225 14263 2283 14269
rect 2225 14260 2237 14263
rect 2004 14232 2237 14260
rect 2004 14220 2010 14232
rect 2225 14229 2237 14232
rect 2271 14229 2283 14263
rect 2225 14223 2283 14229
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 3602 14260 3608 14272
rect 3559 14232 3608 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3752 14232 3801 14260
rect 3752 14220 3758 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 3789 14223 3847 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6089 14263 6147 14269
rect 6089 14229 6101 14263
rect 6135 14260 6147 14263
rect 6454 14260 6460 14272
rect 6135 14232 6460 14260
rect 6135 14229 6147 14232
rect 6089 14223 6147 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 7834 14260 7840 14272
rect 7331 14232 7840 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 8168 14232 8585 14260
rect 8168 14220 8174 14232
rect 8573 14229 8585 14232
rect 8619 14260 8631 14263
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8619 14232 8953 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8941 14229 8953 14232
rect 8987 14260 8999 14263
rect 9122 14260 9128 14272
rect 8987 14232 9128 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9122 14220 9128 14232
rect 9180 14260 9186 14272
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 9180 14232 9413 14260
rect 9180 14220 9186 14232
rect 9401 14229 9413 14232
rect 9447 14260 9459 14263
rect 10229 14263 10287 14269
rect 10229 14260 10241 14263
rect 9447 14232 10241 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10229 14229 10241 14232
rect 10275 14260 10287 14263
rect 10336 14260 10364 14359
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 14792 14368 15761 14396
rect 14792 14356 14798 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16114 14396 16120 14408
rect 15979 14368 16120 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 12434 14328 12440 14340
rect 11992 14300 12440 14328
rect 10962 14260 10968 14272
rect 10275 14232 10968 14260
rect 10275 14229 10287 14232
rect 10229 14223 10287 14229
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 11514 14260 11520 14272
rect 11020 14232 11520 14260
rect 11020 14220 11026 14232
rect 11514 14220 11520 14232
rect 11572 14260 11578 14272
rect 11992 14269 12020 14300
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 12805 14331 12863 14337
rect 12805 14328 12817 14331
rect 12492 14300 12817 14328
rect 12492 14288 12498 14300
rect 12805 14297 12817 14300
rect 12851 14297 12863 14331
rect 15010 14328 15016 14340
rect 14971 14300 15016 14328
rect 12805 14291 12863 14297
rect 15010 14288 15016 14300
rect 15068 14288 15074 14340
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11572 14232 11989 14260
rect 11572 14220 11578 14232
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 11977 14223 12035 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15654 14260 15660 14272
rect 15335 14232 15660 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15988 14232 16313 14260
rect 15988 14220 15994 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 16684 14269 16712 14504
rect 16758 14492 16764 14504
rect 16816 14532 16822 14544
rect 16816 14504 17448 14532
rect 16816 14492 16822 14504
rect 17218 14464 17224 14476
rect 17179 14436 17224 14464
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17420 14405 17448 14504
rect 21358 14492 21364 14544
rect 21416 14541 21422 14544
rect 21416 14535 21480 14541
rect 21416 14501 21434 14535
rect 21468 14501 21480 14535
rect 21416 14495 21480 14501
rect 21416 14492 21422 14495
rect 22094 14492 22100 14544
rect 22152 14532 22158 14544
rect 22646 14532 22652 14544
rect 22152 14504 22652 14532
rect 22152 14492 22158 14504
rect 22646 14492 22652 14504
rect 22704 14492 22710 14544
rect 23198 14492 23204 14544
rect 23256 14532 23262 14544
rect 23256 14504 23980 14532
rect 23256 14492 23262 14504
rect 23952 14476 23980 14504
rect 18874 14473 18880 14476
rect 18868 14464 18880 14473
rect 18787 14436 18880 14464
rect 18868 14427 18880 14436
rect 18932 14464 18938 14476
rect 19426 14464 19432 14476
rect 18932 14436 19432 14464
rect 18874 14424 18880 14427
rect 18932 14424 18938 14436
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 23109 14467 23167 14473
rect 21192 14436 23060 14464
rect 17313 14399 17371 14405
rect 17313 14396 17325 14399
rect 17000 14368 17325 14396
rect 17000 14356 17006 14368
rect 17313 14365 17325 14368
rect 17359 14365 17371 14399
rect 17313 14359 17371 14365
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17328 14328 17356 14359
rect 18230 14356 18236 14408
rect 18288 14396 18294 14408
rect 18598 14396 18604 14408
rect 18288 14368 18604 14396
rect 18288 14356 18294 14368
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 21192 14405 21220 14436
rect 23032 14408 23060 14436
rect 23109 14433 23121 14467
rect 23155 14464 23167 14467
rect 23641 14467 23699 14473
rect 23641 14464 23653 14467
rect 23155 14436 23653 14464
rect 23155 14433 23167 14436
rect 23109 14427 23167 14433
rect 23641 14433 23653 14436
rect 23687 14433 23699 14467
rect 23641 14427 23699 14433
rect 23934 14424 23940 14476
rect 23992 14424 23998 14476
rect 21177 14399 21235 14405
rect 21177 14396 21189 14399
rect 20772 14368 21189 14396
rect 20772 14356 20778 14368
rect 21177 14365 21189 14368
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 23014 14356 23020 14408
rect 23072 14396 23078 14408
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 23072 14368 23397 14396
rect 23072 14356 23078 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 18322 14328 18328 14340
rect 17328 14300 18328 14328
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 22370 14288 22376 14340
rect 22428 14328 22434 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 22428 14300 22569 14328
rect 22428 14288 22434 14300
rect 22557 14297 22569 14300
rect 22603 14328 22615 14331
rect 23109 14331 23167 14337
rect 23109 14328 23121 14331
rect 22603 14300 23121 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 23109 14297 23121 14300
rect 23155 14297 23167 14331
rect 23109 14291 23167 14297
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16448 14232 16681 14260
rect 16448 14220 16454 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 16853 14263 16911 14269
rect 16853 14229 16865 14263
rect 16899 14260 16911 14263
rect 17586 14260 17592 14272
rect 16899 14232 17592 14260
rect 16899 14229 16911 14232
rect 16853 14223 16911 14229
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 19981 14263 20039 14269
rect 19981 14229 19993 14263
rect 20027 14260 20039 14263
rect 20070 14260 20076 14272
rect 20027 14232 20076 14260
rect 20027 14229 20039 14232
rect 19981 14223 20039 14229
rect 20070 14220 20076 14232
rect 20128 14260 20134 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20128 14232 20269 14260
rect 20128 14220 20134 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 21910 14220 21916 14272
rect 21968 14260 21974 14272
rect 22388 14260 22416 14288
rect 21968 14232 22416 14260
rect 21968 14220 21974 14232
rect 23382 14220 23388 14272
rect 23440 14260 23446 14272
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 23440 14232 24777 14260
rect 23440 14220 23446 14232
rect 24765 14229 24777 14232
rect 24811 14229 24823 14263
rect 25038 14260 25044 14272
rect 24999 14232 25044 14260
rect 24765 14223 24823 14229
rect 25038 14220 25044 14232
rect 25096 14220 25102 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 3050 14056 3056 14068
rect 1811 14028 3056 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 3050 14016 3056 14028
rect 3108 14056 3114 14068
rect 3329 14059 3387 14065
rect 3108 14028 3280 14056
rect 3108 14016 3114 14028
rect 3252 13997 3280 14028
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3375 14028 3617 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 3605 14025 3617 14028
rect 3651 14056 3663 14059
rect 5813 14059 5871 14065
rect 5813 14056 5825 14059
rect 3651 14028 5825 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 5813 14025 5825 14028
rect 5859 14056 5871 14059
rect 6086 14056 6092 14068
rect 5859 14028 6092 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6880 14028 7205 14056
rect 6880 14016 6886 14028
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8294 14056 8300 14068
rect 7984 14028 8300 14056
rect 7984 14016 7990 14028
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 8941 14059 8999 14065
rect 8941 14056 8953 14059
rect 8352 14028 8953 14056
rect 8352 14016 8358 14028
rect 8941 14025 8953 14028
rect 8987 14056 8999 14059
rect 9030 14056 9036 14068
rect 8987 14028 9036 14056
rect 8987 14025 8999 14028
rect 8941 14019 8999 14025
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12802 14056 12808 14068
rect 12483 14028 12808 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 13044 14028 13461 14056
rect 13044 14016 13050 14028
rect 13449 14025 13461 14028
rect 13495 14025 13507 14059
rect 13449 14019 13507 14025
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 15013 14059 15071 14065
rect 15013 14056 15025 14059
rect 14792 14028 15025 14056
rect 14792 14016 14798 14028
rect 15013 14025 15025 14028
rect 15059 14025 15071 14059
rect 15470 14056 15476 14068
rect 15431 14028 15476 14056
rect 15013 14019 15071 14025
rect 15470 14016 15476 14028
rect 15528 14056 15534 14068
rect 21358 14056 21364 14068
rect 15528 14028 16068 14056
rect 21319 14028 21364 14056
rect 15528 14016 15534 14028
rect 3237 13991 3295 13997
rect 3237 13957 3249 13991
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 3252 13920 3280 13951
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3252 13892 3985 13920
rect 3973 13889 3985 13892
rect 4019 13920 4031 13923
rect 7101 13923 7159 13929
rect 4019 13892 4200 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13821 4123 13855
rect 4172 13852 4200 13892
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7147 13892 7757 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7745 13889 7757 13892
rect 7791 13920 7803 13923
rect 8754 13920 8760 13932
rect 7791 13892 8760 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 11054 13920 11060 13932
rect 9447 13892 9628 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 4321 13855 4379 13861
rect 4321 13852 4333 13855
rect 4172 13824 4333 13852
rect 4065 13815 4123 13821
rect 4321 13821 4333 13824
rect 4367 13821 4379 13855
rect 6178 13852 6184 13864
rect 6139 13824 6184 13852
rect 4321 13815 4379 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 2102 13787 2160 13793
rect 2102 13784 2114 13787
rect 1728 13756 2114 13784
rect 1728 13744 1734 13756
rect 2102 13753 2114 13756
rect 2148 13753 2160 13787
rect 4080 13784 4108 13815
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13852 6607 13855
rect 6638 13852 6644 13864
rect 6595 13824 6644 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 7834 13852 7840 13864
rect 7699 13824 7840 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8202 13852 8208 13864
rect 8163 13824 8208 13852
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8312 13824 8585 13852
rect 4890 13784 4896 13796
rect 4080 13756 4896 13784
rect 2102 13747 2160 13753
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 7248 13756 7573 13784
rect 7248 13744 7254 13756
rect 7561 13753 7573 13756
rect 7607 13784 7619 13787
rect 8312 13784 8340 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9180 13824 9505 13852
rect 9180 13812 9186 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9600 13852 9628 13892
rect 10796 13892 11060 13920
rect 9749 13855 9807 13861
rect 9749 13852 9761 13855
rect 9600 13824 9761 13852
rect 9493 13815 9551 13821
rect 9749 13821 9761 13824
rect 9795 13852 9807 13855
rect 10796 13852 10824 13892
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11808 13920 11836 14016
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 15746 13988 15752 14000
rect 15620 13960 15752 13988
rect 15620 13948 15626 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 16040 13988 16068 14028
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 22370 14016 22376 14068
rect 22428 14056 22434 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22428 14028 23397 14056
rect 22428 14016 22434 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 16666 13988 16672 14000
rect 16040 13960 16672 13988
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 11808 13892 13001 13920
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14182 13920 14188 13932
rect 13955 13892 14188 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14182 13880 14188 13892
rect 14240 13920 14246 13932
rect 16040 13929 16068 13960
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 19426 13988 19432 14000
rect 19339 13960 19432 13988
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 23198 13948 23204 14000
rect 23256 13988 23262 14000
rect 24397 13991 24455 13997
rect 24397 13988 24409 13991
rect 23256 13960 24409 13988
rect 23256 13948 23262 13960
rect 24397 13957 24409 13960
rect 24443 13957 24455 13991
rect 24397 13951 24455 13957
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14240 13892 14565 13920
rect 14240 13880 14246 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13889 16083 13923
rect 16206 13920 16212 13932
rect 16167 13892 16212 13920
rect 16025 13883 16083 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 19444 13920 19472 13948
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19444 13892 19809 13920
rect 19797 13889 19809 13892
rect 19843 13920 19855 13923
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 19843 13892 20821 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 21729 13923 21787 13929
rect 21729 13889 21741 13923
rect 21775 13920 21787 13923
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 21775 13892 22477 13920
rect 21775 13889 21787 13892
rect 21729 13883 21787 13889
rect 22465 13889 22477 13892
rect 22511 13920 22523 13923
rect 23382 13920 23388 13932
rect 22511 13892 23388 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 24026 13880 24032 13932
rect 24084 13920 24090 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24084 13892 25053 13920
rect 24084 13880 24090 13892
rect 25041 13889 25053 13892
rect 25087 13920 25099 13923
rect 25409 13923 25467 13929
rect 25409 13920 25421 13923
rect 25087 13892 25421 13920
rect 25087 13889 25099 13892
rect 25041 13883 25099 13889
rect 25409 13889 25421 13892
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 9795 13824 10824 13852
rect 10888 13824 11161 13852
rect 9795 13821 9807 13824
rect 9749 13815 9807 13821
rect 7607 13756 8340 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 10888 13728 10916 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11149 13815 11207 13821
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12584 13824 12909 13852
rect 12584 13812 12590 13824
rect 12897 13821 12909 13824
rect 12943 13852 12955 13855
rect 13446 13852 13452 13864
rect 12943 13824 13452 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 15160 13824 16865 13852
rect 15160 13812 15166 13824
rect 16853 13821 16865 13824
rect 16899 13852 16911 13855
rect 16942 13852 16948 13864
rect 16899 13824 16948 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17218 13852 17224 13864
rect 17179 13824 17224 13852
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18138 13852 18144 13864
rect 18095 13824 18144 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 22112 13824 22293 13852
rect 13538 13744 13544 13796
rect 13596 13784 13602 13796
rect 14369 13787 14427 13793
rect 14369 13784 14381 13787
rect 13596 13756 14381 13784
rect 13596 13744 13602 13756
rect 14369 13753 14381 13756
rect 14415 13784 14427 13787
rect 18294 13787 18352 13793
rect 18294 13784 18306 13787
rect 14415 13756 14688 13784
rect 14415 13753 14427 13756
rect 14369 13747 14427 13753
rect 2222 13676 2228 13728
rect 2280 13716 2286 13728
rect 3329 13719 3387 13725
rect 3329 13716 3341 13719
rect 2280 13688 3341 13716
rect 2280 13676 2286 13688
rect 3329 13685 3341 13688
rect 3375 13685 3387 13719
rect 3329 13679 3387 13685
rect 5445 13719 5503 13725
rect 5445 13685 5457 13719
rect 5491 13716 5503 13719
rect 5534 13716 5540 13728
rect 5491 13688 5540 13716
rect 5491 13685 5503 13688
rect 5445 13679 5503 13685
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 10870 13716 10876 13728
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12802 13716 12808 13728
rect 12299 13688 12808 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13964 13688 14013 13716
rect 13964 13676 13970 13688
rect 14001 13685 14013 13688
rect 14047 13685 14059 13719
rect 14458 13716 14464 13728
rect 14419 13688 14464 13716
rect 14001 13679 14059 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 14660 13716 14688 13756
rect 18156 13756 18306 13784
rect 18156 13728 18184 13756
rect 18294 13753 18306 13756
rect 18340 13753 18352 13787
rect 18294 13747 18352 13753
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13784 20223 13787
rect 20625 13787 20683 13793
rect 20625 13784 20637 13787
rect 20211 13756 20637 13784
rect 20211 13753 20223 13756
rect 20165 13747 20223 13753
rect 20625 13753 20637 13756
rect 20671 13784 20683 13787
rect 20990 13784 20996 13796
rect 20671 13756 20996 13784
rect 20671 13753 20683 13756
rect 20625 13747 20683 13753
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 21358 13744 21364 13796
rect 21416 13784 21422 13796
rect 22112 13784 22140 13824
rect 22281 13821 22293 13824
rect 22327 13852 22339 13855
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22327 13824 22845 13852
rect 22327 13821 22339 13824
rect 22281 13815 22339 13821
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 21416 13756 22140 13784
rect 21416 13744 21422 13756
rect 24118 13744 24124 13796
rect 24176 13784 24182 13796
rect 24305 13787 24363 13793
rect 24305 13784 24317 13787
rect 24176 13756 24317 13784
rect 24176 13744 24182 13756
rect 24305 13753 24317 13756
rect 24351 13784 24363 13787
rect 24351 13756 24900 13784
rect 24351 13753 24363 13756
rect 24305 13747 24363 13753
rect 15565 13719 15623 13725
rect 15565 13716 15577 13719
rect 14660 13688 15577 13716
rect 15565 13685 15577 13688
rect 15611 13685 15623 13719
rect 15930 13716 15936 13728
rect 15891 13688 15936 13716
rect 15565 13679 15623 13685
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 17865 13719 17923 13725
rect 17865 13685 17877 13719
rect 17911 13716 17923 13719
rect 18138 13716 18144 13728
rect 17911 13688 18144 13716
rect 17911 13685 17923 13688
rect 17865 13679 17923 13685
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 20254 13716 20260 13728
rect 20215 13688 20260 13716
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 20717 13719 20775 13725
rect 20717 13716 20729 13719
rect 20588 13688 20729 13716
rect 20588 13676 20594 13688
rect 20717 13685 20729 13688
rect 20763 13685 20775 13719
rect 20717 13679 20775 13685
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 22189 13719 22247 13725
rect 22189 13716 22201 13719
rect 21784 13688 22201 13716
rect 21784 13676 21790 13688
rect 22189 13685 22201 13688
rect 22235 13685 22247 13719
rect 23842 13716 23848 13728
rect 23803 13688 23848 13716
rect 22189 13679 22247 13685
rect 23842 13676 23848 13688
rect 23900 13716 23906 13728
rect 24872 13725 24900 13756
rect 24765 13719 24823 13725
rect 24765 13716 24777 13719
rect 23900 13688 24777 13716
rect 23900 13676 23906 13688
rect 24765 13685 24777 13688
rect 24811 13685 24823 13719
rect 24765 13679 24823 13685
rect 24857 13719 24915 13725
rect 24857 13685 24869 13719
rect 24903 13716 24915 13719
rect 25774 13716 25780 13728
rect 24903 13688 25780 13716
rect 24903 13685 24915 13688
rect 24857 13679 24915 13685
rect 25774 13676 25780 13688
rect 25832 13676 25838 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3421 13515 3479 13521
rect 3421 13512 3433 13515
rect 3200 13484 3433 13512
rect 3200 13472 3206 13484
rect 3421 13481 3433 13484
rect 3467 13481 3479 13515
rect 3421 13475 3479 13481
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4062 13512 4068 13524
rect 3927 13484 4068 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5442 13512 5448 13524
rect 4571 13484 5448 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6144 13484 6285 13512
rect 6144 13472 6150 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 6273 13475 6331 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9030 13512 9036 13524
rect 8991 13484 9036 13512
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 12115 13484 12756 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 2032 13447 2090 13453
rect 2032 13413 2044 13447
rect 2078 13444 2090 13447
rect 2222 13444 2228 13456
rect 2078 13416 2228 13444
rect 2078 13413 2090 13416
rect 2032 13407 2090 13413
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 7285 13447 7343 13453
rect 7285 13413 7297 13447
rect 7331 13444 7343 13447
rect 7622 13447 7680 13453
rect 7622 13444 7634 13447
rect 7331 13416 7634 13444
rect 7331 13413 7343 13416
rect 7285 13407 7343 13413
rect 7622 13413 7634 13416
rect 7668 13444 7680 13447
rect 7742 13444 7748 13456
rect 7668 13416 7748 13444
rect 7668 13413 7680 13416
rect 7622 13407 7680 13413
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 12158 13404 12164 13456
rect 12216 13444 12222 13456
rect 12437 13447 12495 13453
rect 12437 13444 12449 13447
rect 12216 13416 12449 13444
rect 12216 13404 12222 13416
rect 12437 13413 12449 13416
rect 12483 13444 12495 13447
rect 12618 13444 12624 13456
rect 12483 13416 12624 13444
rect 12483 13413 12495 13416
rect 12437 13407 12495 13413
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 12728 13444 12756 13484
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12986 13512 12992 13524
rect 12860 13484 12992 13512
rect 12860 13472 12866 13484
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13538 13512 13544 13524
rect 13499 13484 13544 13512
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 18693 13515 18751 13521
rect 13688 13484 13733 13512
rect 13688 13472 13694 13484
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 18874 13512 18880 13524
rect 18739 13484 18880 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19300 13484 19441 13512
rect 19300 13472 19306 13484
rect 19429 13481 19441 13484
rect 19475 13512 19487 13515
rect 20254 13512 20260 13524
rect 19475 13484 20260 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20622 13512 20628 13524
rect 20496 13484 20628 13512
rect 20496 13472 20502 13484
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21358 13512 21364 13524
rect 21319 13484 21364 13512
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21692 13484 21833 13512
rect 21692 13472 21698 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 21821 13475 21879 13481
rect 22465 13515 22523 13521
rect 22465 13481 22477 13515
rect 22511 13512 22523 13515
rect 22646 13512 22652 13524
rect 22511 13484 22652 13512
rect 22511 13481 22523 13484
rect 22465 13475 22523 13481
rect 22646 13472 22652 13484
rect 22704 13512 22710 13524
rect 24026 13512 24032 13524
rect 22704 13484 24032 13512
rect 22704 13472 22710 13484
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 25866 13512 25872 13524
rect 25547 13484 25872 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 14458 13444 14464 13456
rect 12728 13416 14464 13444
rect 14458 13404 14464 13416
rect 14516 13444 14522 13456
rect 14645 13447 14703 13453
rect 14645 13444 14657 13447
rect 14516 13416 14657 13444
rect 14516 13404 14522 13416
rect 14645 13413 14657 13416
rect 14691 13413 14703 13447
rect 14645 13407 14703 13413
rect 14734 13404 14740 13456
rect 14792 13444 14798 13456
rect 19334 13444 19340 13456
rect 14792 13416 17172 13444
rect 19295 13416 19340 13444
rect 14792 13404 14798 13416
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 1854 13376 1860 13388
rect 1811 13348 1860 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4890 13376 4896 13388
rect 4672 13348 4896 13376
rect 4672 13336 4678 13348
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5160 13379 5218 13385
rect 5160 13345 5172 13379
rect 5206 13376 5218 13379
rect 5442 13376 5448 13388
rect 5206 13348 5448 13376
rect 5206 13345 5218 13348
rect 5160 13339 5218 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7466 13376 7472 13388
rect 7423 13348 7472 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7466 13336 7472 13348
rect 7524 13376 7530 13388
rect 8110 13376 8116 13388
rect 7524 13348 8116 13376
rect 7524 13336 7530 13348
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 9674 13376 9680 13388
rect 8812 13348 9680 13376
rect 8812 13336 8818 13348
rect 9674 13336 9680 13348
rect 9732 13376 9738 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 9732 13348 10241 13376
rect 9732 13336 9738 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 12526 13376 12532 13388
rect 12487 13348 12532 13376
rect 10229 13339 10287 13345
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 14001 13339 14059 13345
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 15102 13376 15108 13388
rect 14139 13348 15108 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 10134 13308 10140 13320
rect 9539 13280 10140 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 10134 13268 10140 13280
rect 10192 13308 10198 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 10192 13280 10333 13308
rect 10192 13268 10198 13280
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10870 13308 10876 13320
rect 10468 13280 10876 13308
rect 10468 13268 10474 13280
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 12897 13311 12955 13317
rect 12897 13308 12909 13311
rect 12759 13280 12909 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 12897 13277 12909 13280
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 14108 13308 14136 13339
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15378 13376 15384 13388
rect 15335 13348 15384 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15378 13336 15384 13348
rect 15436 13376 15442 13388
rect 15562 13376 15568 13388
rect 15436 13348 15568 13376
rect 15436 13336 15442 13348
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 15930 13336 15936 13388
rect 15988 13376 15994 13388
rect 16482 13376 16488 13388
rect 15988 13348 16488 13376
rect 15988 13336 15994 13348
rect 16482 13336 16488 13348
rect 16540 13376 16546 13388
rect 17017 13379 17075 13385
rect 17017 13376 17029 13379
rect 16540 13348 17029 13376
rect 16540 13336 16546 13348
rect 17017 13345 17029 13348
rect 17063 13345 17075 13379
rect 17144 13376 17172 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 23382 13453 23388 13456
rect 23376 13444 23388 13453
rect 23343 13416 23388 13444
rect 23376 13407 23388 13416
rect 23382 13404 23388 13407
rect 23440 13404 23446 13456
rect 21542 13376 21548 13388
rect 17144 13348 21548 13376
rect 17017 13339 17075 13345
rect 21542 13336 21548 13348
rect 21600 13376 21606 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 21600 13348 21741 13376
rect 21600 13336 21606 13348
rect 21729 13345 21741 13348
rect 21775 13345 21787 13379
rect 25314 13376 25320 13388
rect 25275 13348 25320 13376
rect 21729 13339 21787 13345
rect 25314 13336 25320 13348
rect 25372 13336 25378 13388
rect 13219 13280 14136 13308
rect 14277 13311 14335 13317
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 16632 13280 16773 13308
rect 16632 13268 16638 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 20070 13308 20076 13320
rect 19659 13280 20076 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 20070 13268 20076 13280
rect 20128 13308 20134 13320
rect 20622 13308 20628 13320
rect 20128 13280 20628 13308
rect 20128 13268 20134 13280
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21910 13308 21916 13320
rect 21140 13280 21916 13308
rect 21140 13268 21146 13280
rect 21910 13268 21916 13280
rect 21968 13268 21974 13320
rect 23109 13311 23167 13317
rect 23109 13277 23121 13311
rect 23155 13277 23167 13311
rect 23109 13271 23167 13277
rect 11977 13243 12035 13249
rect 11977 13209 11989 13243
rect 12023 13240 12035 13243
rect 12023 13212 12296 13240
rect 12023 13209 12035 13212
rect 11977 13203 12035 13209
rect 1210 13132 1216 13184
rect 1268 13172 1274 13184
rect 2038 13172 2044 13184
rect 1268 13144 2044 13172
rect 1268 13132 1274 13144
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 3145 13175 3203 13181
rect 3145 13141 3157 13175
rect 3191 13172 3203 13175
rect 3234 13172 3240 13184
rect 3191 13144 3240 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 6546 13172 6552 13184
rect 6507 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 10870 13132 10876 13144
rect 10928 13172 10934 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 10928 13144 11253 13172
rect 10928 13132 10934 13144
rect 11241 13141 11253 13144
rect 11287 13141 11299 13175
rect 12268 13172 12296 13212
rect 19886 13200 19892 13252
rect 19944 13240 19950 13252
rect 20717 13243 20775 13249
rect 20717 13240 20729 13243
rect 19944 13212 20729 13240
rect 19944 13200 19950 13212
rect 20717 13209 20729 13212
rect 20763 13240 20775 13243
rect 20763 13212 22232 13240
rect 20763 13209 20775 13212
rect 20717 13203 20775 13209
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12268 13144 12909 13172
rect 11241 13135 11299 13141
rect 12897 13141 12909 13144
rect 12943 13172 12955 13175
rect 13170 13172 13176 13184
rect 12943 13144 13176 13172
rect 12943 13141 12955 13144
rect 12897 13135 12955 13141
rect 13170 13132 13176 13144
rect 13228 13172 13234 13184
rect 15105 13175 15163 13181
rect 15105 13172 15117 13175
rect 13228 13144 15117 13172
rect 13228 13132 13234 13144
rect 15105 13141 15117 13144
rect 15151 13172 15163 13175
rect 16206 13172 16212 13184
rect 15151 13144 16212 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 16206 13132 16212 13144
rect 16264 13172 16270 13184
rect 16393 13175 16451 13181
rect 16393 13172 16405 13175
rect 16264 13144 16405 13172
rect 16264 13132 16270 13144
rect 16393 13141 16405 13144
rect 16439 13141 16451 13175
rect 18138 13172 18144 13184
rect 18099 13144 18144 13172
rect 16393 13135 16451 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 18966 13172 18972 13184
rect 18927 13144 18972 13172
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 20254 13172 20260 13184
rect 20215 13144 20260 13172
rect 20254 13132 20260 13144
rect 20312 13172 20318 13184
rect 20530 13172 20536 13184
rect 20312 13144 20536 13172
rect 20312 13132 20318 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 21726 13172 21732 13184
rect 21315 13144 21732 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 22204 13172 22232 13212
rect 22278 13200 22284 13252
rect 22336 13240 22342 13252
rect 22741 13243 22799 13249
rect 22741 13240 22753 13243
rect 22336 13212 22753 13240
rect 22336 13200 22342 13212
rect 22741 13209 22753 13212
rect 22787 13240 22799 13243
rect 23014 13240 23020 13252
rect 22787 13212 23020 13240
rect 22787 13209 22799 13212
rect 22741 13203 22799 13209
rect 23014 13200 23020 13212
rect 23072 13240 23078 13252
rect 23124 13240 23152 13271
rect 25774 13240 25780 13252
rect 23072 13212 23152 13240
rect 24044 13212 25780 13240
rect 23072 13200 23078 13212
rect 24044 13172 24072 13212
rect 25774 13200 25780 13212
rect 25832 13200 25838 13252
rect 22204 13144 24072 13172
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24489 13175 24547 13181
rect 24489 13172 24501 13175
rect 24176 13144 24501 13172
rect 24176 13132 24182 13144
rect 24489 13141 24501 13144
rect 24535 13172 24547 13175
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 24535 13144 24777 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 24765 13141 24777 13144
rect 24811 13141 24823 13175
rect 24765 13135 24823 13141
rect 24946 13132 24952 13184
rect 25004 13172 25010 13184
rect 25133 13175 25191 13181
rect 25133 13172 25145 13175
rect 25004 13144 25145 13172
rect 25004 13132 25010 13144
rect 25133 13141 25145 13144
rect 25179 13141 25191 13175
rect 25133 13135 25191 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 2682 12968 2688 12980
rect 1903 12940 2688 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3476 12940 3617 12968
rect 3476 12928 3482 12940
rect 3605 12937 3617 12940
rect 3651 12937 3663 12971
rect 3605 12931 3663 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5350 12968 5356 12980
rect 4755 12940 5356 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 7190 12968 7196 12980
rect 7151 12940 7196 12968
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10410 12968 10416 12980
rect 9999 12940 10416 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12584 12940 12633 12968
rect 12584 12928 12590 12940
rect 12621 12937 12633 12940
rect 12667 12968 12679 12971
rect 13538 12968 13544 12980
rect 12667 12940 13544 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 15930 12968 15936 12980
rect 15891 12940 15936 12968
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 16724 12940 17785 12968
rect 16724 12928 16730 12940
rect 17773 12937 17785 12940
rect 17819 12968 17831 12971
rect 18506 12968 18512 12980
rect 17819 12940 18512 12968
rect 17819 12937 17831 12940
rect 17773 12931 17831 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 20622 12968 20628 12980
rect 20583 12940 20628 12968
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 21082 12968 21088 12980
rect 21043 12940 21088 12968
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21453 12971 21511 12977
rect 21453 12937 21465 12971
rect 21499 12968 21511 12971
rect 21542 12968 21548 12980
rect 21499 12940 21548 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 23109 12971 23167 12977
rect 23109 12937 23121 12971
rect 23155 12968 23167 12971
rect 23382 12968 23388 12980
rect 23155 12940 23388 12968
rect 23155 12937 23167 12940
rect 23109 12931 23167 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25314 12968 25320 12980
rect 25275 12940 25320 12968
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2038 12900 2044 12912
rect 1811 12872 2044 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 2038 12860 2044 12872
rect 2096 12900 2102 12912
rect 2222 12900 2228 12912
rect 2096 12872 2228 12900
rect 2096 12860 2102 12872
rect 2222 12860 2228 12872
rect 2280 12860 2286 12912
rect 5368 12900 5396 12928
rect 5626 12900 5632 12912
rect 5368 12872 5632 12900
rect 5626 12860 5632 12872
rect 5684 12900 5690 12912
rect 6914 12900 6920 12912
rect 5684 12872 6920 12900
rect 5684 12860 5690 12872
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 16390 12900 16396 12912
rect 16264 12872 16396 12900
rect 16264 12860 16270 12872
rect 16390 12860 16396 12872
rect 16448 12900 16454 12912
rect 16448 12872 18736 12900
rect 16448 12860 16454 12872
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 1728 12804 2421 12832
rect 1728 12792 1734 12804
rect 2409 12801 2421 12804
rect 2455 12832 2467 12835
rect 2455 12804 3004 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2976 12773 3004 12804
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3602 12832 3608 12844
rect 3476 12804 3608 12832
rect 3476 12792 3482 12804
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 3234 12764 3240 12776
rect 3007 12736 3240 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3234 12724 3240 12736
rect 3292 12764 3298 12776
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3292 12736 3525 12764
rect 3292 12724 3298 12736
rect 3513 12733 3525 12736
rect 3559 12764 3571 12767
rect 4172 12764 4200 12795
rect 5350 12792 5356 12844
rect 5408 12832 5414 12844
rect 5534 12832 5540 12844
rect 5408 12804 5540 12832
rect 5408 12792 5414 12804
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5592 12804 5733 12832
rect 5592 12792 5598 12804
rect 5721 12801 5733 12804
rect 5767 12832 5779 12835
rect 6181 12835 6239 12841
rect 6181 12832 6193 12835
rect 5767 12804 6193 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6181 12801 6193 12804
rect 6227 12801 6239 12835
rect 6822 12832 6828 12844
rect 6783 12804 6828 12832
rect 6181 12795 6239 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12832 7806 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7800 12804 8217 12832
rect 7800 12792 7806 12804
rect 8205 12801 8217 12804
rect 8251 12832 8263 12835
rect 8386 12832 8392 12844
rect 8251 12804 8392 12832
rect 8251 12801 8263 12804
rect 8205 12795 8263 12801
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12832 12955 12835
rect 13722 12832 13728 12844
rect 12943 12804 13728 12832
rect 12943 12801 12955 12804
rect 12897 12795 12955 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16347 12804 16957 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16945 12801 16957 12804
rect 16991 12832 17003 12835
rect 18138 12832 18144 12844
rect 16991 12804 18144 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18708 12832 18736 12872
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 19613 12903 19671 12909
rect 19613 12900 19625 12903
rect 19116 12872 19625 12900
rect 19116 12860 19122 12872
rect 19613 12869 19625 12872
rect 19659 12869 19671 12903
rect 19613 12863 19671 12869
rect 20070 12832 20076 12844
rect 18708 12804 20076 12832
rect 20070 12792 20076 12804
rect 20128 12832 20134 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 20128 12804 20177 12832
rect 20128 12792 20134 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 22646 12832 22652 12844
rect 22607 12804 22652 12832
rect 20165 12795 20223 12801
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 24118 12792 24124 12844
rect 24176 12832 24182 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24176 12804 24593 12832
rect 24176 12792 24182 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 24912 12804 25605 12832
rect 24912 12792 24918 12804
rect 25593 12801 25605 12804
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 3559 12736 4200 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5040 12736 6561 12764
rect 5040 12724 5046 12736
rect 6549 12733 6561 12736
rect 6595 12764 6607 12767
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 6595 12736 7665 12764
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 8849 12767 8907 12773
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 8938 12764 8944 12776
rect 8895 12736 8944 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 8938 12724 8944 12736
rect 8996 12764 9002 12776
rect 9858 12764 9864 12776
rect 8996 12736 9864 12764
rect 8996 12724 9002 12736
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10870 12764 10876 12776
rect 10183 12736 10876 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 13998 12764 14004 12776
rect 13955 12736 14004 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14182 12773 14188 12776
rect 14176 12764 14188 12773
rect 14143 12736 14188 12764
rect 14176 12727 14188 12736
rect 14182 12724 14188 12727
rect 14240 12724 14246 12776
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12764 17555 12767
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 17543 12736 18429 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18417 12733 18429 12736
rect 18463 12764 18475 12767
rect 18690 12764 18696 12776
rect 18463 12736 18696 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 21910 12764 21916 12776
rect 21823 12736 21916 12764
rect 21910 12724 21916 12736
rect 21968 12764 21974 12776
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 21968 12736 22477 12764
rect 21968 12724 21974 12736
rect 22465 12733 22477 12736
rect 22511 12764 22523 12767
rect 23382 12764 23388 12776
rect 22511 12736 23388 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 23477 12767 23535 12773
rect 23477 12733 23489 12767
rect 23523 12764 23535 12767
rect 24489 12767 24547 12773
rect 24489 12764 24501 12767
rect 23523 12736 24501 12764
rect 23523 12733 23535 12736
rect 23477 12727 23535 12733
rect 24489 12733 24501 12736
rect 24535 12764 24547 12767
rect 24670 12764 24676 12776
rect 24535 12736 24676 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 5074 12696 5080 12708
rect 2832 12668 3280 12696
rect 4987 12668 5080 12696
rect 2832 12656 2838 12668
rect 3252 12640 3280 12668
rect 5074 12656 5080 12668
rect 5132 12696 5138 12708
rect 5537 12699 5595 12705
rect 5537 12696 5549 12699
rect 5132 12668 5549 12696
rect 5132 12656 5138 12668
rect 5537 12665 5549 12668
rect 5583 12696 5595 12699
rect 6825 12699 6883 12705
rect 6825 12696 6837 12699
rect 5583 12668 6837 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 6825 12665 6837 12668
rect 6871 12665 6883 12699
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 6825 12659 6883 12665
rect 7024 12668 7573 12696
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 2372 12600 2417 12628
rect 2372 12588 2378 12600
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 3970 12628 3976 12640
rect 3931 12600 3976 12628
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5626 12628 5632 12640
rect 5587 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7024 12637 7052 12668
rect 7561 12665 7573 12668
rect 7607 12665 7619 12699
rect 9122 12696 9128 12708
rect 9083 12668 9128 12696
rect 7561 12659 7619 12665
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 10404 12699 10462 12705
rect 10404 12665 10416 12699
rect 10450 12696 10462 12699
rect 10778 12696 10784 12708
rect 10450 12668 10784 12696
rect 10450 12665 10462 12668
rect 10404 12659 10462 12665
rect 10778 12656 10784 12668
rect 10836 12656 10842 12708
rect 18506 12696 18512 12708
rect 16776 12668 18092 12696
rect 18467 12668 18512 12696
rect 16776 12640 16804 12668
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6972 12600 7021 12628
rect 6972 12588 6978 12600
rect 7009 12597 7021 12600
rect 7055 12597 7067 12631
rect 7009 12591 7067 12597
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11112 12600 11529 12628
rect 11112 12588 11118 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 12032 12600 12081 12628
rect 12032 12588 12038 12600
rect 12069 12597 12081 12600
rect 12115 12628 12127 12631
rect 12158 12628 12164 12640
rect 12115 12600 12164 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 13725 12631 13783 12637
rect 13725 12597 13737 12631
rect 13771 12628 13783 12631
rect 14458 12628 14464 12640
rect 13771 12600 14464 12628
rect 13771 12597 13783 12600
rect 13725 12591 13783 12597
rect 14458 12588 14464 12600
rect 14516 12628 14522 12640
rect 15286 12628 15292 12640
rect 14516 12600 15292 12628
rect 14516 12588 14522 12600
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 16390 12628 16396 12640
rect 16351 12600 16396 12628
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 16758 12628 16764 12640
rect 16719 12600 16764 12628
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 16942 12628 16948 12640
rect 16899 12600 16948 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 18064 12637 18092 12668
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 19153 12699 19211 12705
rect 19153 12665 19165 12699
rect 19199 12696 19211 12699
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 19199 12668 19993 12696
rect 19199 12665 19211 12668
rect 19153 12659 19211 12665
rect 19981 12665 19993 12668
rect 20027 12696 20039 12699
rect 20162 12696 20168 12708
rect 20027 12668 20168 12696
rect 20027 12665 20039 12668
rect 19981 12659 20039 12665
rect 20162 12656 20168 12668
rect 20220 12656 20226 12708
rect 24397 12699 24455 12705
rect 24397 12696 24409 12699
rect 23860 12668 24409 12696
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12597 18107 12631
rect 18049 12591 18107 12597
rect 19521 12631 19579 12637
rect 19521 12597 19533 12631
rect 19567 12628 19579 12631
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19567 12600 20085 12628
rect 19567 12597 19579 12600
rect 19521 12591 19579 12597
rect 20073 12597 20085 12600
rect 20119 12628 20131 12631
rect 20622 12628 20628 12640
rect 20119 12600 20628 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 22002 12628 22008 12640
rect 21963 12600 22008 12628
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22373 12631 22431 12637
rect 22373 12628 22385 12631
rect 22244 12600 22385 12628
rect 22244 12588 22250 12600
rect 22373 12597 22385 12600
rect 22419 12597 22431 12631
rect 22373 12591 22431 12597
rect 23658 12588 23664 12640
rect 23716 12628 23722 12640
rect 23860 12637 23888 12668
rect 24397 12665 24409 12668
rect 24443 12665 24455 12699
rect 24397 12659 24455 12665
rect 23845 12631 23903 12637
rect 23845 12628 23857 12631
rect 23716 12600 23857 12628
rect 23716 12588 23722 12600
rect 23845 12597 23857 12600
rect 23891 12597 23903 12631
rect 24026 12628 24032 12640
rect 23987 12600 24032 12628
rect 23845 12591 23903 12597
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1394 12384 1400 12436
rect 1452 12424 1458 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1452 12396 1593 12424
rect 1452 12384 1458 12396
rect 1581 12393 1593 12396
rect 1627 12424 1639 12427
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 1627 12396 2145 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 6454 12424 6460 12436
rect 6415 12396 6460 12424
rect 2133 12387 2191 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 8386 12424 8392 12436
rect 8347 12396 8392 12424
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 8938 12424 8944 12436
rect 8899 12396 8944 12424
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11698 12424 11704 12436
rect 11659 12396 11704 12424
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 13354 12424 13360 12436
rect 12820 12396 13360 12424
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2096 12328 2789 12356
rect 2096 12316 2102 12328
rect 2148 12220 2176 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 4614 12356 4620 12368
rect 2777 12319 2835 12325
rect 4080 12328 4620 12356
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2498 12288 2504 12300
rect 2271 12260 2504 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2498 12248 2504 12260
rect 2556 12288 2562 12300
rect 2866 12288 2872 12300
rect 2556 12260 2872 12288
rect 2556 12248 2562 12260
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 4080 12297 4108 12328
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 7558 12356 7564 12368
rect 7024 12328 7564 12356
rect 4338 12297 4344 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4332 12251 4344 12297
rect 4396 12288 4402 12300
rect 6086 12288 6092 12300
rect 4396 12260 4432 12288
rect 6047 12260 6092 12288
rect 4338 12248 4344 12251
rect 4396 12248 4402 12260
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 7024 12297 7052 12328
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11609 12359 11667 12365
rect 11609 12356 11621 12359
rect 11388 12328 11621 12356
rect 11388 12316 11394 12328
rect 11609 12325 11621 12328
rect 11655 12356 11667 12359
rect 12820 12356 12848 12396
rect 13354 12384 13360 12396
rect 13412 12424 13418 12436
rect 14734 12424 14740 12436
rect 13412 12396 14740 12424
rect 13412 12384 13418 12396
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 15841 12427 15899 12433
rect 15841 12424 15853 12427
rect 15804 12396 15853 12424
rect 15804 12384 15810 12396
rect 15841 12393 15853 12396
rect 15887 12393 15899 12427
rect 15841 12387 15899 12393
rect 16485 12427 16543 12433
rect 16485 12393 16497 12427
rect 16531 12424 16543 12427
rect 16942 12424 16948 12436
rect 16531 12396 16948 12424
rect 16531 12393 16543 12396
rect 16485 12387 16543 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 18877 12427 18935 12433
rect 18877 12393 18889 12427
rect 18923 12424 18935 12427
rect 19242 12424 19248 12436
rect 18923 12396 19248 12424
rect 18923 12393 18935 12396
rect 18877 12387 18935 12393
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19334 12384 19340 12436
rect 19392 12384 19398 12436
rect 20070 12424 20076 12436
rect 20031 12396 20076 12424
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 21174 12424 21180 12436
rect 20220 12396 21180 12424
rect 20220 12384 20226 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 21634 12424 21640 12436
rect 21595 12396 21640 12424
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22097 12427 22155 12433
rect 22097 12393 22109 12427
rect 22143 12424 22155 12427
rect 22186 12424 22192 12436
rect 22143 12396 22192 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 22186 12384 22192 12396
rect 22244 12384 22250 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22336 12396 23305 12424
rect 22336 12384 22342 12396
rect 23293 12393 23305 12396
rect 23339 12424 23351 12427
rect 23382 12424 23388 12436
rect 23339 12396 23388 12424
rect 23339 12393 23351 12396
rect 23293 12387 23351 12393
rect 23382 12384 23388 12396
rect 23440 12424 23446 12436
rect 23661 12427 23719 12433
rect 23661 12424 23673 12427
rect 23440 12396 23673 12424
rect 23440 12384 23446 12396
rect 23661 12393 23673 12396
rect 23707 12393 23719 12427
rect 23661 12387 23719 12393
rect 13998 12356 14004 12368
rect 11655 12328 12848 12356
rect 12912 12328 14004 12356
rect 11655 12325 11667 12328
rect 11609 12319 11667 12325
rect 7282 12297 7288 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12257 7067 12291
rect 7276 12288 7288 12297
rect 7243 12260 7288 12288
rect 7009 12251 7067 12257
rect 7276 12251 7288 12260
rect 7282 12248 7288 12251
rect 7340 12248 7346 12300
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9766 12288 9772 12300
rect 9456 12260 9772 12288
rect 9456 12248 9462 12260
rect 9766 12248 9772 12260
rect 9824 12288 9830 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9824 12260 10057 12288
rect 9824 12248 9830 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 11054 12288 11060 12300
rect 10045 12251 10103 12257
rect 10336 12260 11060 12288
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2148 12192 2329 12220
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 6914 12220 6920 12232
rect 6875 12192 6920 12220
rect 2317 12183 2375 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10336 12229 10364 12260
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 12912 12297 12940 12328
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 16758 12316 16764 12368
rect 16816 12356 16822 12368
rect 17028 12359 17086 12365
rect 17028 12356 17040 12359
rect 16816 12328 17040 12356
rect 16816 12316 16822 12328
rect 17028 12325 17040 12328
rect 17074 12325 17086 12359
rect 19352 12356 19380 12384
rect 20349 12359 20407 12365
rect 20349 12356 20361 12359
rect 19352 12328 20361 12356
rect 17028 12319 17086 12325
rect 20349 12325 20361 12328
rect 20395 12325 20407 12359
rect 20349 12319 20407 12325
rect 22554 12316 22560 12368
rect 22612 12356 22618 12368
rect 23676 12356 23704 12387
rect 24946 12356 24952 12368
rect 22612 12328 23152 12356
rect 22612 12316 22618 12328
rect 13170 12297 13176 12300
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 13164 12288 13176 12297
rect 13131 12260 13176 12288
rect 12897 12251 12955 12257
rect 13164 12251 13176 12260
rect 13170 12248 13176 12251
rect 13228 12248 13234 12300
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14792 12260 15669 12288
rect 14792 12248 14798 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 19334 12288 19340 12300
rect 19295 12260 19340 12288
rect 15657 12251 15715 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20438 12288 20444 12300
rect 20128 12260 20444 12288
rect 20128 12248 20134 12260
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12257 20775 12291
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20717 12251 20775 12257
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10778 12220 10784 12232
rect 10691 12192 10784 12220
rect 10321 12183 10379 12189
rect 10778 12180 10784 12192
rect 10836 12220 10842 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 10836 12192 11161 12220
rect 10836 12180 10842 12192
rect 11149 12189 11161 12192
rect 11195 12220 11207 12223
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11195 12192 11897 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11885 12189 11897 12192
rect 11931 12220 11943 12223
rect 12066 12220 12072 12232
rect 11931 12192 12072 12220
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16632 12192 16773 12220
rect 16632 12180 16638 12192
rect 16761 12189 16773 12192
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18506 12220 18512 12232
rect 18288 12192 18512 12220
rect 18288 12180 18294 12192
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 20732 12220 20760 12251
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22370 12248 22376 12300
rect 22428 12248 22434 12300
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12288 22707 12291
rect 23014 12288 23020 12300
rect 22695 12260 23020 12288
rect 22695 12257 22707 12260
rect 22649 12251 22707 12257
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 20990 12220 20996 12232
rect 19576 12192 19621 12220
rect 20732 12192 20996 12220
rect 19576 12180 19582 12192
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 22388 12220 22416 12248
rect 22554 12220 22560 12232
rect 21140 12192 21185 12220
rect 22388 12192 22560 12220
rect 21140 12180 21146 12192
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12220 22799 12223
rect 22830 12220 22836 12232
rect 22787 12192 22836 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 1765 12155 1823 12161
rect 1765 12121 1777 12155
rect 1811 12152 1823 12155
rect 2222 12152 2228 12164
rect 1811 12124 2228 12152
rect 1811 12121 1823 12124
rect 1765 12115 1823 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 2424 12124 3801 12152
rect 2424 12096 2452 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 17770 12112 17776 12164
rect 17828 12152 17834 12164
rect 18969 12155 19027 12161
rect 18969 12152 18981 12155
rect 17828 12124 18981 12152
rect 17828 12112 17834 12124
rect 18969 12121 18981 12124
rect 19015 12121 19027 12155
rect 18969 12115 19027 12121
rect 22646 12112 22652 12164
rect 22704 12152 22710 12164
rect 22756 12152 22784 12183
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 22925 12223 22983 12229
rect 22925 12189 22937 12223
rect 22971 12220 22983 12223
rect 23124 12220 23152 12328
rect 23676 12328 24952 12356
rect 23676 12288 23704 12328
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 24118 12297 24124 12300
rect 23845 12291 23903 12297
rect 23845 12288 23857 12291
rect 23676 12260 23857 12288
rect 23845 12257 23857 12260
rect 23891 12257 23903 12291
rect 24112 12288 24124 12297
rect 24079 12260 24124 12288
rect 23845 12251 23903 12257
rect 24112 12251 24124 12260
rect 24118 12248 24124 12251
rect 24176 12248 24182 12300
rect 22971 12192 23152 12220
rect 22971 12189 22983 12192
rect 22925 12183 22983 12189
rect 22704 12124 22784 12152
rect 22704 12112 22710 12124
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2406 12084 2412 12096
rect 2188 12056 2412 12084
rect 2188 12044 2194 12056
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3970 12084 3976 12096
rect 3559 12056 3976 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3970 12044 3976 12056
rect 4028 12084 4034 12096
rect 5442 12084 5448 12096
rect 4028 12056 5448 12084
rect 4028 12044 4034 12056
rect 5442 12044 5448 12056
rect 5500 12084 5506 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5500 12056 5733 12084
rect 5500 12044 5506 12056
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 5721 12047 5779 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 11238 12084 11244 12096
rect 11199 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 14240 12056 14289 12084
rect 14240 12044 14246 12056
rect 14277 12053 14289 12056
rect 14323 12084 14335 12087
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14323 12056 14657 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14645 12053 14657 12056
rect 14691 12084 14703 12087
rect 15562 12084 15568 12096
rect 14691 12056 15568 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 16632 12056 18153 12084
rect 16632 12044 16638 12056
rect 18141 12053 18153 12056
rect 18187 12084 18199 12087
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 18187 12056 18429 12084
rect 18187 12053 18199 12056
rect 18141 12047 18199 12053
rect 18417 12053 18429 12056
rect 18463 12084 18475 12087
rect 18598 12084 18604 12096
rect 18463 12056 18604 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 20530 12084 20536 12096
rect 20491 12056 20536 12084
rect 20530 12044 20536 12056
rect 20588 12084 20594 12096
rect 20714 12084 20720 12096
rect 20588 12056 20720 12084
rect 20588 12044 20594 12056
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 22278 12084 22284 12096
rect 22239 12056 22284 12084
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22830 12044 22836 12096
rect 22888 12084 22894 12096
rect 22940 12084 22968 12183
rect 25222 12084 25228 12096
rect 22888 12056 22968 12084
rect 25183 12056 25228 12084
rect 22888 12044 22894 12056
rect 25222 12044 25228 12056
rect 25280 12044 25286 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 2314 11880 2320 11892
rect 1811 11852 2320 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 4522 11880 4528 11892
rect 3467 11852 4528 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 9766 11880 9772 11892
rect 9355 11852 9772 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 9950 11880 9956 11892
rect 9911 11852 9956 11880
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10192 11852 10241 11880
rect 10192 11840 10198 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 11330 11880 11336 11892
rect 11291 11852 11336 11880
rect 10229 11843 10287 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11698 11880 11704 11892
rect 11659 11852 11704 11880
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12802 11880 12808 11892
rect 12299 11852 12808 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13170 11840 13176 11892
rect 13228 11880 13234 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13228 11852 13461 11880
rect 13228 11840 13234 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 13449 11843 13507 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 16264 11852 16313 11880
rect 16264 11840 16270 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 16301 11843 16359 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 17770 11880 17776 11892
rect 17644 11852 17776 11880
rect 17644 11840 17650 11852
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18414 11880 18420 11892
rect 18375 11852 18420 11880
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 20165 11883 20223 11889
rect 20165 11880 20177 11883
rect 19484 11852 20177 11880
rect 19484 11840 19490 11852
rect 20165 11849 20177 11852
rect 20211 11849 20223 11883
rect 20165 11843 20223 11849
rect 22465 11883 22523 11889
rect 22465 11849 22477 11883
rect 22511 11880 22523 11883
rect 22646 11880 22652 11892
rect 22511 11852 22652 11880
rect 22511 11849 22523 11852
rect 22465 11843 22523 11849
rect 22646 11840 22652 11852
rect 22704 11880 22710 11892
rect 24854 11880 24860 11892
rect 22704 11852 24860 11880
rect 22704 11840 22710 11852
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 2038 11772 2044 11824
rect 2096 11812 2102 11824
rect 2096 11784 2360 11812
rect 2096 11772 2102 11784
rect 2332 11756 2360 11784
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 4338 11812 4344 11824
rect 4120 11784 4344 11812
rect 4120 11772 4126 11784
rect 4338 11772 4344 11784
rect 4396 11812 4402 11824
rect 4433 11815 4491 11821
rect 4433 11812 4445 11815
rect 4396 11784 4445 11812
rect 4396 11772 4402 11784
rect 4433 11781 4445 11784
rect 4479 11781 4491 11815
rect 4433 11775 4491 11781
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 4890 11812 4896 11824
rect 4764 11784 4896 11812
rect 4764 11772 4770 11784
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 5997 11815 6055 11821
rect 5997 11812 6009 11815
rect 5460 11784 6009 11812
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 3970 11744 3976 11756
rect 2372 11716 2465 11744
rect 3931 11716 3976 11744
rect 2372 11704 2378 11716
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5460 11753 5488 11784
rect 5997 11781 6009 11784
rect 6043 11781 6055 11815
rect 7742 11812 7748 11824
rect 7703 11784 7748 11812
rect 5997 11775 6055 11781
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 11238 11812 11244 11824
rect 10704 11784 11244 11812
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5224 11716 5457 11744
rect 5224 11704 5230 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 5537 11707 5595 11713
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3375 11648 3801 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3789 11645 3801 11648
rect 3835 11676 3847 11679
rect 3878 11676 3884 11688
rect 3835 11648 3884 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 4522 11676 4528 11688
rect 4396 11648 4528 11676
rect 4396 11636 4402 11648
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 5552 11676 5580 11707
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 10704 11753 10732 11784
rect 11238 11772 11244 11784
rect 11296 11772 11302 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 19889 11815 19947 11821
rect 12492 11784 12537 11812
rect 12492 11772 12498 11784
rect 19889 11781 19901 11815
rect 19935 11812 19947 11815
rect 19978 11812 19984 11824
rect 19935 11784 19984 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 19978 11772 19984 11784
rect 20036 11812 20042 11824
rect 20438 11812 20444 11824
rect 20036 11784 20444 11812
rect 20036 11772 20042 11784
rect 20438 11772 20444 11784
rect 20496 11772 20502 11824
rect 25314 11812 25320 11824
rect 25275 11784 25320 11812
rect 25314 11772 25320 11784
rect 25372 11772 25378 11824
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 9548 11716 10701 11744
rect 9548 11704 9554 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 11054 11744 11060 11756
rect 10919 11716 11060 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 7374 11676 7380 11688
rect 4939 11648 5580 11676
rect 7335 11648 7380 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 5460 11620 5488 11648
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8220 11676 8248 11704
rect 8297 11679 8355 11685
rect 8297 11676 8309 11679
rect 8220 11648 8309 11676
rect 8297 11645 8309 11648
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9088 11648 9597 11676
rect 9088 11636 9094 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 5442 11568 5448 11620
rect 5500 11568 5506 11620
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 6641 11611 6699 11617
rect 6641 11608 6653 11611
rect 6236 11580 6653 11608
rect 6236 11568 6242 11580
rect 6641 11577 6653 11580
rect 6687 11608 6699 11611
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 6687 11580 8217 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 8205 11577 8217 11580
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 8941 11611 8999 11617
rect 8941 11577 8953 11611
rect 8987 11608 8999 11611
rect 10888 11608 10916 11707
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12584 11716 13001 11744
rect 12584 11704 12590 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 18506 11744 18512 11756
rect 18467 11716 18512 11744
rect 12989 11707 13047 11713
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23440 11716 23949 11744
rect 23440 11704 23446 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12676 11648 12817 11676
rect 12676 11636 12682 11648
rect 12805 11645 12817 11648
rect 12851 11676 12863 11679
rect 13262 11676 13268 11688
rect 12851 11648 13268 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14918 11676 14924 11688
rect 14056 11648 14924 11676
rect 14056 11636 14062 11648
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11676 17371 11679
rect 18322 11676 18328 11688
rect 17359 11648 18328 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18765 11679 18823 11685
rect 18765 11676 18777 11679
rect 18472 11648 18777 11676
rect 18472 11636 18478 11648
rect 18765 11645 18777 11648
rect 18811 11645 18823 11679
rect 18765 11639 18823 11645
rect 20530 11636 20536 11688
rect 20588 11676 20594 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20588 11648 20729 11676
rect 20588 11636 20594 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 24204 11679 24262 11685
rect 24204 11645 24216 11679
rect 24250 11676 24262 11679
rect 25222 11676 25228 11688
rect 24250 11648 25228 11676
rect 24250 11645 24262 11648
rect 24204 11639 24262 11645
rect 24320 11620 24348 11648
rect 25222 11636 25228 11648
rect 25280 11636 25286 11688
rect 8987 11580 10916 11608
rect 15188 11611 15246 11617
rect 8987 11577 8999 11580
rect 8941 11571 8999 11577
rect 9968 11552 9996 11580
rect 15188 11577 15200 11611
rect 15234 11608 15246 11611
rect 15286 11608 15292 11620
rect 15234 11580 15292 11608
rect 15234 11577 15246 11580
rect 15188 11571 15246 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 20962 11611 21020 11617
rect 20962 11608 20974 11611
rect 20548 11580 20974 11608
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1673 11543 1731 11549
rect 1673 11540 1685 11543
rect 1636 11512 1685 11540
rect 1636 11500 1642 11512
rect 1673 11509 1685 11512
rect 1719 11540 1731 11543
rect 2038 11540 2044 11552
rect 1719 11512 2044 11540
rect 1719 11509 1731 11512
rect 1673 11503 1731 11509
rect 2038 11500 2044 11512
rect 2096 11540 2102 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 2096 11512 2145 11540
rect 2096 11500 2102 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2133 11503 2191 11509
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4948 11512 4997 11540
rect 4948 11500 4954 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5132 11512 5365 11540
rect 5132 11500 5138 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 9398 11540 9404 11552
rect 7616 11512 9404 11540
rect 7616 11500 7622 11512
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9950 11500 9956 11552
rect 10008 11500 10014 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10192 11512 10609 11540
rect 10192 11500 10198 11512
rect 10597 11509 10609 11512
rect 10643 11540 10655 11543
rect 10778 11540 10784 11552
rect 10643 11512 10784 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12860 11512 12909 11540
rect 12860 11500 12866 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13320 11512 14197 11540
rect 13320 11500 13326 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20548 11549 20576 11580
rect 20962 11577 20974 11580
rect 21008 11608 21020 11611
rect 21082 11608 21088 11620
rect 21008 11580 21088 11608
rect 21008 11577 21020 11580
rect 20962 11571 21020 11577
rect 21082 11568 21088 11580
rect 21140 11568 21146 11620
rect 23477 11611 23535 11617
rect 23477 11577 23489 11611
rect 23523 11608 23535 11611
rect 24302 11608 24308 11620
rect 23523 11580 24308 11608
rect 23523 11577 23535 11580
rect 23477 11571 23535 11577
rect 24302 11568 24308 11580
rect 24360 11568 24366 11620
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 20496 11512 20545 11540
rect 20496 11500 20502 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 21324 11512 22109 11540
rect 21324 11500 21330 11512
rect 22097 11509 22109 11512
rect 22143 11540 22155 11543
rect 22554 11540 22560 11552
rect 22143 11512 22560 11540
rect 22143 11509 22155 11512
rect 22097 11503 22155 11509
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 22833 11543 22891 11549
rect 22833 11509 22845 11543
rect 22879 11540 22891 11543
rect 23014 11540 23020 11552
rect 22879 11512 23020 11540
rect 22879 11509 22891 11512
rect 22833 11503 22891 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 25682 11540 25688 11552
rect 25643 11512 25688 11540
rect 25682 11500 25688 11512
rect 25740 11540 25746 11552
rect 25961 11543 26019 11549
rect 25961 11540 25973 11543
rect 25740 11512 25973 11540
rect 25740 11500 25746 11512
rect 25961 11509 25973 11512
rect 26007 11509 26019 11543
rect 25961 11503 26019 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1486 11296 1492 11348
rect 1544 11336 1550 11348
rect 1765 11339 1823 11345
rect 1765 11336 1777 11339
rect 1544 11308 1777 11336
rect 1544 11296 1550 11308
rect 1765 11305 1777 11308
rect 1811 11305 1823 11339
rect 1765 11299 1823 11305
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 2682 11336 2688 11348
rect 2271 11308 2688 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 3200 11308 3525 11336
rect 3200 11296 3206 11308
rect 3513 11305 3525 11308
rect 3559 11336 3571 11339
rect 3878 11336 3884 11348
rect 3559 11308 3884 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4488 11308 4629 11336
rect 4488 11296 4494 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 6178 11336 6184 11348
rect 6139 11308 6184 11336
rect 4617 11299 4675 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 8113 11339 8171 11345
rect 8113 11305 8125 11339
rect 8159 11336 8171 11339
rect 8478 11336 8484 11348
rect 8159 11308 8484 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 10686 11336 10692 11348
rect 9723 11308 10692 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 13262 11336 13268 11348
rect 12176 11308 13268 11336
rect 1578 11268 1584 11280
rect 1539 11240 1584 11268
rect 1578 11228 1584 11240
rect 1636 11228 1642 11280
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 2372 11240 2789 11268
rect 2372 11228 2378 11240
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 2777 11231 2835 11237
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4890 11268 4896 11280
rect 4212 11240 4896 11268
rect 4212 11228 4218 11240
rect 4890 11228 4896 11240
rect 4948 11268 4954 11280
rect 5077 11271 5135 11277
rect 5077 11268 5089 11271
rect 4948 11240 5089 11268
rect 4948 11228 4954 11240
rect 5077 11237 5089 11240
rect 5123 11237 5135 11271
rect 5077 11231 5135 11237
rect 6549 11271 6607 11277
rect 6549 11237 6561 11271
rect 6595 11268 6607 11271
rect 6638 11268 6644 11280
rect 6595 11240 6644 11268
rect 6595 11237 6607 11240
rect 6549 11231 6607 11237
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 7285 11271 7343 11277
rect 7285 11237 7297 11271
rect 7331 11268 7343 11271
rect 8202 11268 8208 11280
rect 7331 11240 8208 11268
rect 7331 11237 7343 11240
rect 7285 11231 7343 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 9950 11268 9956 11280
rect 9539 11240 9956 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 12176 11268 12204 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 15013 11339 15071 11345
rect 13495 11308 14964 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 10796 11240 12204 11268
rect 12529 11271 12587 11277
rect 1210 11160 1216 11212
rect 1268 11200 1274 11212
rect 1486 11200 1492 11212
rect 1268 11172 1492 11200
rect 1268 11160 1274 11172
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11200 2191 11203
rect 2406 11200 2412 11212
rect 2179 11172 2412 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3878 11200 3884 11212
rect 3839 11172 3884 11200
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2280 11104 2329 11132
rect 2280 11092 2286 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 3697 11067 3755 11073
rect 3697 11064 3709 11067
rect 1912 11036 3709 11064
rect 1912 11024 1918 11036
rect 3697 11033 3709 11036
rect 3743 11064 3755 11067
rect 4522 11064 4528 11076
rect 3743 11036 4108 11064
rect 4483 11036 4528 11064
rect 3743 11033 3755 11036
rect 3697 11027 3755 11033
rect 4080 10996 4108 11036
rect 4522 11024 4528 11036
rect 4580 11064 4586 11076
rect 5000 11064 5028 11163
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 9858 11200 9864 11212
rect 9456 11172 9864 11200
rect 9456 11160 9462 11172
rect 9858 11160 9864 11172
rect 9916 11200 9922 11212
rect 10696 11203 10754 11209
rect 10696 11200 10708 11203
rect 9916 11172 10708 11200
rect 9916 11160 9922 11172
rect 10696 11169 10708 11172
rect 10742 11200 10754 11203
rect 10796 11200 10824 11240
rect 12529 11237 12541 11271
rect 12575 11268 12587 11271
rect 12618 11268 12624 11280
rect 12575 11240 12624 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13998 11268 14004 11280
rect 13280 11240 14004 11268
rect 13280 11212 13308 11240
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14936 11268 14964 11308
rect 15013 11305 15025 11339
rect 15059 11336 15071 11339
rect 15286 11336 15292 11348
rect 15059 11308 15292 11336
rect 15059 11305 15071 11308
rect 15013 11299 15071 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18322 11336 18328 11348
rect 18235 11308 18328 11336
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18840 11308 19257 11336
rect 18840 11296 18846 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19392 11308 19625 11336
rect 19392 11296 19398 11308
rect 19613 11305 19625 11308
rect 19659 11336 19671 11339
rect 20254 11336 20260 11348
rect 19659 11308 20260 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 21085 11339 21143 11345
rect 21085 11336 21097 11339
rect 20956 11308 21097 11336
rect 20956 11296 20962 11308
rect 21085 11305 21097 11308
rect 21131 11305 21143 11339
rect 21085 11299 21143 11305
rect 21726 11296 21732 11348
rect 21784 11336 21790 11348
rect 22094 11336 22100 11348
rect 21784 11308 22100 11336
rect 21784 11296 21790 11308
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 23845 11339 23903 11345
rect 23845 11336 23857 11339
rect 23532 11308 23857 11336
rect 23532 11296 23538 11308
rect 23845 11305 23857 11308
rect 23891 11305 23903 11339
rect 23845 11299 23903 11305
rect 23937 11339 23995 11345
rect 23937 11305 23949 11339
rect 23983 11336 23995 11339
rect 24026 11336 24032 11348
rect 23983 11308 24032 11336
rect 23983 11305 23995 11308
rect 23937 11299 23995 11305
rect 15746 11268 15752 11280
rect 14936 11240 15752 11268
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 16301 11271 16359 11277
rect 16301 11237 16313 11271
rect 16347 11268 16359 11271
rect 18340 11268 18368 11296
rect 20625 11271 20683 11277
rect 20625 11268 20637 11271
rect 16347 11240 20637 11268
rect 16347 11237 16359 11240
rect 16301 11231 16359 11237
rect 20625 11237 20637 11240
rect 20671 11268 20683 11271
rect 20990 11268 20996 11280
rect 20671 11240 20996 11268
rect 20671 11237 20683 11240
rect 20625 11231 20683 11237
rect 20990 11228 20996 11240
rect 21048 11228 21054 11280
rect 22462 11268 22468 11280
rect 21100 11240 22468 11268
rect 10962 11209 10968 11212
rect 10956 11200 10968 11209
rect 10742 11172 10824 11200
rect 10923 11172 10968 11200
rect 10742 11169 10754 11172
rect 10696 11163 10754 11169
rect 10956 11163 10968 11172
rect 10962 11160 10968 11163
rect 11020 11160 11026 11212
rect 13262 11160 13268 11212
rect 13320 11160 13326 11212
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 13814 11200 13820 11212
rect 13412 11172 13820 11200
rect 13412 11160 13418 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16114 11200 16120 11212
rect 15703 11172 16120 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17586 11200 17592 11212
rect 17175 11172 17592 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 18380 11172 18521 11200
rect 18380 11160 18386 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18748 11172 19073 11200
rect 18748 11160 18754 11172
rect 19061 11169 19073 11172
rect 19107 11200 19119 11203
rect 19518 11200 19524 11212
rect 19107 11172 19524 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 19702 11200 19708 11212
rect 19615 11172 19708 11200
rect 19702 11160 19708 11172
rect 19760 11200 19766 11212
rect 21100 11200 21128 11240
rect 22462 11228 22468 11240
rect 22520 11228 22526 11280
rect 22186 11200 22192 11212
rect 19760 11172 21128 11200
rect 22147 11172 22192 11200
rect 19760 11160 19766 11172
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 22281 11203 22339 11209
rect 22281 11169 22293 11203
rect 22327 11200 22339 11203
rect 22646 11200 22652 11212
rect 22327 11172 22652 11200
rect 22327 11169 22339 11172
rect 22281 11163 22339 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 5166 11132 5172 11144
rect 5127 11104 5172 11132
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5592 11104 6132 11132
rect 5592 11092 5598 11104
rect 4580 11036 5028 11064
rect 4580 11024 4586 11036
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 6104 11073 6132 11104
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6512 11104 6653 11132
rect 6512 11092 6518 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7374 11132 7380 11144
rect 6779 11104 7380 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5132 11036 5641 11064
rect 5132 11024 5138 11036
rect 5629 11033 5641 11036
rect 5675 11033 5687 11067
rect 5629 11027 5687 11033
rect 6089 11067 6147 11073
rect 6089 11033 6101 11067
rect 6135 11064 6147 11067
rect 6748 11064 6776 11095
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 8110 11132 8116 11144
rect 7708 11104 8116 11132
rect 7708 11092 7714 11104
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 8168 11104 8217 11132
rect 8168 11092 8174 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 13722 11132 13728 11144
rect 12943 11104 13728 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 6135 11036 6776 11064
rect 6135 11033 6147 11036
rect 6089 11027 6147 11033
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 6880 11036 7757 11064
rect 6880 11024 6886 11036
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 8312 11064 8340 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 7745 11027 7803 11033
rect 7852 11036 8340 11064
rect 7852 11008 7880 11036
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 10192 11036 10241 11064
rect 10192 11024 10198 11036
rect 10229 11033 10241 11036
rect 10275 11033 10287 11067
rect 10229 11027 10287 11033
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 11756 11036 12848 11064
rect 11756 11024 11762 11036
rect 12820 11008 12848 11036
rect 4430 10996 4436 11008
rect 4080 10968 4436 10996
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10996 7711 10999
rect 7834 10996 7840 11008
rect 7699 10968 7840 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 9030 10996 9036 11008
rect 8991 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 12066 10996 12072 11008
rect 9732 10968 12072 10996
rect 9732 10956 9738 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13924 10996 13952 11095
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14366 11132 14372 11144
rect 14056 11104 14372 11132
rect 14056 11092 14062 11104
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14424 11104 14473 11132
rect 14424 11092 14430 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 16632 11104 17325 11132
rect 16632 11092 16638 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20438 11132 20444 11144
rect 19843 11104 20444 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 15470 11024 15476 11076
rect 15528 11064 15534 11076
rect 15841 11067 15899 11073
rect 15841 11064 15853 11067
rect 15528 11036 15853 11064
rect 15528 11024 15534 11036
rect 15841 11033 15853 11036
rect 15887 11033 15899 11067
rect 15841 11027 15899 11033
rect 19426 11024 19432 11076
rect 19484 11064 19490 11076
rect 19812 11064 19840 11095
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 22462 11132 22468 11144
rect 21775 11104 22468 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22462 11092 22468 11104
rect 22520 11132 22526 11144
rect 22848 11132 22876 11296
rect 23385 11271 23443 11277
rect 23385 11237 23397 11271
rect 23431 11268 23443 11271
rect 23952 11268 23980 11299
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24489 11339 24547 11345
rect 24489 11336 24501 11339
rect 24176 11308 24501 11336
rect 24176 11296 24182 11308
rect 24489 11305 24501 11308
rect 24535 11305 24547 11339
rect 24489 11299 24547 11305
rect 25225 11339 25283 11345
rect 25225 11305 25237 11339
rect 25271 11336 25283 11339
rect 25406 11336 25412 11348
rect 25271 11308 25412 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 24946 11268 24952 11280
rect 23431 11240 23980 11268
rect 24907 11240 24952 11268
rect 23431 11237 23443 11240
rect 23385 11231 23443 11237
rect 24946 11228 24952 11240
rect 25004 11268 25010 11280
rect 25682 11268 25688 11280
rect 25004 11240 25688 11268
rect 25004 11228 25010 11240
rect 25682 11228 25688 11240
rect 25740 11228 25746 11280
rect 25041 11203 25099 11209
rect 25041 11169 25053 11203
rect 25087 11200 25099 11203
rect 25590 11200 25596 11212
rect 25087 11172 25596 11200
rect 25087 11169 25099 11172
rect 25041 11163 25099 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 22520 11104 22876 11132
rect 22520 11092 22526 11104
rect 23934 11092 23940 11144
rect 23992 11132 23998 11144
rect 24121 11135 24179 11141
rect 24121 11132 24133 11135
rect 23992 11104 24133 11132
rect 23992 11092 23998 11104
rect 24121 11101 24133 11104
rect 24167 11132 24179 11135
rect 24302 11132 24308 11144
rect 24167 11104 24308 11132
rect 24167 11101 24179 11104
rect 24121 11095 24179 11101
rect 24302 11092 24308 11104
rect 24360 11092 24366 11144
rect 21818 11064 21824 11076
rect 19484 11036 19840 11064
rect 21779 11036 21824 11064
rect 19484 11024 19490 11036
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 23477 11067 23535 11073
rect 23477 11033 23489 11067
rect 23523 11064 23535 11067
rect 23750 11064 23756 11076
rect 23523 11036 23756 11064
rect 23523 11033 23535 11036
rect 23477 11027 23535 11033
rect 23750 11024 23756 11036
rect 23808 11024 23814 11076
rect 14366 10996 14372 11008
rect 12860 10968 14372 10996
rect 12860 10956 12866 10968
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16669 10999 16727 11005
rect 16669 10965 16681 10999
rect 16715 10996 16727 10999
rect 16942 10996 16948 11008
rect 16715 10968 16948 10996
rect 16715 10965 16727 10968
rect 16669 10959 16727 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 20346 10956 20352 11008
rect 20404 10996 20410 11008
rect 25038 10996 25044 11008
rect 20404 10968 25044 10996
rect 20404 10956 20410 10968
rect 25038 10956 25044 10968
rect 25096 10956 25102 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2222 10792 2228 10804
rect 1811 10764 2228 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2222 10752 2228 10764
rect 2280 10792 2286 10804
rect 4062 10792 4068 10804
rect 2280 10764 3280 10792
rect 4023 10764 4068 10792
rect 2280 10752 2286 10764
rect 3252 10733 3280 10764
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4890 10792 4896 10804
rect 4479 10764 4896 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4890 10752 4896 10764
rect 4948 10792 4954 10804
rect 5166 10792 5172 10804
rect 4948 10764 5172 10792
rect 4948 10752 4954 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5905 10795 5963 10801
rect 5905 10792 5917 10795
rect 5500 10764 5917 10792
rect 5500 10752 5506 10764
rect 5905 10761 5917 10764
rect 5951 10761 5963 10795
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 5905 10755 5963 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9306 10792 9312 10804
rect 9263 10764 9312 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 10042 10792 10048 10804
rect 10003 10764 10048 10792
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10318 10792 10324 10804
rect 10279 10764 10324 10792
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 12066 10792 12072 10804
rect 11979 10764 12072 10792
rect 12066 10752 12072 10764
rect 12124 10792 12130 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12124 10764 12173 10792
rect 12124 10752 12130 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 14826 10792 14832 10804
rect 14787 10764 14832 10792
rect 12161 10755 12219 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 15378 10792 15384 10804
rect 15335 10764 15384 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 16482 10792 16488 10804
rect 16439 10764 16488 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 17218 10792 17224 10804
rect 16807 10764 17224 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 19245 10795 19303 10801
rect 19245 10761 19257 10795
rect 19291 10792 19303 10795
rect 19426 10792 19432 10804
rect 19291 10764 19432 10792
rect 19291 10761 19303 10764
rect 19245 10755 19303 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 21082 10792 21088 10804
rect 19576 10764 20668 10792
rect 21043 10764 21088 10792
rect 19576 10752 19582 10764
rect 3237 10727 3295 10733
rect 3237 10693 3249 10727
rect 3283 10724 3295 10727
rect 3970 10724 3976 10736
rect 3283 10696 3976 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 6638 10724 6644 10736
rect 6599 10696 6644 10724
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 1854 10656 1860 10668
rect 1815 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 4430 10616 4436 10668
rect 4488 10656 4494 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4488 10628 4537 10656
rect 4488 10616 4494 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 4525 10619 4583 10625
rect 9048 10628 9689 10656
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4792 10591 4850 10597
rect 4792 10588 4804 10591
rect 4672 10560 4804 10588
rect 4672 10548 4678 10560
rect 4792 10557 4804 10560
rect 4838 10588 4850 10591
rect 5350 10588 5356 10600
rect 4838 10560 5356 10588
rect 4838 10557 4850 10560
rect 4792 10551 4850 10557
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 7374 10588 7380 10600
rect 6871 10560 7380 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 7374 10548 7380 10560
rect 7432 10588 7438 10600
rect 8110 10588 8116 10600
rect 7432 10560 8116 10588
rect 7432 10548 7438 10560
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 9048 10597 9076 10628
rect 9677 10625 9689 10628
rect 9723 10656 9735 10659
rect 10226 10656 10232 10668
rect 9723 10628 10232 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10336 10656 10364 10752
rect 10778 10684 10784 10736
rect 10836 10724 10842 10736
rect 10836 10696 11192 10724
rect 10836 10684 10842 10696
rect 11164 10665 11192 10696
rect 11606 10684 11612 10736
rect 11664 10724 11670 10736
rect 17494 10724 17500 10736
rect 11664 10696 17500 10724
rect 11664 10684 11670 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 20640 10724 20668 10764
rect 21082 10752 21088 10764
rect 21140 10752 21146 10804
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 20640 10696 21588 10724
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10336 10628 10977 10656
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 12526 10656 12532 10668
rect 11195 10628 12532 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 13446 10616 13452 10668
rect 13504 10656 13510 10668
rect 13998 10656 14004 10668
rect 13504 10628 14004 10656
rect 13504 10616 13510 10628
rect 13998 10616 14004 10628
rect 14056 10656 14062 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 14056 10628 14289 10656
rect 14056 10616 14062 10628
rect 14277 10625 14289 10628
rect 14323 10656 14335 10659
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14323 10628 15117 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15620 10628 15853 10656
rect 15620 10616 15626 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17368 10628 17877 10656
rect 17368 10616 17374 10628
rect 17865 10625 17877 10628
rect 17911 10656 17923 10659
rect 18690 10656 18696 10668
rect 17911 10628 18696 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8260 10560 9045 10588
rect 8260 10548 8266 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10100 10560 10885 10588
rect 10100 10548 10106 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10588 12127 10591
rect 12621 10591 12679 10597
rect 12621 10588 12633 10591
rect 12115 10560 12633 10588
rect 12115 10557 12127 10560
rect 12069 10551 12127 10557
rect 12621 10557 12633 10560
rect 12667 10557 12679 10591
rect 12621 10551 12679 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14826 10588 14832 10600
rect 14139 10560 14832 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15654 10588 15660 10600
rect 15615 10560 15660 10588
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 16942 10588 16948 10600
rect 16899 10560 16948 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18104 10560 18429 10588
rect 18104 10548 18110 10560
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 19058 10588 19064 10600
rect 18564 10560 19064 10588
rect 18564 10548 18570 10560
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20530 10588 20536 10600
rect 19751 10560 20536 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 21560 10597 21588 10696
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 22557 10659 22615 10665
rect 22557 10656 22569 10659
rect 22520 10628 22569 10656
rect 22520 10616 22526 10628
rect 22557 10625 22569 10628
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 23566 10616 23572 10668
rect 23624 10616 23630 10668
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10588 21603 10591
rect 23584 10588 23612 10616
rect 21591 10560 23612 10588
rect 23937 10591 23995 10597
rect 21591 10557 21603 10560
rect 21545 10551 21603 10557
rect 2124 10523 2182 10529
rect 2124 10489 2136 10523
rect 2170 10520 2182 10523
rect 2682 10520 2688 10532
rect 2170 10492 2688 10520
rect 2170 10489 2182 10492
rect 2124 10483 2182 10489
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 3418 10520 3424 10532
rect 2740 10492 3424 10520
rect 2740 10480 2746 10492
rect 3418 10480 3424 10492
rect 3476 10520 3482 10532
rect 3513 10523 3571 10529
rect 3513 10520 3525 10523
rect 3476 10492 3525 10520
rect 3476 10480 3482 10492
rect 3513 10489 3525 10492
rect 3559 10489 3571 10523
rect 3513 10483 3571 10489
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6972 10492 7082 10520
rect 6972 10480 6978 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 11146 10520 11152 10532
rect 7070 10483 7128 10489
rect 10060 10492 11152 10520
rect 10060 10464 10088 10492
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 15286 10480 15292 10532
rect 15344 10520 15350 10532
rect 17402 10520 17408 10532
rect 15344 10492 17408 10520
rect 15344 10480 15350 10492
rect 17402 10480 17408 10492
rect 17460 10480 17466 10532
rect 19978 10529 19984 10532
rect 19613 10523 19671 10529
rect 19613 10489 19625 10523
rect 19659 10520 19671 10523
rect 19972 10520 19984 10529
rect 19659 10492 19984 10520
rect 19659 10489 19671 10492
rect 19613 10483 19671 10489
rect 19972 10483 19984 10492
rect 19978 10480 19984 10483
rect 20036 10480 20042 10532
rect 22480 10529 22508 10560
rect 23937 10557 23949 10591
rect 23983 10588 23995 10591
rect 24946 10588 24952 10600
rect 23983 10560 24952 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24946 10548 24952 10560
rect 25004 10588 25010 10600
rect 25961 10591 26019 10597
rect 25961 10588 25973 10591
rect 25004 10560 25973 10588
rect 25004 10548 25010 10560
rect 25961 10557 25973 10560
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 22373 10523 22431 10529
rect 22373 10520 22385 10523
rect 21836 10492 22385 10520
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6454 10452 6460 10464
rect 6319 10424 6460 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 7834 10412 7840 10464
rect 7892 10452 7898 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7892 10424 8217 10452
rect 7892 10412 7898 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 10686 10452 10692 10464
rect 10551 10424 10692 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11112 10424 11621 10452
rect 11112 10412 11118 10424
rect 11609 10421 11621 10424
rect 11655 10452 11667 10455
rect 11974 10452 11980 10464
rect 11655 10424 11980 10452
rect 11655 10421 11667 10424
rect 11609 10415 11667 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 13412 10424 13461 10452
rect 13412 10412 13418 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13449 10415 13507 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 15838 10452 15844 10464
rect 15795 10424 15844 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 17126 10452 17132 10464
rect 17083 10424 17132 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17497 10455 17555 10461
rect 17497 10421 17509 10455
rect 17543 10452 17555 10455
rect 17586 10452 17592 10464
rect 17543 10424 17592 10452
rect 17543 10421 17555 10424
rect 17497 10415 17555 10421
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17920 10424 18061 10452
rect 17920 10412 17926 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 21836 10461 21864 10492
rect 22373 10489 22385 10492
rect 22419 10489 22431 10523
rect 22373 10483 22431 10489
rect 22465 10523 22523 10529
rect 22465 10489 22477 10523
rect 22511 10489 22523 10523
rect 22465 10483 22523 10489
rect 22830 10480 22836 10532
rect 22888 10520 22894 10532
rect 23566 10520 23572 10532
rect 22888 10492 23572 10520
rect 22888 10480 22894 10492
rect 23566 10480 23572 10492
rect 23624 10480 23630 10532
rect 24210 10529 24216 10532
rect 24204 10483 24216 10529
rect 24268 10520 24274 10532
rect 24268 10492 24304 10520
rect 24210 10480 24216 10483
rect 24268 10480 24274 10492
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 21784 10424 21833 10452
rect 21784 10412 21790 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21968 10424 22017 10452
rect 21968 10412 21974 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22646 10412 22652 10464
rect 22704 10452 22710 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22704 10424 23029 10452
rect 22704 10412 22710 10424
rect 23017 10421 23029 10424
rect 23063 10421 23075 10455
rect 25314 10452 25320 10464
rect 25275 10424 25320 10452
rect 23017 10415 23075 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2740 10220 3065 10248
rect 2740 10208 2746 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 4614 10248 4620 10260
rect 4575 10220 4620 10248
rect 3053 10211 3111 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 4948 10220 6285 10248
rect 4948 10208 4954 10220
rect 6273 10217 6285 10220
rect 6319 10248 6331 10251
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6319 10220 6837 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6825 10217 6837 10220
rect 6871 10248 6883 10251
rect 6914 10248 6920 10260
rect 6871 10220 6920 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7098 10248 7104 10260
rect 7059 10220 7104 10248
rect 7098 10208 7104 10220
rect 7156 10248 7162 10260
rect 9030 10248 9036 10260
rect 7156 10220 9036 10248
rect 7156 10208 7162 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10778 10248 10784 10260
rect 10551 10220 10784 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 12115 10220 14105 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 14366 10248 14372 10260
rect 14323 10220 14372 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 15654 10248 15660 10260
rect 14783 10220 15660 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18506 10248 18512 10260
rect 18187 10220 18512 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 19242 10248 19248 10260
rect 18831 10220 19248 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 19705 10251 19763 10257
rect 19705 10217 19717 10251
rect 19751 10248 19763 10251
rect 20162 10248 20168 10260
rect 19751 10220 20168 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 22002 10248 22008 10260
rect 20763 10220 22008 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22244 10220 22293 10248
rect 22244 10208 22250 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 23201 10251 23259 10257
rect 23201 10248 23213 10251
rect 22704 10220 23213 10248
rect 22704 10208 22710 10220
rect 23201 10217 23213 10220
rect 23247 10248 23259 10251
rect 23290 10248 23296 10260
rect 23247 10220 23296 10248
rect 23247 10217 23259 10220
rect 23201 10211 23259 10217
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 23934 10248 23940 10260
rect 23895 10220 23940 10248
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 24210 10248 24216 10260
rect 24171 10220 24216 10248
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 24857 10251 24915 10257
rect 24857 10248 24869 10251
rect 24360 10220 24869 10248
rect 24360 10208 24366 10220
rect 24857 10217 24869 10220
rect 24903 10248 24915 10251
rect 25222 10248 25228 10260
rect 24903 10220 25228 10248
rect 24903 10217 24915 10220
rect 24857 10211 24915 10217
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 25774 10248 25780 10260
rect 25735 10220 25780 10248
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 1854 10140 1860 10192
rect 1912 10140 1918 10192
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 3697 10183 3755 10189
rect 3697 10180 3709 10183
rect 2832 10152 3709 10180
rect 2832 10140 2838 10152
rect 3697 10149 3709 10152
rect 3743 10149 3755 10183
rect 3697 10143 3755 10149
rect 5160 10183 5218 10189
rect 5160 10149 5172 10183
rect 5206 10180 5218 10183
rect 5442 10180 5448 10192
rect 5206 10152 5448 10180
rect 5206 10149 5218 10152
rect 5160 10143 5218 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 14458 10180 14464 10192
rect 10100 10152 14464 10180
rect 10100 10140 10106 10152
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1872 10112 1900 10140
rect 1719 10084 1900 10112
rect 1940 10115 1998 10121
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 1940 10081 1952 10115
rect 1986 10112 1998 10115
rect 2958 10112 2964 10124
rect 1986 10084 2964 10112
rect 1986 10081 1998 10084
rect 1940 10075 1998 10081
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3510 10112 3516 10124
rect 3467 10084 3516 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4488 10084 4905 10112
rect 4488 10072 4494 10084
rect 4893 10081 4905 10084
rect 4939 10112 4951 10115
rect 7282 10112 7288 10124
rect 4939 10084 6592 10112
rect 7243 10084 7288 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 6564 10044 6592 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7650 10121 7656 10124
rect 7644 10112 7656 10121
rect 7611 10084 7656 10112
rect 7644 10075 7656 10084
rect 7650 10072 7656 10075
rect 7708 10072 7714 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10870 10121 10876 10124
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 10008 10084 10609 10112
rect 10008 10072 10014 10084
rect 10597 10081 10609 10084
rect 10643 10081 10655 10115
rect 10864 10112 10876 10121
rect 10831 10084 10876 10112
rect 10597 10075 10655 10081
rect 10864 10075 10876 10084
rect 10870 10072 10876 10075
rect 10928 10072 10934 10124
rect 12066 10072 12072 10124
rect 12124 10112 12130 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12124 10084 13185 10112
rect 12124 10072 12130 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 15948 10112 15976 10208
rect 16660 10183 16718 10189
rect 16660 10149 16672 10183
rect 16706 10180 16718 10183
rect 17310 10180 17316 10192
rect 16706 10152 17316 10180
rect 16706 10149 16718 10152
rect 16660 10143 16718 10149
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 17770 10180 17776 10192
rect 17552 10152 17776 10180
rect 17552 10140 17558 10152
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 18966 10140 18972 10192
rect 19024 10180 19030 10192
rect 19061 10183 19119 10189
rect 19061 10180 19073 10183
rect 19024 10152 19073 10180
rect 19024 10140 19030 10152
rect 19061 10149 19073 10152
rect 19107 10149 19119 10183
rect 19061 10143 19119 10149
rect 22922 10140 22928 10192
rect 22980 10180 22986 10192
rect 24228 10180 24256 10208
rect 22980 10152 23336 10180
rect 24228 10152 24992 10180
rect 22980 10140 22986 10152
rect 16390 10112 16396 10124
rect 15335 10084 15976 10112
rect 16351 10084 16396 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 20346 10112 20352 10124
rect 19659 10084 20352 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 21174 10072 21180 10124
rect 21232 10072 21238 10124
rect 21358 10072 21364 10124
rect 21416 10112 21422 10124
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21416 10084 21649 10112
rect 21416 10072 21422 10084
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 22462 10112 22468 10124
rect 21637 10075 21695 10081
rect 21928 10084 22468 10112
rect 7374 10044 7380 10056
rect 6564 10016 7380 10044
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 12676 10016 13277 10044
rect 12676 10004 12682 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10044 15163 10047
rect 15838 10044 15844 10056
rect 15151 10016 15844 10044
rect 15151 10013 15163 10016
rect 15105 10007 15163 10013
rect 8754 9976 8760 9988
rect 8715 9948 8760 9976
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 12069 9979 12127 9985
rect 12069 9976 12081 9979
rect 9732 9948 10640 9976
rect 9732 9936 9738 9948
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 3142 9908 3148 9920
rect 2372 9880 3148 9908
rect 2372 9868 2378 9880
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 8570 9908 8576 9920
rect 4856 9880 8576 9908
rect 4856 9868 4862 9880
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 9398 9908 9404 9920
rect 9359 9880 9404 9908
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10042 9908 10048 9920
rect 9999 9880 10048 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10612 9908 10640 9948
rect 11808 9948 12081 9976
rect 11808 9908 11836 9948
rect 12069 9945 12081 9948
rect 12115 9945 12127 9979
rect 12069 9939 12127 9945
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 12805 9979 12863 9985
rect 12805 9976 12817 9979
rect 12400 9948 12817 9976
rect 12400 9936 12406 9948
rect 12805 9945 12817 9948
rect 12851 9945 12863 9979
rect 12805 9939 12863 9945
rect 11974 9908 11980 9920
rect 10612 9880 11836 9908
rect 11935 9880 11980 9908
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12253 9911 12311 9917
rect 12253 9908 12265 9911
rect 12216 9880 12265 9908
rect 12216 9868 12222 9880
rect 12253 9877 12265 9880
rect 12299 9877 12311 9911
rect 12253 9871 12311 9877
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12584 9880 12633 9908
rect 12584 9868 12590 9880
rect 12621 9877 12633 9880
rect 12667 9908 12679 9911
rect 13372 9908 13400 10007
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19576 10016 19809 10044
rect 19576 10004 19582 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19978 10004 19984 10056
rect 20036 10044 20042 10056
rect 21192 10044 21220 10072
rect 20036 10016 21220 10044
rect 20036 10004 20042 10016
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 21928 10053 21956 10084
rect 22462 10072 22468 10084
rect 22520 10112 22526 10124
rect 22649 10115 22707 10121
rect 22649 10112 22661 10115
rect 22520 10084 22661 10112
rect 22520 10072 22526 10084
rect 22649 10081 22661 10084
rect 22695 10112 22707 10115
rect 23308 10112 23336 10152
rect 22695 10084 23244 10112
rect 23308 10084 23428 10112
rect 22695 10081 22707 10084
rect 22649 10075 22707 10081
rect 21729 10047 21787 10053
rect 21729 10044 21741 10047
rect 21324 10016 21741 10044
rect 21324 10004 21330 10016
rect 21729 10013 21741 10016
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 14093 9979 14151 9985
rect 14093 9945 14105 9979
rect 14139 9976 14151 9979
rect 15286 9976 15292 9988
rect 14139 9948 15292 9976
rect 14139 9945 14151 9948
rect 14093 9939 14151 9945
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 21177 9979 21235 9985
rect 21177 9945 21189 9979
rect 21223 9976 21235 9979
rect 21928 9976 21956 10007
rect 21223 9948 21956 9976
rect 21223 9945 21235 9948
rect 21177 9939 21235 9945
rect 12667 9880 13400 9908
rect 13909 9911 13967 9917
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 13909 9877 13921 9911
rect 13955 9908 13967 9911
rect 14182 9908 14188 9920
rect 13955 9880 14188 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 14182 9868 14188 9880
rect 14240 9908 14246 9920
rect 15378 9908 15384 9920
rect 14240 9880 15384 9908
rect 14240 9868 14246 9880
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 15473 9911 15531 9917
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 15930 9908 15936 9920
rect 15519 9880 15936 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16209 9911 16267 9917
rect 16209 9908 16221 9911
rect 16172 9880 16221 9908
rect 16172 9868 16178 9880
rect 16209 9877 16221 9880
rect 16255 9877 16267 9911
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 16209 9871 16267 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 19242 9908 19248 9920
rect 19203 9880 19248 9908
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 20254 9908 20260 9920
rect 20215 9880 20260 9908
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 21269 9911 21327 9917
rect 21269 9877 21281 9911
rect 21315 9908 21327 9911
rect 21634 9908 21640 9920
rect 21315 9880 21640 9908
rect 21315 9877 21327 9880
rect 21269 9871 21327 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 22830 9908 22836 9920
rect 22791 9880 22836 9908
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 23216 9908 23244 10084
rect 23400 10053 23428 10084
rect 23934 10072 23940 10124
rect 23992 10112 23998 10124
rect 24765 10115 24823 10121
rect 24765 10112 24777 10115
rect 23992 10084 24777 10112
rect 23992 10072 23998 10084
rect 24765 10081 24777 10084
rect 24811 10112 24823 10115
rect 24854 10112 24860 10124
rect 24811 10084 24860 10112
rect 24811 10081 24823 10084
rect 24765 10075 24823 10081
rect 24854 10072 24860 10084
rect 24912 10072 24918 10124
rect 24964 10056 24992 10152
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10013 23351 10047
rect 23293 10007 23351 10013
rect 23385 10047 23443 10053
rect 23385 10013 23397 10047
rect 23431 10013 23443 10047
rect 23385 10007 23443 10013
rect 23308 9976 23336 10007
rect 24946 10004 24952 10056
rect 25004 10044 25010 10056
rect 25004 10016 25097 10044
rect 25004 10004 25010 10016
rect 23308 9948 24440 9976
rect 24210 9908 24216 9920
rect 23216 9880 24216 9908
rect 24210 9868 24216 9880
rect 24268 9868 24274 9920
rect 24412 9917 24440 9948
rect 24397 9911 24455 9917
rect 24397 9877 24409 9911
rect 24443 9908 24455 9911
rect 24762 9908 24768 9920
rect 24443 9880 24768 9908
rect 24443 9877 24455 9880
rect 24397 9871 24455 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 25501 9911 25559 9917
rect 25501 9877 25513 9911
rect 25547 9908 25559 9911
rect 25590 9908 25596 9920
rect 25547 9880 25596 9908
rect 25547 9877 25559 9880
rect 25501 9871 25559 9877
rect 25590 9868 25596 9880
rect 25648 9868 25654 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 5721 9707 5779 9713
rect 5721 9704 5733 9707
rect 5500 9676 5733 9704
rect 5500 9664 5506 9676
rect 5721 9673 5733 9676
rect 5767 9673 5779 9707
rect 7282 9704 7288 9716
rect 5721 9667 5779 9673
rect 6840 9676 7288 9704
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9636 1639 9639
rect 1946 9636 1952 9648
rect 1627 9608 1952 9636
rect 1627 9605 1639 9608
rect 1581 9599 1639 9605
rect 1946 9596 1952 9608
rect 2004 9596 2010 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4580 9608 4721 9636
rect 4580 9596 4586 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 4709 9599 4767 9605
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9568 2194 9580
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2188 9540 3801 9568
rect 2188 9528 2194 9540
rect 3789 9537 3801 9540
rect 3835 9568 3847 9571
rect 3878 9568 3884 9580
rect 3835 9540 3884 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4663 9540 5365 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 5353 9537 5365 9540
rect 5399 9568 5411 9571
rect 5460 9568 5488 9664
rect 6641 9639 6699 9645
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 6840 9636 6868 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 12066 9664 12072 9716
rect 12124 9664 12130 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 12676 9676 13001 9704
rect 12676 9664 12682 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 12989 9667 13047 9673
rect 16945 9707 17003 9713
rect 16945 9673 16957 9707
rect 16991 9704 17003 9707
rect 17310 9704 17316 9716
rect 16991 9676 17316 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 19797 9707 19855 9713
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 20162 9704 20168 9716
rect 19843 9676 20168 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 23934 9664 23940 9716
rect 23992 9704 23998 9716
rect 24026 9704 24032 9716
rect 23992 9676 24032 9704
rect 23992 9664 23998 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 24670 9664 24676 9716
rect 24728 9704 24734 9716
rect 25222 9704 25228 9716
rect 24728 9676 25228 9704
rect 24728 9664 24734 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 25774 9664 25780 9716
rect 25832 9704 25838 9716
rect 26145 9707 26203 9713
rect 26145 9704 26157 9707
rect 25832 9676 26157 9704
rect 25832 9664 25838 9676
rect 26145 9673 26157 9676
rect 26191 9673 26203 9707
rect 26145 9667 26203 9673
rect 6687 9608 6868 9636
rect 10229 9639 10287 9645
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 10229 9605 10241 9639
rect 10275 9636 10287 9639
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 10275 9608 10609 9636
rect 10275 9605 10287 9608
rect 10229 9599 10287 9605
rect 10597 9605 10609 9608
rect 10643 9636 10655 9639
rect 10870 9636 10876 9648
rect 10643 9608 10876 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 10870 9596 10876 9608
rect 10928 9636 10934 9648
rect 12084 9636 12112 9664
rect 12158 9636 12164 9648
rect 10928 9608 11376 9636
rect 12084 9608 12164 9636
rect 10928 9596 10934 9608
rect 7558 9568 7564 9580
rect 5399 9540 5488 9568
rect 7519 9540 7564 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 11348 9577 11376 9608
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13170 9636 13176 9648
rect 12860 9608 13176 9636
rect 12860 9596 12866 9608
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 14458 9636 14464 9648
rect 14419 9608 14464 9636
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19484 9608 20269 9636
rect 19484 9596 19490 9608
rect 20257 9605 20269 9608
rect 20303 9605 20315 9639
rect 20257 9599 20315 9605
rect 24946 9596 24952 9648
rect 25004 9636 25010 9648
rect 25133 9639 25191 9645
rect 25133 9636 25145 9639
rect 25004 9608 25145 9636
rect 25004 9596 25010 9608
rect 25133 9605 25145 9608
rect 25179 9636 25191 9639
rect 25409 9639 25467 9645
rect 25409 9636 25421 9639
rect 25179 9608 25421 9636
rect 25179 9605 25191 9608
rect 25133 9599 25191 9605
rect 25409 9605 25421 9608
rect 25455 9605 25467 9639
rect 25409 9599 25467 9605
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 11333 9571 11391 9577
rect 9907 9540 11192 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3016 9472 4169 9500
rect 3016 9460 3022 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 11164 9509 11192 9540
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 12066 9568 12072 9580
rect 11379 9540 12072 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 15519 9540 15700 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 10744 9472 11069 9500
rect 10744 9460 10750 9472
rect 11057 9469 11069 9472
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 12342 9500 12348 9512
rect 11195 9472 12348 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 13170 9500 13176 9512
rect 12492 9472 13176 9500
rect 12492 9460 12498 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15672 9500 15700 9540
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 18012 9540 18061 9568
rect 18012 9528 18018 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 20898 9568 20904 9580
rect 20859 9540 20904 9568
rect 18049 9531 18107 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 22830 9568 22836 9580
rect 22695 9540 22836 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 24854 9528 24860 9580
rect 24912 9568 24918 9580
rect 25777 9571 25835 9577
rect 25777 9568 25789 9571
rect 24912 9540 25789 9568
rect 24912 9528 24918 9540
rect 25777 9537 25789 9540
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 15832 9503 15890 9509
rect 15832 9500 15844 9503
rect 15672 9472 15844 9500
rect 15565 9463 15623 9469
rect 15832 9469 15844 9472
rect 15878 9500 15890 9503
rect 16206 9500 16212 9512
rect 15878 9472 16212 9500
rect 15878 9469 15890 9472
rect 15832 9463 15890 9469
rect 1949 9435 2007 9441
rect 1949 9401 1961 9435
rect 1995 9432 2007 9435
rect 3053 9435 3111 9441
rect 1995 9404 2728 9432
rect 1995 9401 2007 9404
rect 1949 9395 2007 9401
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2700 9373 2728 9404
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 3099 9404 3648 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 3620 9376 3648 9404
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4948 9404 5089 9432
rect 4948 9392 4954 9404
rect 5077 9401 5089 9404
rect 5123 9432 5135 9435
rect 6089 9435 6147 9441
rect 6089 9432 6101 9435
rect 5123 9404 6101 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 6089 9401 6101 9404
rect 6135 9401 6147 9435
rect 6089 9395 6147 9401
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 7101 9435 7159 9441
rect 7101 9432 7113 9435
rect 6420 9404 7113 9432
rect 6420 9392 6426 9404
rect 7101 9401 7113 9404
rect 7147 9432 7159 9435
rect 7828 9435 7886 9441
rect 7828 9432 7840 9435
rect 7147 9404 7840 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7828 9401 7840 9404
rect 7874 9432 7886 9435
rect 8662 9432 8668 9444
rect 7874 9404 8668 9432
rect 7874 9401 7886 9404
rect 7828 9395 7886 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 12158 9432 12164 9444
rect 12119 9404 12164 9432
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 15580 9432 15608 9463
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 20622 9500 20628 9512
rect 19392 9472 20628 9500
rect 19392 9460 19398 9472
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 22152 9472 22385 9500
rect 22152 9460 22158 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 23753 9503 23811 9509
rect 23753 9500 23765 9503
rect 23440 9472 23765 9500
rect 23440 9460 23446 9472
rect 23753 9469 23765 9472
rect 23799 9500 23811 9503
rect 25590 9500 25596 9512
rect 23799 9472 25596 9500
rect 23799 9469 23811 9472
rect 23753 9463 23811 9469
rect 25590 9460 25596 9472
rect 25648 9460 25654 9512
rect 16390 9432 16396 9444
rect 15580 9404 16396 9432
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 17788 9404 18306 9432
rect 17788 9376 17816 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 20254 9432 20260 9444
rect 18294 9395 18352 9401
rect 19352 9404 20260 9432
rect 19352 9376 19380 9404
rect 20254 9392 20260 9404
rect 20312 9432 20318 9444
rect 20717 9435 20775 9441
rect 20717 9432 20729 9435
rect 20312 9404 20729 9432
rect 20312 9392 20318 9404
rect 20717 9401 20729 9404
rect 20763 9401 20775 9435
rect 20717 9395 20775 9401
rect 23290 9392 23296 9444
rect 23348 9392 23354 9444
rect 23477 9435 23535 9441
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 23934 9432 23940 9444
rect 23523 9404 23940 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 23934 9392 23940 9404
rect 23992 9441 23998 9444
rect 23992 9435 24056 9441
rect 23992 9401 24010 9435
rect 24044 9401 24056 9435
rect 23992 9395 24056 9401
rect 23992 9392 23998 9395
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 2866 9364 2872 9376
rect 2731 9336 2872 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3142 9364 3148 9376
rect 3103 9336 3148 9364
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 3476 9336 3525 9364
rect 3476 9324 3482 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 5169 9367 5227 9373
rect 3660 9336 3705 9364
rect 3660 9324 3666 9336
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5442 9364 5448 9376
rect 5215 9336 5448 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9364 7527 9367
rect 7650 9364 7656 9376
rect 7515 9336 7656 9364
rect 7515 9333 7527 9336
rect 7469 9327 7527 9333
rect 7650 9324 7656 9336
rect 7708 9364 7714 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 7708 9336 8953 9364
rect 7708 9324 7714 9336
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 8941 9327 8999 9333
rect 9309 9367 9367 9373
rect 9309 9333 9321 9367
rect 9355 9364 9367 9367
rect 9398 9364 9404 9376
rect 9355 9336 9404 9364
rect 9355 9333 9367 9336
rect 9309 9327 9367 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10778 9364 10784 9376
rect 10735 9336 10784 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11790 9364 11796 9376
rect 11112 9336 11796 9364
rect 11112 9324 11118 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12943 9336 13001 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 12989 9333 13001 9336
rect 13035 9364 13047 9367
rect 14826 9364 14832 9376
rect 13035 9336 14832 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17770 9364 17776 9376
rect 17368 9336 17776 9364
rect 17368 9324 17374 9336
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 19334 9324 19340 9376
rect 19392 9324 19398 9376
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19518 9364 19524 9376
rect 19475 9336 19524 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 20165 9367 20223 9373
rect 20165 9333 20177 9367
rect 20211 9364 20223 9367
rect 20346 9364 20352 9376
rect 20211 9336 20352 9364
rect 20211 9333 20223 9336
rect 20165 9327 20223 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 21637 9367 21695 9373
rect 21637 9364 21649 9367
rect 21416 9336 21649 9364
rect 21416 9324 21422 9336
rect 21637 9333 21649 9336
rect 21683 9333 21695 9367
rect 22002 9364 22008 9376
rect 21963 9336 22008 9364
rect 21637 9327 21695 9333
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 22462 9364 22468 9376
rect 22423 9336 22468 9364
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 22554 9324 22560 9376
rect 22612 9364 22618 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22612 9336 23029 9364
rect 22612 9324 22618 9336
rect 23017 9333 23029 9336
rect 23063 9364 23075 9367
rect 23308 9364 23336 9392
rect 23063 9336 23336 9364
rect 23063 9333 23075 9336
rect 23017 9327 23075 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2188 9132 2237 9160
rect 2188 9120 2194 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2225 9123 2283 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4982 9160 4988 9172
rect 4203 9132 4988 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 6822 9160 6828 9172
rect 6227 9132 6828 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 9214 9160 9220 9172
rect 9079 9132 9220 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 10686 9160 10692 9172
rect 10643 9132 10692 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 11848 9132 12909 9160
rect 11848 9120 11854 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 13872 9132 15025 9160
rect 13872 9120 13878 9132
rect 15013 9129 15025 9132
rect 15059 9129 15071 9163
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15013 9123 15071 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16850 9160 16856 9172
rect 15804 9132 15849 9160
rect 16811 9132 16856 9160
rect 15804 9120 15810 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17862 9160 17868 9172
rect 17359 9132 17868 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18322 9160 18328 9172
rect 18283 9132 18328 9160
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 20622 9160 20628 9172
rect 20583 9132 20628 9160
rect 19245 9123 19303 9129
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 20898 9120 20904 9172
rect 20956 9160 20962 9172
rect 21085 9163 21143 9169
rect 21085 9160 21097 9163
rect 20956 9132 21097 9160
rect 20956 9120 20962 9132
rect 21085 9129 21097 9132
rect 21131 9129 21143 9163
rect 22922 9160 22928 9172
rect 22883 9132 22928 9160
rect 21085 9123 21143 9129
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 23842 9120 23848 9172
rect 23900 9160 23906 9172
rect 23937 9163 23995 9169
rect 23937 9160 23949 9163
rect 23900 9132 23949 9160
rect 23900 9120 23906 9132
rect 23937 9129 23949 9132
rect 23983 9160 23995 9163
rect 24854 9160 24860 9172
rect 23983 9132 24716 9160
rect 24815 9132 24860 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 1397 9095 1455 9101
rect 1397 9061 1409 9095
rect 1443 9092 1455 9095
rect 2498 9092 2504 9104
rect 1443 9064 2504 9092
rect 1443 9061 1455 9064
rect 1397 9055 1455 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 4617 9095 4675 9101
rect 2599 9064 3915 9092
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2038 9024 2044 9036
rect 1995 8996 2044 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2038 8984 2044 8996
rect 2096 9024 2102 9036
rect 2599 9024 2627 9064
rect 2096 8996 2627 9024
rect 2777 9027 2835 9033
rect 2096 8984 2102 8996
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 3142 9024 3148 9036
rect 2823 8996 3148 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3099 8928 3249 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 2740 8860 3801 8888
rect 2740 8848 2746 8860
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 3887 8888 3915 9064
rect 4617 9061 4629 9095
rect 4663 9092 4675 9095
rect 4706 9092 4712 9104
rect 4663 9064 4712 9092
rect 4663 9061 4675 9064
rect 4617 9055 4675 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 10870 9052 10876 9104
rect 10928 9101 10934 9104
rect 10928 9095 10992 9101
rect 10928 9061 10946 9095
rect 10980 9061 10992 9095
rect 10928 9055 10992 9061
rect 10928 9052 10934 9055
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 16761 9095 16819 9101
rect 13044 9064 13216 9092
rect 13044 9052 13050 9064
rect 4522 9024 4528 9036
rect 4483 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6822 9024 6828 9036
rect 6135 8996 6828 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7374 9024 7380 9036
rect 7331 8996 7380 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7552 9027 7610 9033
rect 7552 8993 7564 9027
rect 7598 9024 7610 9027
rect 7834 9024 7840 9036
rect 7598 8996 7840 9024
rect 7598 8993 7610 8996
rect 7552 8987 7610 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10008 8996 10701 9024
rect 10008 8984 10014 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4028 8928 4813 8956
rect 4028 8916 4034 8928
rect 4801 8925 4813 8928
rect 4847 8956 4859 8959
rect 5534 8956 5540 8968
rect 4847 8928 5540 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 6362 8956 6368 8968
rect 6323 8928 6368 8956
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 12986 8956 12992 8968
rect 12483 8928 12992 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13188 8956 13216 9064
rect 16761 9061 16773 9095
rect 16807 9092 16819 9095
rect 17221 9095 17279 9101
rect 17221 9092 17233 9095
rect 16807 9064 17233 9092
rect 16807 9061 16819 9064
rect 16761 9055 16819 9061
rect 17221 9061 17233 9064
rect 17267 9092 17279 9095
rect 17678 9092 17684 9104
rect 17267 9064 17684 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 20162 9052 20168 9104
rect 20220 9092 20226 9104
rect 20349 9095 20407 9101
rect 20349 9092 20361 9095
rect 20220 9064 20361 9092
rect 20220 9052 20226 9064
rect 20349 9061 20361 9064
rect 20395 9092 20407 9095
rect 20916 9092 20944 9120
rect 21726 9092 21732 9104
rect 20395 9064 20944 9092
rect 21639 9064 21732 9092
rect 20395 9061 20407 9064
rect 20349 9055 20407 9061
rect 21726 9052 21732 9064
rect 21784 9092 21790 9104
rect 24688 9092 24716 9132
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 25225 9163 25283 9169
rect 25225 9160 25237 9163
rect 25188 9132 25237 9160
rect 25188 9120 25194 9132
rect 25225 9129 25237 9132
rect 25271 9129 25283 9163
rect 25590 9160 25596 9172
rect 25551 9132 25596 9160
rect 25225 9123 25283 9129
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 25682 9092 25688 9104
rect 21784 9064 24155 9092
rect 24688 9064 25688 9092
rect 21784 9052 21790 9064
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13320 8996 13369 9024
rect 13320 8984 13326 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 13613 9027 13671 9033
rect 13613 9024 13625 9027
rect 13504 8996 13625 9024
rect 13504 8984 13510 8996
rect 13613 8993 13625 8996
rect 13659 8993 13671 9027
rect 13613 8987 13671 8993
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19484 8996 19625 9024
rect 19484 8984 19490 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 19978 9024 19984 9036
rect 19751 8996 19984 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 13188 8928 13308 8956
rect 13081 8919 13139 8925
rect 5721 8891 5779 8897
rect 3887 8860 4844 8888
rect 3789 8851 3847 8857
rect 4816 8832 4844 8860
rect 5721 8857 5733 8891
rect 5767 8888 5779 8891
rect 7098 8888 7104 8900
rect 5767 8860 7104 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 13096 8888 13124 8919
rect 13280 8900 13308 8928
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15896 8928 15941 8956
rect 15896 8916 15902 8928
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17368 8928 17417 8956
rect 17368 8916 17374 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 19720 8956 19748 8987
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 23845 9027 23903 9033
rect 23845 9024 23857 9027
rect 23532 8996 23857 9024
rect 23532 8984 23538 8996
rect 23845 8993 23857 8996
rect 23891 8993 23903 9027
rect 23845 8987 23903 8993
rect 19886 8956 19892 8968
rect 18831 8928 19748 8956
rect 19847 8928 19892 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21818 8956 21824 8968
rect 21508 8928 21824 8956
rect 21508 8916 21514 8928
rect 21818 8916 21824 8928
rect 21876 8916 21882 8968
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 12084 8860 13124 8888
rect 12084 8832 12112 8860
rect 13262 8848 13268 8900
rect 13320 8848 13326 8900
rect 14366 8848 14372 8900
rect 14424 8888 14430 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 14424 8860 14749 8888
rect 14424 8848 14430 8860
rect 14737 8857 14749 8860
rect 14783 8888 14795 8891
rect 15856 8888 15884 8916
rect 21928 8888 21956 8919
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 24029 8959 24087 8965
rect 24029 8956 24041 8959
rect 22888 8928 24041 8956
rect 22888 8916 22894 8928
rect 24029 8925 24041 8928
rect 24075 8925 24087 8959
rect 24127 8956 24155 9064
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 25038 9024 25044 9036
rect 24999 8996 25044 9024
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 25866 8956 25872 8968
rect 24127 8928 25872 8956
rect 24029 8919 24087 8925
rect 25866 8916 25872 8928
rect 25924 8916 25930 8968
rect 14783 8860 15884 8888
rect 19536 8860 21956 8888
rect 23293 8891 23351 8897
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 19536 8832 19564 8860
rect 23293 8857 23305 8891
rect 23339 8888 23351 8891
rect 24210 8888 24216 8900
rect 23339 8860 24216 8888
rect 23339 8857 23351 8860
rect 23293 8851 23351 8857
rect 24210 8848 24216 8860
rect 24268 8848 24274 8900
rect 24302 8848 24308 8900
rect 24360 8888 24366 8900
rect 24854 8888 24860 8900
rect 24360 8860 24860 8888
rect 24360 8848 24366 8860
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 3513 8823 3571 8829
rect 3513 8820 3525 8823
rect 3283 8792 3525 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3513 8789 3525 8792
rect 3559 8820 3571 8823
rect 3878 8820 3884 8832
rect 3559 8792 3884 8820
rect 3559 8789 3571 8792
rect 3513 8783 3571 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5500 8792 5549 8820
rect 5500 8780 5506 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 8662 8820 8668 8832
rect 8623 8792 8668 8820
rect 5537 8783 5595 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 10226 8820 10232 8832
rect 10187 8792 10232 8820
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 12066 8820 12072 8832
rect 12027 8792 12072 8820
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12216 8792 12541 8820
rect 12216 8780 12222 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 12529 8783 12587 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16390 8820 16396 8832
rect 16351 8792 16396 8820
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 19058 8820 19064 8832
rect 19019 8792 19064 8820
rect 19058 8780 19064 8792
rect 19116 8820 19122 8832
rect 19518 8820 19524 8832
rect 19116 8792 19524 8820
rect 19116 8780 19122 8792
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21361 8823 21419 8829
rect 21361 8820 21373 8823
rect 20772 8792 21373 8820
rect 20772 8780 20778 8792
rect 21361 8789 21373 8792
rect 21407 8789 21419 8823
rect 21361 8783 21419 8789
rect 22465 8823 22523 8829
rect 22465 8789 22477 8823
rect 22511 8820 22523 8823
rect 22830 8820 22836 8832
rect 22511 8792 22836 8820
rect 22511 8789 22523 8792
rect 22465 8783 22523 8789
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 23382 8780 23388 8832
rect 23440 8820 23446 8832
rect 23477 8823 23535 8829
rect 23477 8820 23489 8823
rect 23440 8792 23489 8820
rect 23440 8780 23446 8792
rect 23477 8789 23489 8792
rect 23523 8789 23535 8823
rect 23477 8783 23535 8789
rect 23842 8780 23848 8832
rect 23900 8820 23906 8832
rect 24026 8820 24032 8832
rect 23900 8792 24032 8820
rect 23900 8780 23906 8792
rect 24026 8780 24032 8792
rect 24084 8820 24090 8832
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 24084 8792 24501 8820
rect 24084 8780 24090 8792
rect 24489 8789 24501 8792
rect 24535 8789 24547 8823
rect 24489 8783 24547 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2866 8616 2872 8628
rect 1811 8588 2872 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3016 8588 3249 8616
rect 3016 8576 3022 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 4709 8619 4767 8625
rect 4709 8616 4721 8619
rect 4672 8588 4721 8616
rect 4672 8576 4678 8588
rect 4709 8585 4721 8588
rect 4755 8585 4767 8619
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4709 8579 4767 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8754 8616 8760 8628
rect 8715 8588 8760 8616
rect 8754 8576 8760 8588
rect 8812 8616 8818 8628
rect 10321 8619 10379 8625
rect 8812 8588 9444 8616
rect 8812 8576 8818 8588
rect 2884 8548 2912 8576
rect 4062 8548 4068 8560
rect 2884 8520 4068 8548
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 5905 8551 5963 8557
rect 5905 8548 5917 8551
rect 4580 8520 5917 8548
rect 4580 8508 4586 8520
rect 5905 8517 5917 8520
rect 5951 8517 5963 8551
rect 5905 8511 5963 8517
rect 6641 8551 6699 8557
rect 6641 8517 6653 8551
rect 6687 8548 6699 8551
rect 6687 8520 7696 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 7668 8492 7696 8520
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 5408 8452 5457 8480
rect 5408 8440 5414 8452
rect 5445 8449 5457 8452
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 7156 8452 7481 8480
rect 7156 8440 7162 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7650 8480 7656 8492
rect 7611 8452 7656 8480
rect 7469 8443 7527 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 9416 8489 9444 8588
rect 10321 8585 10333 8619
rect 10367 8616 10379 8619
rect 10870 8616 10876 8628
rect 10367 8588 10876 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11882 8616 11888 8628
rect 11843 8588 11888 8616
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12124 8588 12173 8616
rect 12124 8576 12130 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12161 8579 12219 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 15838 8616 15844 8628
rect 15427 8588 15844 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17862 8616 17868 8628
rect 17727 8588 17868 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18693 8619 18751 8625
rect 18693 8585 18705 8619
rect 18739 8616 18751 8619
rect 19886 8616 19892 8628
rect 18739 8588 19892 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20162 8616 20168 8628
rect 20123 8588 20168 8616
rect 20162 8576 20168 8588
rect 20220 8576 20226 8628
rect 20901 8619 20959 8625
rect 20901 8585 20913 8619
rect 20947 8616 20959 8619
rect 21726 8616 21732 8628
rect 20947 8588 21732 8616
rect 20947 8585 20959 8588
rect 20901 8579 20959 8585
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 22152 8588 22385 8616
rect 22152 8576 22158 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22373 8579 22431 8585
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 23992 8588 25053 8616
rect 23992 8576 23998 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 25682 8616 25688 8628
rect 25643 8588 25688 8616
rect 25041 8579 25099 8585
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 9824 8520 10793 8548
rect 9824 8508 9830 8520
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 11900 8548 11928 8576
rect 11900 8520 12480 8548
rect 10781 8511 10839 8517
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 10735 8452 11345 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 11333 8449 11345 8452
rect 11379 8480 11391 8483
rect 11974 8480 11980 8492
rect 11379 8452 11980 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2130 8421 2136 8424
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1728 8384 1869 8412
rect 1728 8372 1734 8384
rect 1857 8381 1869 8384
rect 1903 8381 1915 8415
rect 2124 8412 2136 8421
rect 2091 8384 2136 8412
rect 1857 8375 1915 8381
rect 2124 8375 2136 8384
rect 2130 8372 2136 8375
rect 2188 8372 2194 8424
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4706 8412 4712 8424
rect 4295 8384 4712 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 9272 8384 9321 8412
rect 9272 8372 9278 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 3200 8316 3525 8344
rect 3200 8304 3206 8316
rect 3513 8313 3525 8316
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 4614 8304 4620 8356
rect 4672 8344 4678 8356
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 4672 8316 5365 8344
rect 4672 8304 4678 8316
rect 5353 8313 5365 8316
rect 5399 8313 5411 8347
rect 5353 8307 5411 8313
rect 8481 8347 8539 8353
rect 8481 8313 8493 8347
rect 8527 8344 8539 8347
rect 8846 8344 8852 8356
rect 8527 8316 8852 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 8846 8304 8852 8316
rect 8904 8344 8910 8356
rect 9508 8344 9536 8443
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 10778 8412 10784 8424
rect 10284 8384 10784 8412
rect 10284 8372 10290 8384
rect 10778 8372 10784 8384
rect 10836 8412 10842 8424
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10836 8384 11161 8412
rect 10836 8372 10842 8384
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 12158 8412 12164 8424
rect 11287 8384 12164 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 8904 8316 9536 8344
rect 8904 8304 8910 8316
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11256 8344 11284 8375
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12452 8421 12480 8520
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 16574 8480 16580 8492
rect 16448 8452 16580 8480
rect 16448 8440 16454 8452
rect 16574 8440 16580 8452
rect 16632 8480 16638 8492
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 16632 8452 16773 8480
rect 16632 8440 16638 8452
rect 16761 8449 16773 8452
rect 16807 8449 16819 8483
rect 23290 8480 23296 8492
rect 23203 8452 23296 8480
rect 16761 8443 16819 8449
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 13808 8415 13866 8421
rect 13587 8384 13768 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 13740 8356 13768 8384
rect 13808 8381 13820 8415
rect 13854 8412 13866 8415
rect 14366 8412 14372 8424
rect 13854 8384 14372 8412
rect 13854 8381 13866 8384
rect 13808 8375 13866 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16666 8412 16672 8424
rect 15795 8384 16672 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 18831 8384 19288 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 11020 8316 11284 8344
rect 11020 8304 11026 8316
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 13078 8344 13084 8356
rect 12860 8316 13084 8344
rect 12860 8304 12866 8316
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 13722 8304 13728 8356
rect 13780 8304 13786 8356
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 13964 8316 16129 8344
rect 13964 8304 13970 8316
rect 16117 8313 16129 8316
rect 16163 8344 16175 8347
rect 18230 8344 18236 8356
rect 16163 8316 16620 8344
rect 18191 8316 18236 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 5258 8276 5264 8288
rect 5219 8248 5264 8276
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 7374 8276 7380 8288
rect 7335 8248 7380 8276
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8021 8279 8079 8285
rect 8021 8276 8033 8279
rect 7892 8248 8033 8276
rect 7892 8236 7898 8248
rect 8021 8245 8033 8248
rect 8067 8245 8079 8279
rect 8021 8239 8079 8245
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9214 8276 9220 8288
rect 8987 8248 9220 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 13630 8276 13636 8288
rect 12492 8248 13636 8276
rect 12492 8236 12498 8248
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 13872 8248 14933 8276
rect 13872 8236 13878 8248
rect 14921 8245 14933 8248
rect 14967 8245 14979 8279
rect 16206 8276 16212 8288
rect 16167 8248 16212 8276
rect 14921 8239 14979 8245
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 16592 8285 16620 8316
rect 18230 8304 18236 8316
rect 18288 8344 18294 8356
rect 19058 8353 19064 8356
rect 19030 8347 19064 8353
rect 19030 8344 19042 8347
rect 18288 8316 19042 8344
rect 18288 8304 18294 8316
rect 19030 8313 19042 8316
rect 19116 8344 19122 8356
rect 19116 8316 19178 8344
rect 19030 8307 19064 8313
rect 19058 8304 19064 8307
rect 19116 8304 19122 8316
rect 16577 8279 16635 8285
rect 16577 8245 16589 8279
rect 16623 8276 16635 8279
rect 17862 8276 17868 8288
rect 16623 8248 17868 8276
rect 16623 8245 16635 8248
rect 16577 8239 16635 8245
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 19260 8276 19288 8384
rect 19518 8372 19524 8424
rect 19576 8412 19582 8424
rect 20441 8415 20499 8421
rect 20441 8412 20453 8415
rect 19576 8384 20453 8412
rect 19576 8372 19582 8384
rect 20441 8381 20453 8384
rect 20487 8381 20499 8415
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20441 8375 20499 8381
rect 20824 8384 21005 8412
rect 20824 8344 20852 8384
rect 20993 8381 21005 8384
rect 21039 8412 21051 8415
rect 21082 8412 21088 8424
rect 21039 8384 21088 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21082 8372 21088 8384
rect 21140 8412 21146 8424
rect 23216 8412 23244 8452
rect 23290 8440 23296 8452
rect 23348 8480 23354 8492
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23348 8452 23673 8480
rect 23348 8440 23354 8452
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 25038 8440 25044 8492
rect 25096 8480 25102 8492
rect 25317 8483 25375 8489
rect 25317 8480 25329 8483
rect 25096 8452 25329 8480
rect 25096 8440 25102 8452
rect 25317 8449 25329 8452
rect 25363 8449 25375 8483
rect 25317 8443 25375 8449
rect 23474 8412 23480 8424
rect 21140 8384 23244 8412
rect 23435 8384 23480 8412
rect 21140 8372 21146 8384
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 20640 8316 20852 8344
rect 20346 8276 20352 8288
rect 19208 8248 20352 8276
rect 19208 8236 19214 8248
rect 20346 8236 20352 8248
rect 20404 8276 20410 8288
rect 20640 8276 20668 8316
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 21238 8347 21296 8353
rect 21238 8344 21250 8347
rect 20956 8316 21250 8344
rect 20956 8304 20962 8316
rect 21238 8313 21250 8316
rect 21284 8313 21296 8347
rect 21238 8307 21296 8313
rect 22462 8304 22468 8356
rect 22520 8344 22526 8356
rect 22741 8347 22799 8353
rect 22741 8344 22753 8347
rect 22520 8316 22753 8344
rect 22520 8304 22526 8316
rect 22741 8313 22753 8316
rect 22787 8344 22799 8347
rect 23928 8347 23986 8353
rect 22787 8316 23520 8344
rect 22787 8313 22799 8316
rect 22741 8307 22799 8313
rect 20404 8248 20668 8276
rect 20404 8236 20410 8248
rect 22830 8236 22836 8288
rect 22888 8276 22894 8288
rect 23109 8279 23167 8285
rect 23109 8276 23121 8279
rect 22888 8248 23121 8276
rect 22888 8236 22894 8248
rect 23109 8245 23121 8248
rect 23155 8276 23167 8279
rect 23290 8276 23296 8288
rect 23155 8248 23296 8276
rect 23155 8245 23167 8248
rect 23109 8239 23167 8245
rect 23290 8236 23296 8248
rect 23348 8236 23354 8288
rect 23492 8276 23520 8316
rect 23928 8313 23940 8347
rect 23974 8344 23986 8347
rect 24210 8344 24216 8356
rect 23974 8316 24216 8344
rect 23974 8313 23986 8316
rect 23928 8307 23986 8313
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 24026 8276 24032 8288
rect 23492 8248 24032 8276
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 25682 8236 25688 8288
rect 25740 8276 25746 8288
rect 26053 8279 26111 8285
rect 26053 8276 26065 8279
rect 25740 8248 26065 8276
rect 25740 8236 25746 8248
rect 26053 8245 26065 8248
rect 26099 8245 26111 8279
rect 26053 8239 26111 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2130 8072 2136 8084
rect 1995 8044 2136 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2130 8032 2136 8044
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 3970 8072 3976 8084
rect 3927 8044 3976 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4246 8072 4252 8084
rect 4203 8044 4252 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4890 8072 4896 8084
rect 4571 8044 4896 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5408 8044 5549 8072
rect 5408 8032 5414 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7374 8072 7380 8084
rect 7055 8044 7380 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7374 8032 7380 8044
rect 7432 8072 7438 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 7432 8044 8401 8072
rect 7432 8032 7438 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 8389 8035 8447 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10962 8072 10968 8084
rect 10551 8044 10968 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12345 8075 12403 8081
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12526 8072 12532 8084
rect 12391 8044 12532 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12526 8032 12532 8044
rect 12584 8072 12590 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12584 8044 12817 8072
rect 12584 8032 12590 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 13044 8044 13185 8072
rect 13044 8032 13050 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 14277 8075 14335 8081
rect 13320 8044 13768 8072
rect 13320 8032 13326 8044
rect 2038 7964 2044 8016
rect 2096 8004 2102 8016
rect 3326 8004 3332 8016
rect 2096 7976 3332 8004
rect 2096 7964 2102 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 5166 7964 5172 8016
rect 5224 8004 5230 8016
rect 5261 8007 5319 8013
rect 5261 8004 5273 8007
rect 5224 7976 5273 8004
rect 5224 7964 5230 7976
rect 5261 7973 5273 7976
rect 5307 8004 5319 8007
rect 5626 8004 5632 8016
rect 5307 7976 5632 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 7469 8007 7527 8013
rect 7469 7973 7481 8007
rect 7515 8004 7527 8007
rect 7926 8004 7932 8016
rect 7515 7976 7932 8004
rect 7515 7973 7527 7976
rect 7469 7967 7527 7973
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 13630 8004 13636 8016
rect 9640 7976 13636 8004
rect 9640 7964 9646 7976
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 3510 7936 3516 7948
rect 2823 7908 3004 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2222 7868 2228 7880
rect 1443 7840 2228 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 2406 7800 2412 7812
rect 2367 7772 2412 7800
rect 2406 7760 2412 7772
rect 2464 7760 2470 7812
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 2976 7800 3004 7908
rect 3068 7908 3516 7936
rect 3068 7877 3096 7908
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 6178 7936 6184 7948
rect 5951 7908 6184 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6972 7908 7389 7936
rect 6972 7896 6978 7908
rect 7377 7905 7389 7908
rect 7423 7936 7435 7939
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7423 7908 8033 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 8021 7905 8033 7908
rect 8067 7905 8079 7939
rect 8021 7899 8079 7905
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10318 7936 10324 7948
rect 9907 7908 10324 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 11232 7939 11290 7945
rect 11232 7905 11244 7939
rect 11278 7936 11290 7939
rect 11790 7936 11796 7948
rect 11278 7908 11796 7936
rect 11278 7905 11290 7908
rect 11232 7899 11290 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4028 7840 4629 7868
rect 4028 7828 4034 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4798 7868 4804 7880
rect 4759 7840 4804 7868
rect 4617 7831 4675 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 6595 7840 7665 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 8570 7868 8576 7880
rect 8531 7840 8576 7868
rect 7653 7831 7711 7837
rect 7668 7800 7696 7831
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10008 7840 10977 7868
rect 10008 7828 10014 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 13004 7868 13032 7976
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13446 7936 13452 7948
rect 13127 7908 13452 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13740 7936 13768 8044
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14366 8072 14372 8084
rect 14323 8044 14372 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15712 8044 16129 8072
rect 15712 8032 15718 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16816 8044 17693 8072
rect 16816 8032 16822 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 18932 8044 19349 8072
rect 18932 8032 18938 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 19337 8035 19395 8041
rect 20073 8075 20131 8081
rect 20073 8041 20085 8075
rect 20119 8072 20131 8075
rect 20162 8072 20168 8084
rect 20119 8044 20168 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20404 8044 20545 8072
rect 20404 8032 20410 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 22278 8072 22284 8084
rect 22239 8044 22284 8072
rect 20533 8035 20591 8041
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 22738 8032 22744 8084
rect 22796 8072 22802 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 22796 8044 23397 8072
rect 22796 8032 22802 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 24670 8072 24676 8084
rect 24631 8044 24676 8072
rect 23385 8035 23443 8041
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 25593 8075 25651 8081
rect 25593 8041 25605 8075
rect 25639 8072 25651 8075
rect 25682 8072 25688 8084
rect 25639 8044 25688 8072
rect 25639 8041 25651 8044
rect 25593 8035 25651 8041
rect 25682 8032 25688 8044
rect 25740 8032 25746 8084
rect 15746 8004 15752 8016
rect 15707 7976 15752 8004
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 16574 8013 16580 8016
rect 16568 8004 16580 8013
rect 16535 7976 16580 8004
rect 16568 7967 16580 7976
rect 16574 7964 16580 7967
rect 16632 7964 16638 8016
rect 18601 8007 18659 8013
rect 18601 7973 18613 8007
rect 18647 8004 18659 8007
rect 19426 8004 19432 8016
rect 18647 7976 19432 8004
rect 18647 7973 18659 7976
rect 18601 7967 18659 7973
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 22189 8007 22247 8013
rect 22189 7973 22201 8007
rect 22235 8004 22247 8007
rect 22925 8007 22983 8013
rect 22925 8004 22937 8007
rect 22235 7976 22937 8004
rect 22235 7973 22247 7976
rect 22189 7967 22247 7973
rect 22925 7973 22937 7976
rect 22971 8004 22983 8007
rect 23106 8004 23112 8016
rect 22971 7976 23112 8004
rect 22971 7973 22983 7976
rect 22925 7967 22983 7973
rect 23106 7964 23112 7976
rect 23164 7964 23170 8016
rect 13587 7908 13768 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13262 7868 13268 7880
rect 13004 7840 13268 7868
rect 10965 7831 11023 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13556 7868 13584 7899
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 16850 7936 16856 7948
rect 14884 7908 16856 7936
rect 14884 7896 14890 7908
rect 16850 7896 16856 7908
rect 16908 7936 16914 7948
rect 17770 7936 17776 7948
rect 16908 7908 17776 7936
rect 16908 7896 16914 7908
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 18380 7908 18889 7936
rect 18380 7896 18386 7908
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 20717 7939 20775 7945
rect 19116 7908 19564 7936
rect 19116 7896 19122 7908
rect 13464 7840 13584 7868
rect 13725 7871 13783 7877
rect 13464 7812 13492 7840
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15838 7868 15844 7880
rect 15335 7840 15844 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 8662 7800 8668 7812
rect 2556 7772 6592 7800
rect 7668 7772 8668 7800
rect 2556 7760 2562 7772
rect 6564 7744 6592 7772
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 10192 7772 10916 7800
rect 10192 7760 10198 7772
rect 10888 7744 10916 7772
rect 13446 7760 13452 7812
rect 13504 7760 13510 7812
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 3050 7732 3056 7744
rect 1636 7704 3056 7732
rect 1636 7692 1642 7704
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7732 7070 7744
rect 7190 7732 7196 7744
rect 7064 7704 7196 7732
rect 7064 7692 7070 7704
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 10042 7732 10048 7744
rect 10003 7704 10048 7732
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 12492 7704 12633 7732
rect 12492 7692 12498 7704
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12621 7695 12679 7701
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 13740 7732 13768 7831
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 16080 7840 16313 7868
rect 16080 7828 16086 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 16301 7831 16359 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 19536 7877 19564 7908
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 20898 7936 20904 7948
rect 20763 7908 20904 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 23198 7896 23204 7948
rect 23256 7936 23262 7948
rect 23753 7939 23811 7945
rect 23753 7936 23765 7939
rect 23256 7908 23765 7936
rect 23256 7896 23262 7908
rect 23753 7905 23765 7908
rect 23799 7905 23811 7939
rect 23753 7899 23811 7905
rect 24949 7939 25007 7945
rect 24949 7905 24961 7939
rect 24995 7936 25007 7939
rect 25498 7936 25504 7948
rect 24995 7908 25504 7936
rect 24995 7905 25007 7908
rect 24949 7899 25007 7905
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 22465 7871 22523 7877
rect 22465 7868 22477 7871
rect 21968 7840 22477 7868
rect 21968 7828 21974 7840
rect 22465 7837 22477 7840
rect 22511 7837 22523 7871
rect 22465 7831 22523 7837
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 23658 7868 23664 7880
rect 23339 7840 23664 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 18969 7803 19027 7809
rect 18969 7769 18981 7803
rect 19015 7800 19027 7803
rect 19242 7800 19248 7812
rect 19015 7772 19248 7800
rect 19015 7769 19027 7772
rect 18969 7763 19027 7769
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 20346 7800 20352 7812
rect 20307 7772 20352 7800
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 22480 7800 22508 7831
rect 23658 7828 23664 7840
rect 23716 7868 23722 7880
rect 23845 7871 23903 7877
rect 23845 7868 23857 7871
rect 23716 7840 23857 7868
rect 23716 7828 23722 7840
rect 23845 7837 23857 7840
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 23992 7840 24037 7868
rect 23992 7828 23998 7840
rect 22480 7772 23336 7800
rect 23308 7744 23336 7772
rect 12851 7704 13768 7732
rect 14645 7735 14703 7741
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 14826 7732 14832 7744
rect 14691 7704 14832 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 14826 7692 14832 7704
rect 14884 7732 14890 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14884 7704 14933 7732
rect 14884 7692 14890 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 14921 7695 14979 7701
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18230 7732 18236 7744
rect 18187 7704 18236 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 18690 7732 18696 7744
rect 18651 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 21450 7732 21456 7744
rect 21411 7704 21456 7732
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21818 7732 21824 7744
rect 21779 7704 21824 7732
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 23290 7692 23296 7744
rect 23348 7692 23354 7744
rect 25130 7732 25136 7744
rect 25091 7704 25136 7732
rect 25130 7692 25136 7704
rect 25188 7692 25194 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2866 7528 2872 7540
rect 2363 7500 2872 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3050 7488 3056 7540
rect 3108 7488 3114 7540
rect 3970 7528 3976 7540
rect 3931 7500 3976 7528
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 4982 7528 4988 7540
rect 4755 7500 4988 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 6914 7528 6920 7540
rect 6875 7500 6920 7528
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 8021 7531 8079 7537
rect 8021 7497 8033 7531
rect 8067 7528 8079 7531
rect 8570 7528 8576 7540
rect 8067 7500 8576 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 1949 7463 2007 7469
rect 1949 7429 1961 7463
rect 1995 7460 2007 7463
rect 2498 7460 2504 7472
rect 1995 7432 2504 7460
rect 1995 7429 2007 7432
rect 1949 7423 2007 7429
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 3068 7460 3096 7488
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 3068 7432 6561 7460
rect 6549 7429 6561 7432
rect 6595 7460 6607 7463
rect 6595 7432 7420 7460
rect 6595 7429 6607 7432
rect 6549 7423 6607 7429
rect 3050 7392 3056 7404
rect 3011 7364 3056 7392
rect 3050 7352 3056 7364
rect 3108 7392 3114 7404
rect 3421 7395 3479 7401
rect 3421 7392 3433 7395
rect 3108 7364 3433 7392
rect 3108 7352 3114 7364
rect 3421 7361 3433 7364
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 5258 7392 5264 7404
rect 4203 7364 5264 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5629 7355 5687 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 7392 7401 7420 7432
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7834 7392 7840 7404
rect 7607 7364 7840 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 2866 7324 2872 7336
rect 2823 7296 2872 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 8036 7324 8064 7491
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 10318 7528 10324 7540
rect 8720 7500 8765 7528
rect 10279 7500 10324 7528
rect 8720 7488 8726 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10781 7531 10839 7537
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 11054 7528 11060 7540
rect 10827 7500 11060 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12526 7528 12532 7540
rect 12299 7500 12532 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 12158 7460 12164 7472
rect 10192 7432 12164 7460
rect 10192 7420 10198 7432
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9766 7392 9772 7404
rect 9171 7364 9772 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7392 11483 7395
rect 11698 7392 11704 7404
rect 11471 7364 11704 7392
rect 11471 7361 11483 7364
rect 11425 7355 11483 7361
rect 11698 7352 11704 7364
rect 11756 7392 11762 7404
rect 12268 7392 12296 7491
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 16206 7528 16212 7540
rect 15703 7500 16212 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 18932 7500 19073 7528
rect 18932 7488 18938 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19061 7491 19119 7497
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 19889 7531 19947 7537
rect 19889 7497 19901 7531
rect 19935 7528 19947 7531
rect 19978 7528 19984 7540
rect 19935 7500 19984 7528
rect 19935 7497 19947 7500
rect 19889 7491 19947 7497
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 21910 7528 21916 7540
rect 21871 7500 21916 7528
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 22833 7531 22891 7537
rect 22833 7497 22845 7531
rect 22879 7528 22891 7531
rect 23109 7531 23167 7537
rect 23109 7528 23121 7531
rect 22879 7500 23121 7528
rect 22879 7497 22891 7500
rect 22833 7491 22891 7497
rect 23109 7497 23121 7500
rect 23155 7528 23167 7531
rect 23382 7528 23388 7540
rect 23155 7500 23388 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 23934 7528 23940 7540
rect 23523 7500 23940 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 23934 7488 23940 7500
rect 23992 7488 23998 7540
rect 24026 7488 24032 7540
rect 24084 7528 24090 7540
rect 24581 7531 24639 7537
rect 24581 7528 24593 7531
rect 24084 7500 24593 7528
rect 24084 7488 24090 7500
rect 24581 7497 24593 7500
rect 24627 7497 24639 7531
rect 25958 7528 25964 7540
rect 25919 7500 25964 7528
rect 24581 7491 24639 7497
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 16758 7460 16764 7472
rect 16071 7432 16764 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 16758 7420 16764 7432
rect 16816 7460 16822 7472
rect 21545 7463 21603 7469
rect 16816 7432 16988 7460
rect 16816 7420 16822 7432
rect 11756 7364 12296 7392
rect 11756 7352 11762 7364
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16960 7401 16988 7432
rect 21545 7429 21557 7463
rect 21591 7460 21603 7463
rect 24210 7460 24216 7472
rect 21591 7432 24216 7460
rect 21591 7429 21603 7432
rect 21545 7423 21603 7429
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16264 7364 16865 7392
rect 16264 7352 16270 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 18288 7364 18705 7392
rect 18288 7352 18294 7364
rect 18693 7361 18705 7364
rect 18739 7392 18751 7395
rect 18874 7392 18880 7404
rect 18739 7364 18880 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 22664 7401 22692 7432
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20220 7364 20453 7392
rect 20220 7352 20226 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24728 7364 25053 7392
rect 24728 7352 24734 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 7331 7296 8064 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9272 7296 9597 7324
rect 9272 7284 9278 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 13541 7327 13599 7333
rect 12492 7296 12537 7324
rect 12492 7284 12498 7296
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 13630 7324 13636 7336
rect 13587 7296 13636 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13814 7333 13820 7336
rect 13808 7324 13820 7333
rect 13775 7296 13820 7324
rect 13808 7287 13820 7296
rect 13814 7284 13820 7287
rect 13872 7284 13878 7336
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 16298 7324 16304 7336
rect 15335 7296 16304 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18104 7296 18521 7324
rect 18104 7284 18110 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7324 20407 7327
rect 20622 7324 20628 7336
rect 20395 7296 20628 7324
rect 20395 7293 20407 7296
rect 20349 7287 20407 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7324 22431 7327
rect 22833 7327 22891 7333
rect 22833 7324 22845 7327
rect 22419 7296 22845 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 22833 7293 22845 7296
rect 22879 7293 22891 7327
rect 22833 7287 22891 7293
rect 4338 7216 4344 7268
rect 4396 7256 4402 7268
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 4396 7228 5089 7256
rect 4396 7216 4402 7228
rect 5077 7225 5089 7228
rect 5123 7256 5135 7259
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5123 7228 5549 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 5994 7256 6000 7268
rect 5583 7228 6000 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 10704 7228 11253 7256
rect 10704 7200 10732 7228
rect 11241 7225 11253 7228
rect 11287 7225 11299 7259
rect 13906 7256 13912 7268
rect 11241 7219 11299 7225
rect 11624 7228 13912 7256
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2188 7160 2421 7188
rect 2188 7148 2194 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 3326 7188 3332 7200
rect 2915 7160 3332 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6273 7191 6331 7197
rect 6273 7188 6285 7191
rect 6236 7160 6285 7188
rect 6236 7148 6242 7160
rect 6273 7157 6285 7160
rect 6319 7188 6331 7191
rect 6914 7188 6920 7200
rect 6319 7160 6920 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7892 7160 8309 7188
rect 7892 7148 7898 7160
rect 8297 7157 8309 7160
rect 8343 7157 8355 7191
rect 8297 7151 8355 7157
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9490 7188 9496 7200
rect 9263 7160 9496 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9640 7160 9689 7188
rect 9640 7148 9646 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 9677 7151 9735 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10928 7160 11161 7188
rect 10928 7148 10934 7160
rect 11149 7157 11161 7160
rect 11195 7188 11207 7191
rect 11624 7188 11652 7228
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 16724 7228 16773 7256
rect 16724 7216 16730 7228
rect 16761 7225 16773 7228
rect 16807 7256 16819 7259
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 16807 7228 17417 7256
rect 16807 7225 16819 7228
rect 16761 7219 16819 7225
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 17405 7219 17463 7225
rect 17770 7216 17776 7268
rect 17828 7256 17834 7268
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 17828 7228 18429 7256
rect 17828 7216 17834 7228
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 23290 7216 23296 7268
rect 23348 7256 23354 7268
rect 24029 7259 24087 7265
rect 24029 7256 24041 7259
rect 23348 7228 24041 7256
rect 23348 7216 23354 7228
rect 24029 7225 24041 7228
rect 24075 7256 24087 7259
rect 24854 7256 24860 7268
rect 24075 7228 24860 7256
rect 24075 7225 24087 7228
rect 24029 7219 24087 7225
rect 24854 7216 24860 7228
rect 24912 7256 24918 7268
rect 25148 7256 25176 7355
rect 26142 7256 26148 7268
rect 24912 7228 25176 7256
rect 25240 7228 26148 7256
rect 24912 7216 24918 7228
rect 11790 7188 11796 7200
rect 11195 7160 11652 7188
rect 11751 7160 11796 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 12618 7188 12624 7200
rect 12579 7160 12624 7188
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 12860 7160 13185 7188
rect 12860 7148 12866 7160
rect 13173 7157 13185 7160
rect 13219 7188 13231 7191
rect 13446 7188 13452 7200
rect 13219 7160 13452 7188
rect 13219 7157 13231 7160
rect 13173 7151 13231 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14424 7160 14933 7188
rect 14424 7148 14430 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 14921 7151 14979 7157
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 16022 7188 16028 7200
rect 15620 7160 16028 7188
rect 15620 7148 15626 7160
rect 16022 7148 16028 7160
rect 16080 7188 16086 7200
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 16080 7160 16129 7188
rect 16080 7148 16086 7160
rect 16117 7157 16129 7160
rect 16163 7157 16175 7191
rect 16117 7151 16175 7157
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7188 16451 7191
rect 16482 7188 16488 7200
rect 16439 7160 16488 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18322 7188 18328 7200
rect 18095 7160 18328 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 20257 7191 20315 7197
rect 20257 7157 20269 7191
rect 20303 7188 20315 7191
rect 20346 7188 20352 7200
rect 20303 7160 20352 7188
rect 20303 7157 20315 7160
rect 20257 7151 20315 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 22005 7191 22063 7197
rect 22005 7157 22017 7191
rect 22051 7188 22063 7191
rect 22094 7188 22100 7200
rect 22051 7160 22100 7188
rect 22051 7157 22063 7160
rect 22005 7151 22063 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24949 7191 25007 7197
rect 24949 7188 24961 7191
rect 24535 7160 24961 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24949 7157 24961 7160
rect 24995 7188 25007 7191
rect 25240 7188 25268 7228
rect 26142 7216 26148 7228
rect 26200 7216 26206 7268
rect 24995 7160 25268 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25593 7191 25651 7197
rect 25593 7188 25605 7191
rect 25556 7160 25605 7188
rect 25556 7148 25562 7160
rect 25593 7157 25605 7160
rect 25639 7157 25651 7191
rect 25593 7151 25651 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2961 6987 3019 6993
rect 2961 6953 2973 6987
rect 3007 6984 3019 6987
rect 3418 6984 3424 6996
rect 3007 6956 3424 6984
rect 3007 6953 3019 6956
rect 2961 6947 3019 6953
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 5074 6984 5080 6996
rect 5035 6956 5080 6984
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 5994 6984 6000 6996
rect 5868 6956 6000 6984
rect 5868 6944 5874 6956
rect 5994 6944 6000 6956
rect 6052 6984 6058 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 6052 6956 6101 6984
rect 6052 6944 6058 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 8202 6984 8208 6996
rect 7055 6956 8208 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 1486 6876 1492 6928
rect 1544 6916 1550 6928
rect 2041 6919 2099 6925
rect 2041 6916 2053 6919
rect 1544 6888 2053 6916
rect 1544 6876 1550 6888
rect 2041 6885 2053 6888
rect 2087 6916 2099 6919
rect 2682 6916 2688 6928
rect 2087 6888 2688 6916
rect 2087 6885 2099 6888
rect 2041 6879 2099 6885
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 5445 6919 5503 6925
rect 5445 6885 5457 6919
rect 5491 6916 5503 6919
rect 5534 6916 5540 6928
rect 5491 6888 5540 6916
rect 5491 6885 5503 6888
rect 5445 6879 5503 6885
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 7024 6916 7052 6947
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 11698 6984 11704 6996
rect 11659 6956 11704 6984
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12492 6956 12541 6984
rect 12492 6944 12498 6956
rect 12529 6953 12541 6956
rect 12575 6953 12587 6987
rect 13262 6984 13268 6996
rect 13223 6956 13268 6984
rect 12529 6947 12587 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 16666 6984 16672 6996
rect 14016 6956 16528 6984
rect 16627 6956 16672 6984
rect 6840 6888 7052 6916
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5350 6848 5356 6860
rect 4663 6820 5356 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 6178 6848 6184 6860
rect 5552 6820 6184 6848
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2590 6780 2596 6792
rect 2363 6752 2596 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4212 6752 4905 6780
rect 4212 6740 4218 6752
rect 4893 6749 4905 6752
rect 4939 6780 4951 6783
rect 5258 6780 5264 6792
rect 4939 6752 5264 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1762 6712 1768 6724
rect 1719 6684 1768 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 5368 6712 5396 6808
rect 5552 6789 5580 6820
rect 6178 6808 6184 6820
rect 6236 6848 6242 6860
rect 6454 6848 6460 6860
rect 6236 6820 6460 6848
rect 6236 6808 6242 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6840 6848 6868 6888
rect 9858 6876 9864 6928
rect 9916 6916 9922 6928
rect 14016 6916 14044 6956
rect 9916 6888 14044 6916
rect 9916 6876 9922 6888
rect 14090 6876 14096 6928
rect 14148 6916 14154 6928
rect 14734 6916 14740 6928
rect 14148 6888 14740 6916
rect 14148 6876 14154 6888
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 16500 6916 16528 6956
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 17034 6984 17040 6996
rect 16995 6956 17040 6984
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19576 6956 19625 6984
rect 19576 6944 19582 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 19613 6947 19671 6953
rect 20349 6987 20407 6993
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20622 6984 20628 6996
rect 20395 6956 20628 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22557 6987 22615 6993
rect 22557 6984 22569 6987
rect 22336 6956 22569 6984
rect 22336 6944 22342 6956
rect 22557 6953 22569 6956
rect 22603 6953 22615 6987
rect 22557 6947 22615 6953
rect 17218 6916 17224 6928
rect 16500 6888 17224 6916
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 18230 6916 18236 6928
rect 17880 6888 18236 6916
rect 8386 6848 8392 6860
rect 6696 6820 6868 6848
rect 8347 6820 8392 6848
rect 6696 6808 6702 6820
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8570 6848 8576 6860
rect 8527 6820 8576 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9582 6848 9588 6860
rect 9355 6820 9588 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10226 6857 10232 6860
rect 10209 6851 10232 6857
rect 10209 6848 10221 6851
rect 9824 6820 10221 6848
rect 9824 6808 9830 6820
rect 10209 6817 10221 6820
rect 10284 6848 10290 6860
rect 10284 6820 10357 6848
rect 10209 6811 10232 6817
rect 10226 6808 10232 6811
rect 10284 6808 10290 6820
rect 11422 6808 11428 6860
rect 11480 6848 11486 6860
rect 11698 6848 11704 6860
rect 11480 6820 11704 6848
rect 11480 6808 11486 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 11940 6820 12633 6848
rect 11940 6808 11946 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 13906 6848 13912 6860
rect 13867 6820 13912 6848
rect 12621 6811 12679 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 15286 6848 15292 6860
rect 15247 6820 15292 6848
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6848 16451 6851
rect 16574 6848 16580 6860
rect 16439 6820 16580 6848
rect 16439 6817 16451 6820
rect 16393 6811 16451 6817
rect 16574 6808 16580 6820
rect 16632 6848 16638 6860
rect 17773 6851 17831 6857
rect 16632 6820 17264 6848
rect 16632 6808 16638 6820
rect 17236 6792 17264 6820
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 17880 6848 17908 6888
rect 18230 6876 18236 6888
rect 18288 6876 18294 6928
rect 21100 6888 21680 6916
rect 19058 6848 19064 6860
rect 17819 6820 17908 6848
rect 19019 6820 19064 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19392 6820 19717 6848
rect 19392 6808 19398 6820
rect 19705 6817 19717 6820
rect 19751 6848 19763 6851
rect 20438 6848 20444 6860
rect 19751 6820 20444 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 20990 6848 20996 6860
rect 20947 6820 20996 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 20990 6808 20996 6820
rect 21048 6848 21054 6860
rect 21100 6848 21128 6888
rect 21048 6820 21128 6848
rect 21168 6851 21226 6857
rect 21048 6808 21054 6820
rect 21168 6817 21180 6851
rect 21214 6848 21226 6851
rect 21542 6848 21548 6860
rect 21214 6820 21548 6848
rect 21214 6817 21226 6820
rect 21168 6811 21226 6817
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 21652 6848 21680 6888
rect 21652 6820 21956 6848
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 5629 6743 5687 6749
rect 5644 6712 5672 6743
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 8202 6780 8208 6792
rect 7331 6752 8208 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9950 6780 9956 6792
rect 9911 6752 9956 6780
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12124 6752 12725 6780
rect 12124 6740 12130 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13814 6780 13820 6792
rect 13679 6752 13820 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 15470 6780 15476 6792
rect 15431 6752 15476 6780
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 5368 6684 5672 6712
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11977 6715 12035 6721
rect 11977 6712 11989 6715
rect 11112 6684 11989 6712
rect 11112 6672 11118 6684
rect 11977 6681 11989 6684
rect 12023 6681 12035 6715
rect 12158 6712 12164 6724
rect 12119 6684 12164 6712
rect 11977 6675 12035 6681
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 13832 6712 13860 6740
rect 14182 6712 14188 6724
rect 13832 6684 14188 6712
rect 14182 6672 14188 6684
rect 14240 6672 14246 6724
rect 17144 6712 17172 6743
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 18230 6780 18236 6792
rect 17276 6752 17369 6780
rect 18191 6752 18236 6780
rect 17276 6740 17282 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 20070 6780 20076 6792
rect 19935 6752 20076 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 21928 6780 21956 6820
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 23017 6851 23075 6857
rect 23017 6848 23029 6851
rect 22152 6820 23029 6848
rect 22152 6808 22158 6820
rect 23017 6817 23029 6820
rect 23063 6848 23075 6851
rect 23198 6848 23204 6860
rect 23063 6820 23204 6848
rect 23063 6817 23075 6820
rect 23017 6811 23075 6817
rect 23198 6808 23204 6820
rect 23256 6808 23262 6860
rect 23382 6857 23388 6860
rect 23376 6848 23388 6857
rect 23343 6820 23388 6848
rect 23376 6811 23388 6820
rect 23382 6808 23388 6811
rect 23440 6808 23446 6860
rect 25314 6848 25320 6860
rect 25275 6820 25320 6848
rect 25314 6808 25320 6820
rect 25372 6808 25378 6860
rect 23109 6783 23167 6789
rect 23109 6780 23121 6783
rect 21928 6752 23121 6780
rect 23109 6749 23121 6752
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 17494 6712 17500 6724
rect 17144 6684 17500 6712
rect 17494 6672 17500 6684
rect 17552 6672 17558 6724
rect 19242 6712 19248 6724
rect 19203 6684 19248 6712
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 24118 6672 24124 6724
rect 24176 6712 24182 6724
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 24176 6684 24777 6712
rect 24176 6672 24182 6684
rect 24765 6681 24777 6684
rect 24811 6681 24823 6715
rect 24765 6675 24823 6681
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3418 6644 3424 6656
rect 3375 6616 3424 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6595 6616 6653 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 6641 6613 6653 6616
rect 6687 6644 6699 6647
rect 7098 6644 7104 6656
rect 6687 6616 7104 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7432 6616 7665 6644
rect 7432 6604 7438 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 7984 6616 8033 6644
rect 7984 6604 7990 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 8021 6607 8079 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8662 6644 8668 6656
rect 8623 6616 8668 6644
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 10928 6616 11345 6644
rect 10928 6604 10934 6616
rect 11333 6613 11345 6616
rect 11379 6644 11391 6647
rect 11790 6644 11796 6656
rect 11379 6616 11796 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 14826 6644 14832 6656
rect 14783 6616 14832 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 14826 6604 14832 6616
rect 14884 6644 14890 6656
rect 15105 6647 15163 6653
rect 15105 6644 15117 6647
rect 14884 6616 15117 6644
rect 14884 6604 14890 6616
rect 15105 6613 15117 6616
rect 15151 6644 15163 6647
rect 17310 6644 17316 6656
rect 15151 6616 17316 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 21266 6644 21272 6656
rect 20763 6616 21272 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 22152 6616 22293 6644
rect 22152 6604 22158 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 24210 6604 24216 6656
rect 24268 6644 24274 6656
rect 24489 6647 24547 6653
rect 24489 6644 24501 6647
rect 24268 6616 24501 6644
rect 24268 6604 24274 6616
rect 24489 6613 24501 6616
rect 24535 6644 24547 6647
rect 24670 6644 24676 6656
rect 24535 6616 24676 6644
rect 24535 6613 24547 6616
rect 24489 6607 24547 6613
rect 24670 6604 24676 6616
rect 24728 6604 24734 6656
rect 25130 6644 25136 6656
rect 25091 6616 25136 6644
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 25501 6647 25559 6653
rect 25501 6644 25513 6647
rect 25280 6616 25513 6644
rect 25280 6604 25286 6616
rect 25501 6613 25513 6616
rect 25547 6613 25559 6647
rect 25501 6607 25559 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2314 6440 2320 6452
rect 2087 6412 2320 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6403
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 5169 6443 5227 6449
rect 5169 6409 5181 6443
rect 5215 6440 5227 6443
rect 5442 6440 5448 6452
rect 5215 6412 5448 6440
rect 5215 6409 5227 6412
rect 5169 6403 5227 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8294 6440 8300 6452
rect 7975 6412 8300 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8570 6440 8576 6452
rect 8531 6412 8576 6440
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 8846 6440 8852 6452
rect 8807 6412 8852 6440
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10284 6412 10425 6440
rect 10284 6400 10290 6412
rect 10413 6409 10425 6412
rect 10459 6440 10471 6443
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10459 6412 10701 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 11146 6440 11152 6452
rect 11107 6412 11152 6440
rect 10689 6403 10747 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12342 6440 12348 6452
rect 11931 6412 12348 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 14550 6440 14556 6452
rect 13228 6412 14556 6440
rect 13228 6400 13234 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 17129 6443 17187 6449
rect 17129 6409 17141 6443
rect 17175 6440 17187 6443
rect 17218 6440 17224 6452
rect 17175 6412 17224 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 17218 6400 17224 6412
rect 17276 6440 17282 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17276 6412 17785 6440
rect 17276 6400 17282 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 19334 6440 19340 6452
rect 18555 6412 19340 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 20257 6443 20315 6449
rect 20257 6440 20269 6443
rect 19576 6412 20269 6440
rect 19576 6400 19582 6412
rect 20257 6409 20269 6412
rect 20303 6409 20315 6443
rect 20806 6440 20812 6452
rect 20767 6412 20812 6440
rect 20257 6403 20315 6409
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21542 6400 21548 6452
rect 21600 6440 21606 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21600 6412 21833 6440
rect 21600 6400 21606 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 23658 6440 23664 6452
rect 23619 6412 23664 6440
rect 21821 6403 21879 6409
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 25038 6440 25044 6452
rect 24999 6412 25044 6440
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 25682 6400 25688 6452
rect 25740 6440 25746 6452
rect 26329 6443 26387 6449
rect 26329 6440 26341 6443
rect 25740 6412 26341 6440
rect 25740 6400 25746 6412
rect 26329 6409 26341 6412
rect 26375 6409 26387 6443
rect 26329 6403 26387 6409
rect 4065 6375 4123 6381
rect 4065 6341 4077 6375
rect 4111 6372 4123 6375
rect 5350 6372 5356 6384
rect 4111 6344 5356 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 5350 6332 5356 6344
rect 5408 6372 5414 6384
rect 5408 6344 5764 6372
rect 5408 6332 5414 6344
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 5626 6304 5632 6316
rect 4479 6276 5632 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5736 6313 5764 6344
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 5721 6267 5779 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8864 6304 8892 6400
rect 13725 6375 13783 6381
rect 13725 6341 13737 6375
rect 13771 6372 13783 6375
rect 15286 6372 15292 6384
rect 13771 6344 15292 6372
rect 13771 6341 13783 6344
rect 13725 6335 13783 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 17494 6372 17500 6384
rect 17455 6344 17500 6372
rect 17494 6332 17500 6344
rect 17552 6332 17558 6384
rect 20622 6332 20628 6384
rect 20680 6372 20686 6384
rect 20717 6375 20775 6381
rect 20717 6372 20729 6375
rect 20680 6344 20729 6372
rect 20680 6332 20686 6344
rect 20717 6341 20729 6344
rect 20763 6372 20775 6375
rect 20763 6344 21404 6372
rect 20763 6341 20775 6344
rect 20717 6335 20775 6341
rect 13633 6307 13691 6313
rect 8864 6276 9168 6304
rect 1443 6208 2084 6236
rect 3329 6239 3387 6245
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3510 6236 3516 6248
rect 3375 6208 3516 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 5074 6236 5080 6248
rect 5035 6208 5080 6236
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5316 6208 5549 6236
rect 5316 6196 5322 6208
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 2498 6168 2504 6180
rect 1596 6140 2504 6168
rect 1596 6109 1624 6140
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 4801 6171 4859 6177
rect 2823 6140 3188 6168
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 3160 6112 3188 6140
rect 4801 6137 4813 6171
rect 4847 6168 4859 6171
rect 5442 6168 5448 6180
rect 4847 6140 5448 6168
rect 4847 6137 4859 6140
rect 4801 6131 4859 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5552 6168 5580 6199
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6730 6236 6736 6248
rect 6144 6208 6736 6236
rect 6144 6196 6150 6208
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7156 6208 7297 6236
rect 7156 6196 7162 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 9030 6236 9036 6248
rect 9088 6245 9094 6248
rect 8943 6208 9036 6236
rect 7285 6199 7343 6205
rect 9017 6196 9036 6208
rect 9088 6199 9098 6245
rect 9140 6236 9168 6276
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 14366 6304 14372 6316
rect 13679 6276 14372 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 21266 6304 21272 6316
rect 21227 6276 21272 6304
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21376 6313 21404 6344
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6273 21419 6307
rect 22186 6304 22192 6316
rect 22147 6276 22192 6304
rect 21361 6267 21419 6273
rect 22186 6264 22192 6276
rect 22244 6304 22250 6316
rect 24118 6304 24124 6316
rect 22244 6276 22416 6304
rect 24079 6276 24124 6304
rect 22244 6264 22250 6276
rect 9289 6239 9347 6245
rect 9289 6236 9301 6239
rect 9140 6208 9301 6236
rect 9289 6205 9301 6208
rect 9335 6236 9347 6239
rect 9582 6236 9588 6248
rect 9335 6208 9588 6236
rect 9335 6205 9347 6208
rect 9289 6199 9347 6205
rect 9088 6196 9094 6199
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 11204 6208 11253 6236
rect 11204 6196 11210 6208
rect 11241 6205 11253 6208
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12526 6236 12532 6248
rect 12483 6208 12532 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12526 6196 12532 6208
rect 12584 6236 12590 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12584 6208 13185 6236
rect 12584 6196 12590 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 15620 6208 15761 6236
rect 15620 6196 15626 6208
rect 15749 6205 15761 6208
rect 15795 6236 15807 6239
rect 17954 6236 17960 6248
rect 15795 6208 17960 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 17954 6196 17960 6208
rect 18012 6236 18018 6248
rect 18414 6236 18420 6248
rect 18012 6208 18420 6236
rect 18012 6196 18018 6208
rect 18414 6196 18420 6208
rect 18472 6236 18478 6248
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 18472 6208 18613 6236
rect 18472 6196 18478 6208
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 22388 6245 22416 6276
rect 24118 6264 24124 6276
rect 24176 6264 24182 6316
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6304 24363 6307
rect 24670 6304 24676 6316
rect 24351 6276 24676 6304
rect 24351 6273 24363 6276
rect 24305 6267 24363 6273
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 25406 6304 25412 6316
rect 25367 6276 25412 6304
rect 25406 6264 25412 6276
rect 25464 6264 25470 6316
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 20956 6208 21189 6236
rect 20956 6196 20962 6208
rect 21177 6205 21189 6208
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 22373 6239 22431 6245
rect 22373 6205 22385 6239
rect 22419 6205 22431 6239
rect 24026 6236 24032 6248
rect 23987 6208 24032 6236
rect 22373 6199 22431 6205
rect 24026 6196 24032 6208
rect 24084 6196 24090 6248
rect 25038 6196 25044 6248
rect 25096 6236 25102 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25096 6208 25237 6236
rect 25096 6196 25102 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 9017 6168 9045 6196
rect 10042 6168 10048 6180
rect 5552 6140 6684 6168
rect 9017 6140 10048 6168
rect 6656 6112 6684 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 12713 6171 12771 6177
rect 12713 6137 12725 6171
rect 12759 6137 12771 6171
rect 12713 6131 12771 6137
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 2590 6100 2596 6112
rect 2455 6072 2596 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 2924 6072 2969 6100
rect 2924 6060 2930 6072
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3237 6103 3295 6109
rect 3237 6100 3249 6103
rect 3200 6072 3249 6100
rect 3200 6060 3206 6072
rect 3237 6069 3249 6072
rect 3283 6069 3295 6103
rect 3237 6063 3295 6069
rect 4893 6103 4951 6109
rect 4893 6069 4905 6103
rect 4939 6100 4951 6103
rect 5074 6100 5080 6112
rect 4939 6072 5080 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 6638 6060 6644 6112
rect 6696 6060 6702 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 11422 6100 11428 6112
rect 11383 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12158 6100 12164 6112
rect 11940 6072 12164 6100
rect 11940 6060 11946 6072
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12728 6100 12756 6131
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13688 6140 14105 6168
rect 13688 6128 13694 6140
rect 14093 6137 14105 6140
rect 14139 6168 14151 6171
rect 15105 6171 15163 6177
rect 15105 6168 15117 6171
rect 14139 6140 15117 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 15105 6137 15117 6140
rect 15151 6137 15163 6171
rect 15654 6168 15660 6180
rect 15567 6140 15660 6168
rect 15105 6131 15163 6137
rect 15654 6128 15660 6140
rect 15712 6168 15718 6180
rect 15994 6171 16052 6177
rect 15994 6168 16006 6171
rect 15712 6140 16006 6168
rect 15712 6128 15718 6140
rect 15994 6137 16006 6140
rect 16040 6137 16052 6171
rect 15994 6131 16052 6137
rect 18506 6128 18512 6180
rect 18564 6168 18570 6180
rect 18846 6171 18904 6177
rect 18846 6168 18858 6171
rect 18564 6140 18858 6168
rect 18564 6128 18570 6140
rect 18846 6137 18858 6140
rect 18892 6137 18904 6171
rect 18846 6131 18904 6137
rect 19426 6128 19432 6180
rect 19484 6168 19490 6180
rect 26510 6168 26516 6180
rect 19484 6140 26516 6168
rect 19484 6128 19490 6140
rect 26510 6128 26516 6140
rect 26568 6128 26574 6180
rect 13722 6100 13728 6112
rect 12728 6072 13728 6100
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13872 6072 14197 6100
rect 13872 6060 13878 6072
rect 14185 6069 14197 6072
rect 14231 6100 14243 6103
rect 14737 6103 14795 6109
rect 14737 6100 14749 6103
rect 14231 6072 14749 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14737 6069 14749 6072
rect 14783 6069 14795 6103
rect 14737 6063 14795 6069
rect 19981 6103 20039 6109
rect 19981 6069 19993 6103
rect 20027 6100 20039 6103
rect 20070 6100 20076 6112
rect 20027 6072 20076 6100
rect 20027 6069 20039 6072
rect 19981 6063 20039 6069
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 22554 6100 22560 6112
rect 22515 6072 22560 6100
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 23201 6103 23259 6109
rect 23201 6069 23213 6103
rect 23247 6100 23259 6103
rect 23382 6100 23388 6112
rect 23247 6072 23388 6100
rect 23247 6069 23259 6072
rect 23201 6063 23259 6069
rect 23382 6060 23388 6072
rect 23440 6100 23446 6112
rect 24670 6100 24676 6112
rect 23440 6072 24676 6100
rect 23440 6060 23446 6072
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 25958 6100 25964 6112
rect 25919 6072 25964 6100
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 2924 5868 3709 5896
rect 2924 5856 2930 5868
rect 3697 5865 3709 5868
rect 3743 5865 3755 5899
rect 3697 5859 3755 5865
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4798 5896 4804 5908
rect 3936 5868 4804 5896
rect 3936 5856 3942 5868
rect 4798 5856 4804 5868
rect 4856 5896 4862 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 4856 5868 5457 5896
rect 4856 5856 4862 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 7190 5896 7196 5908
rect 6411 5868 7196 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7432 5868 7849 5896
rect 7432 5856 7438 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 8260 5868 8585 5896
rect 8260 5856 8266 5868
rect 8573 5865 8585 5868
rect 8619 5896 8631 5899
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8619 5868 8953 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 3326 5828 3332 5840
rect 3287 5800 3332 5828
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 5074 5828 5080 5840
rect 4080 5800 5080 5828
rect 1670 5760 1676 5772
rect 1631 5732 1676 5760
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 1946 5769 1952 5772
rect 1940 5760 1952 5769
rect 1907 5732 1952 5760
rect 1940 5723 1952 5732
rect 2004 5760 2010 5772
rect 3418 5760 3424 5772
rect 2004 5732 3424 5760
rect 1946 5720 1952 5723
rect 2004 5720 2010 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4080 5769 4108 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 8297 5831 8355 5837
rect 8297 5797 8309 5831
rect 8343 5828 8355 5831
rect 8386 5828 8392 5840
rect 8343 5800 8392 5828
rect 8343 5797 8355 5800
rect 8297 5791 8355 5797
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4321 5763 4379 5769
rect 4321 5760 4333 5763
rect 4212 5732 4333 5760
rect 4212 5720 4218 5732
rect 4321 5729 4333 5732
rect 4367 5729 4379 5763
rect 4321 5723 4379 5729
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 6724 5763 6782 5769
rect 6724 5760 6736 5763
rect 6328 5732 6736 5760
rect 6328 5720 6334 5732
rect 6724 5729 6736 5732
rect 6770 5760 6782 5763
rect 8202 5760 8208 5772
rect 6770 5732 8208 5760
rect 6770 5729 6782 5732
rect 6724 5723 6782 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 8956 5760 8984 5859
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 9088 5868 9137 5896
rect 9088 5856 9094 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 10321 5899 10379 5905
rect 10321 5896 10333 5899
rect 9548 5868 10333 5896
rect 9548 5856 9554 5868
rect 10321 5865 10333 5868
rect 10367 5865 10379 5899
rect 11974 5896 11980 5908
rect 11935 5868 11980 5896
rect 10321 5859 10379 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13357 5899 13415 5905
rect 13357 5896 13369 5899
rect 13044 5868 13369 5896
rect 13044 5856 13050 5868
rect 13357 5865 13369 5868
rect 13403 5865 13415 5899
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 13357 5859 13415 5865
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8956 5732 9321 5760
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 11882 5760 11888 5772
rect 11572 5732 11888 5760
rect 11572 5720 11578 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 13372 5760 13400 5859
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14093 5899 14151 5905
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14642 5896 14648 5908
rect 14139 5868 14648 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14642 5856 14648 5868
rect 14700 5896 14706 5908
rect 15010 5896 15016 5908
rect 14700 5868 15016 5896
rect 14700 5856 14706 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15286 5896 15292 5908
rect 15151 5868 15292 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 17034 5896 17040 5908
rect 16995 5868 17040 5896
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 20901 5899 20959 5905
rect 20901 5865 20913 5899
rect 20947 5896 20959 5899
rect 21266 5896 21272 5908
rect 20947 5868 21272 5896
rect 20947 5865 20959 5868
rect 20901 5859 20959 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 22373 5899 22431 5905
rect 22373 5865 22385 5899
rect 22419 5896 22431 5899
rect 22462 5896 22468 5908
rect 22419 5868 22468 5896
rect 22419 5865 22431 5868
rect 22373 5859 22431 5865
rect 22462 5856 22468 5868
rect 22520 5896 22526 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 22520 5868 24041 5896
rect 22520 5856 22526 5868
rect 24029 5865 24041 5868
rect 24075 5865 24087 5899
rect 24029 5859 24087 5865
rect 24118 5856 24124 5908
rect 24176 5896 24182 5908
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 24176 5868 25053 5896
rect 24176 5856 24182 5868
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25041 5859 25099 5865
rect 25130 5856 25136 5908
rect 25188 5896 25194 5908
rect 25409 5899 25467 5905
rect 25409 5896 25421 5899
rect 25188 5868 25421 5896
rect 25188 5856 25194 5868
rect 25409 5865 25421 5868
rect 25455 5865 25467 5899
rect 25409 5859 25467 5865
rect 25682 5856 25688 5908
rect 25740 5896 25746 5908
rect 25777 5899 25835 5905
rect 25777 5896 25789 5899
rect 25740 5868 25789 5896
rect 25740 5856 25746 5868
rect 25777 5865 25789 5868
rect 25823 5865 25835 5899
rect 25777 5859 25835 5865
rect 14366 5788 14372 5840
rect 14424 5828 14430 5840
rect 15534 5831 15592 5837
rect 15534 5828 15546 5831
rect 14424 5800 15546 5828
rect 14424 5788 14430 5800
rect 15534 5797 15546 5800
rect 15580 5797 15592 5831
rect 15534 5791 15592 5797
rect 20530 5788 20536 5840
rect 20588 5828 20594 5840
rect 20588 5800 22968 5828
rect 20588 5788 20594 5800
rect 22940 5772 22968 5800
rect 23658 5788 23664 5840
rect 23716 5828 23722 5840
rect 24397 5831 24455 5837
rect 24397 5828 24409 5831
rect 23716 5800 24409 5828
rect 23716 5788 23722 5800
rect 24397 5797 24409 5800
rect 24443 5828 24455 5831
rect 24854 5828 24860 5840
rect 24443 5800 24860 5828
rect 24443 5797 24455 5800
rect 24397 5791 24455 5797
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 13630 5760 13636 5772
rect 13372 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17451 5732 17785 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 17773 5729 17785 5732
rect 17819 5760 17831 5763
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 17819 5732 18337 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 18325 5729 18337 5732
rect 18371 5760 18383 5763
rect 18414 5760 18420 5772
rect 18371 5732 18420 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 18414 5720 18420 5732
rect 18472 5720 18478 5772
rect 18598 5769 18604 5772
rect 18592 5760 18604 5769
rect 18559 5732 18604 5760
rect 18592 5723 18604 5732
rect 18598 5720 18604 5723
rect 18656 5720 18662 5772
rect 21266 5760 21272 5772
rect 21227 5732 21272 5760
rect 21266 5720 21272 5732
rect 21324 5760 21330 5772
rect 21913 5763 21971 5769
rect 21913 5760 21925 5763
rect 21324 5732 21925 5760
rect 21324 5720 21330 5732
rect 21913 5729 21925 5732
rect 21959 5729 21971 5763
rect 21913 5723 21971 5729
rect 22370 5720 22376 5772
rect 22428 5760 22434 5772
rect 22738 5760 22744 5772
rect 22428 5732 22744 5760
rect 22428 5720 22434 5732
rect 22738 5720 22744 5732
rect 22796 5760 22802 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 22796 5732 22845 5760
rect 22796 5720 22802 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 22922 5720 22928 5772
rect 22980 5760 22986 5772
rect 26142 5760 26148 5772
rect 22980 5732 26148 5760
rect 22980 5720 22986 5732
rect 26142 5720 26148 5732
rect 26200 5720 26206 5772
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 6457 5695 6515 5701
rect 6457 5692 6469 5695
rect 5132 5664 6469 5692
rect 5132 5652 5138 5664
rect 6457 5661 6469 5664
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3050 5556 3056 5568
rect 2832 5528 3056 5556
rect 2832 5516 2838 5528
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6178 5556 6184 5568
rect 5859 5528 6184 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6472 5556 6500 5655
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 9824 5664 10425 5692
rect 9824 5652 9830 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10778 5692 10784 5704
rect 10643 5664 10784 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12124 5664 12541 5692
rect 12124 5652 12130 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 14182 5692 14188 5704
rect 14143 5664 14188 5692
rect 12529 5655 12587 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14642 5692 14648 5704
rect 14603 5664 14648 5692
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 21358 5692 21364 5704
rect 20763 5664 21364 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 9950 5624 9956 5636
rect 9911 5596 9956 5624
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 11054 5584 11060 5636
rect 11112 5624 11118 5636
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 11112 5596 11529 5624
rect 11112 5584 11118 5596
rect 11517 5593 11529 5596
rect 11563 5593 11575 5627
rect 11517 5587 11575 5593
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12952 5596 13093 5624
rect 12952 5584 12958 5596
rect 13081 5593 13093 5596
rect 13127 5624 13139 5627
rect 14200 5624 14228 5652
rect 13127 5596 14228 5624
rect 13127 5593 13139 5596
rect 13081 5587 13139 5593
rect 6730 5556 6736 5568
rect 6472 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5556 6794 5568
rect 7098 5556 7104 5568
rect 6788 5528 7104 5556
rect 6788 5516 6794 5528
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 10965 5559 11023 5565
rect 10965 5525 10977 5559
rect 11011 5556 11023 5559
rect 11146 5556 11152 5568
rect 11011 5528 11152 5556
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11146 5516 11152 5528
rect 11204 5556 11210 5568
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 11204 5528 11437 5556
rect 11204 5516 11210 5528
rect 11425 5525 11437 5528
rect 11471 5556 11483 5559
rect 11790 5556 11796 5568
rect 11471 5528 11796 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 15304 5556 15332 5655
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 23106 5692 23112 5704
rect 23067 5664 23112 5692
rect 21453 5655 21511 5661
rect 21468 5624 21496 5655
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 23624 5664 24501 5692
rect 23624 5652 23630 5664
rect 24489 5661 24501 5664
rect 24535 5661 24547 5695
rect 24670 5692 24676 5704
rect 24583 5664 24676 5692
rect 24489 5655 24547 5661
rect 20088 5596 21496 5624
rect 24504 5624 24532 5655
rect 24670 5652 24676 5664
rect 24728 5692 24734 5704
rect 24946 5692 24952 5704
rect 24728 5664 24952 5692
rect 24728 5652 24734 5664
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 25406 5624 25412 5636
rect 24504 5596 25412 5624
rect 20088 5568 20116 5596
rect 25406 5584 25412 5596
rect 25464 5584 25470 5636
rect 15562 5556 15568 5568
rect 15304 5528 15568 5556
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 16666 5556 16672 5568
rect 16627 5528 16672 5556
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 18233 5559 18291 5565
rect 18233 5525 18245 5559
rect 18279 5556 18291 5559
rect 18506 5556 18512 5568
rect 18279 5528 18512 5556
rect 18279 5525 18291 5528
rect 18233 5519 18291 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 20070 5556 20076 5568
rect 20031 5528 20076 5556
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 22465 5559 22523 5565
rect 22465 5525 22477 5559
rect 22511 5556 22523 5559
rect 23382 5556 23388 5568
rect 22511 5528 23388 5556
rect 22511 5525 22523 5528
rect 22465 5519 22523 5525
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 23658 5556 23664 5568
rect 23619 5528 23664 5556
rect 23658 5516 23664 5528
rect 23716 5516 23722 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2590 5312 2596 5364
rect 2648 5352 2654 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 2648 5324 3709 5352
rect 2648 5312 2654 5324
rect 3697 5321 3709 5324
rect 3743 5352 3755 5355
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 3743 5324 4353 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4341 5321 4353 5324
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 5994 5352 6000 5364
rect 5951 5324 6000 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 4065 5287 4123 5293
rect 4065 5253 4077 5287
rect 4111 5284 4123 5287
rect 4154 5284 4160 5296
rect 4111 5256 4160 5284
rect 4111 5253 4123 5256
rect 4065 5247 4123 5253
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 1728 5188 2329 5216
rect 1728 5176 1734 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 4356 5216 4384 5315
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6270 5352 6276 5364
rect 6231 5324 6276 5352
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 7248 5324 7297 5352
rect 7248 5312 7254 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 7285 5315 7343 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10778 5352 10784 5364
rect 10739 5324 10784 5352
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 12032 5324 12173 5352
rect 12032 5312 12038 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12161 5315 12219 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 13814 5352 13820 5364
rect 13403 5324 13820 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14424 5324 14933 5352
rect 14424 5312 14430 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 15838 5352 15844 5364
rect 15795 5324 15844 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16724 5324 16865 5352
rect 16724 5312 16730 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 16853 5315 16911 5321
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18693 5355 18751 5361
rect 18693 5352 18705 5355
rect 18656 5324 18705 5352
rect 18656 5312 18662 5324
rect 18693 5321 18705 5324
rect 18739 5352 18751 5355
rect 20622 5352 20628 5364
rect 18739 5324 20628 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 21358 5312 21364 5364
rect 21416 5352 21422 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21416 5324 21557 5352
rect 21416 5312 21422 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 21545 5315 21603 5321
rect 22738 5312 22744 5364
rect 22796 5352 22802 5364
rect 22925 5355 22983 5361
rect 22925 5352 22937 5355
rect 22796 5324 22937 5352
rect 22796 5312 22802 5324
rect 22925 5321 22937 5324
rect 22971 5321 22983 5355
rect 22925 5315 22983 5321
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 23293 5355 23351 5361
rect 23293 5352 23305 5355
rect 23164 5324 23305 5352
rect 23164 5312 23170 5324
rect 23293 5321 23305 5324
rect 23339 5321 23351 5355
rect 23293 5315 23351 5321
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25041 5355 25099 5361
rect 25041 5352 25053 5355
rect 25004 5324 25053 5352
rect 25004 5312 25010 5324
rect 25041 5321 25053 5324
rect 25087 5352 25099 5355
rect 25317 5355 25375 5361
rect 25317 5352 25329 5355
rect 25087 5324 25329 5352
rect 25087 5321 25099 5324
rect 25041 5315 25099 5321
rect 25317 5321 25329 5324
rect 25363 5321 25375 5355
rect 25317 5315 25375 5321
rect 25406 5312 25412 5364
rect 25464 5352 25470 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 25464 5324 25697 5352
rect 25464 5312 25470 5324
rect 25685 5321 25697 5324
rect 25731 5321 25743 5355
rect 25685 5315 25743 5321
rect 25774 5312 25780 5364
rect 25832 5352 25838 5364
rect 26053 5355 26111 5361
rect 26053 5352 26065 5355
rect 25832 5324 26065 5352
rect 25832 5312 25838 5324
rect 26053 5321 26065 5324
rect 26099 5321 26111 5355
rect 26053 5315 26111 5321
rect 6178 5244 6184 5296
rect 6236 5284 6242 5296
rect 6454 5284 6460 5296
rect 6236 5256 6460 5284
rect 6236 5244 6242 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6641 5219 6699 5225
rect 4356 5188 4660 5216
rect 2317 5179 2375 5185
rect 2332 5148 2360 5179
rect 2866 5148 2872 5160
rect 2332 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5117 4583 5151
rect 4632 5148 4660 5188
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7558 5216 7564 5228
rect 6687 5188 7564 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 7558 5176 7564 5188
rect 7616 5216 7622 5228
rect 7742 5216 7748 5228
rect 7616 5188 7748 5216
rect 7616 5176 7622 5188
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 8312 5216 8340 5312
rect 9677 5287 9735 5293
rect 9677 5253 9689 5287
rect 9723 5284 9735 5287
rect 10134 5284 10140 5296
rect 9723 5256 10140 5284
rect 9723 5253 9735 5256
rect 9677 5247 9735 5253
rect 10134 5244 10140 5256
rect 10192 5284 10198 5296
rect 14461 5287 14519 5293
rect 10192 5256 10364 5284
rect 10192 5244 10198 5256
rect 10336 5225 10364 5256
rect 14461 5253 14473 5287
rect 14507 5284 14519 5287
rect 15286 5284 15292 5296
rect 14507 5256 15292 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 7975 5188 8340 5216
rect 10321 5219 10379 5225
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 12250 5216 12256 5228
rect 11379 5188 12256 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13688 5188 13829 5216
rect 13688 5176 13694 5188
rect 13817 5185 13829 5188
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14182 5216 14188 5228
rect 14047 5188 14188 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 15856 5216 15884 5312
rect 16298 5216 16304 5228
rect 15856 5188 16304 5216
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5216 16543 5219
rect 16684 5216 16712 5312
rect 17586 5244 17592 5296
rect 17644 5284 17650 5296
rect 18233 5287 18291 5293
rect 18233 5284 18245 5287
rect 17644 5256 18245 5284
rect 17644 5244 17650 5256
rect 18233 5253 18245 5256
rect 18279 5253 18291 5287
rect 23658 5284 23664 5296
rect 18233 5247 18291 5253
rect 23492 5256 23664 5284
rect 16531 5188 16712 5216
rect 19153 5219 19211 5225
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 19153 5185 19165 5219
rect 19199 5216 19211 5219
rect 19199 5188 19380 5216
rect 19199 5185 19211 5188
rect 19153 5179 19211 5185
rect 4781 5151 4839 5157
rect 4781 5148 4793 5151
rect 4632 5120 4793 5148
rect 4525 5111 4583 5117
rect 4781 5117 4793 5120
rect 4827 5117 4839 5151
rect 4781 5111 4839 5117
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9355 5120 10241 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10962 5148 10968 5160
rect 10275 5120 10968 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 2590 5089 2596 5092
rect 2584 5080 2596 5089
rect 2551 5052 2596 5080
rect 2584 5043 2596 5052
rect 2590 5040 2596 5043
rect 2648 5040 2654 5092
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 4540 5080 4568 5111
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 15381 5151 15439 5157
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 15427 5120 16221 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 16209 5117 16221 5120
rect 16255 5148 16267 5151
rect 16390 5148 16396 5160
rect 16255 5120 16396 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17788 5120 18061 5148
rect 17788 5092 17816 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5117 19303 5151
rect 19352 5148 19380 5188
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22649 5219 22707 5225
rect 22152 5188 22197 5216
rect 22152 5176 22158 5188
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 22922 5216 22928 5228
rect 22695 5188 22928 5216
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 22922 5176 22928 5188
rect 22980 5176 22986 5228
rect 19512 5151 19570 5157
rect 19512 5148 19524 5151
rect 19352 5120 19524 5148
rect 19245 5111 19303 5117
rect 19512 5117 19524 5120
rect 19558 5148 19570 5151
rect 20070 5148 20076 5160
rect 19558 5120 20076 5148
rect 19558 5117 19570 5120
rect 19512 5111 19570 5117
rect 5074 5080 5080 5092
rect 4120 5052 5080 5080
rect 4120 5040 4126 5052
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 8941 5083 8999 5089
rect 8941 5049 8953 5083
rect 8987 5080 8999 5083
rect 9858 5080 9864 5092
rect 8987 5052 9864 5080
rect 8987 5049 8999 5052
rect 8941 5043 8999 5049
rect 9858 5040 9864 5052
rect 9916 5080 9922 5092
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 9916 5052 10149 5080
rect 9916 5040 9922 5052
rect 10137 5049 10149 5052
rect 10183 5049 10195 5083
rect 10137 5043 10195 5049
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 11793 5083 11851 5089
rect 11793 5080 11805 5083
rect 11112 5052 11805 5080
rect 11112 5040 11118 5052
rect 11793 5049 11805 5052
rect 11839 5080 11851 5083
rect 11882 5080 11888 5092
rect 11839 5052 11888 5080
rect 11839 5049 11851 5052
rect 11793 5043 11851 5049
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 13262 5080 13268 5092
rect 13175 5052 13268 5080
rect 13262 5040 13268 5052
rect 13320 5080 13326 5092
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 13320 5052 13737 5080
rect 13320 5040 13326 5052
rect 13725 5049 13737 5052
rect 13771 5080 13783 5083
rect 17770 5080 17776 5092
rect 13771 5052 16436 5080
rect 17731 5052 17776 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 16408 5024 16436 5052
rect 17770 5040 17776 5052
rect 17828 5040 17834 5092
rect 19150 5040 19156 5092
rect 19208 5080 19214 5092
rect 19260 5080 19288 5111
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5148 21143 5151
rect 21910 5148 21916 5160
rect 21131 5120 21916 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 23290 5108 23296 5160
rect 23348 5148 23354 5160
rect 23492 5148 23520 5256
rect 23658 5244 23664 5256
rect 23716 5244 23722 5296
rect 23348 5120 23520 5148
rect 23348 5108 23354 5120
rect 19208 5052 19288 5080
rect 23492 5080 23520 5120
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 25682 5148 25688 5160
rect 23707 5120 25688 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 25682 5108 25688 5120
rect 25740 5108 25746 5160
rect 23906 5083 23964 5089
rect 23906 5080 23918 5083
rect 23492 5052 23918 5080
rect 19208 5040 19214 5052
rect 23906 5049 23918 5052
rect 23952 5049 23964 5083
rect 23906 5043 23964 5049
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 1946 5012 1952 5024
rect 1719 4984 1952 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 1946 4972 1952 4984
rect 2004 5012 2010 5024
rect 2041 5015 2099 5021
rect 2041 5012 2053 5015
rect 2004 4984 2053 5012
rect 2004 4972 2010 4984
rect 2041 4981 2053 4984
rect 2087 5012 2099 5015
rect 2222 5012 2228 5024
rect 2087 4984 2228 5012
rect 2087 4981 2099 4984
rect 2041 4975 2099 4981
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 7193 5015 7251 5021
rect 7193 4981 7205 5015
rect 7239 5012 7251 5015
rect 7650 5012 7656 5024
rect 7239 4984 7656 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10962 5012 10968 5024
rect 9640 4984 10968 5012
rect 9640 4972 9646 4984
rect 10962 4972 10968 4984
rect 11020 5012 11026 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 11020 4984 11161 5012
rect 11020 4972 11026 4984
rect 11149 4981 11161 4984
rect 11195 5012 11207 5015
rect 12066 5012 12072 5024
rect 11195 4984 12072 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 15841 5015 15899 5021
rect 15841 4981 15853 5015
rect 15887 5012 15899 5015
rect 16114 5012 16120 5024
rect 15887 4984 16120 5012
rect 15887 4981 15899 4984
rect 15841 4975 15899 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16390 4972 16396 5024
rect 16448 4972 16454 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 21453 5015 21511 5021
rect 21453 4981 21465 5015
rect 21499 5012 21511 5015
rect 22005 5015 22063 5021
rect 22005 5012 22017 5015
rect 21499 4984 22017 5012
rect 21499 4981 21511 4984
rect 21453 4975 21511 4981
rect 22005 4981 22017 4984
rect 22051 5012 22063 5015
rect 22738 5012 22744 5024
rect 22051 4984 22744 5012
rect 22051 4981 22063 4984
rect 22005 4975 22063 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 24762 4972 24768 5024
rect 24820 5012 24826 5024
rect 25406 5012 25412 5024
rect 24820 4984 25412 5012
rect 24820 4972 24826 4984
rect 25406 4972 25412 4984
rect 25464 4972 25470 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4982 4808 4988 4820
rect 4943 4780 4988 4808
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 5224 4780 5365 4808
rect 5224 4768 5230 4780
rect 5353 4777 5365 4780
rect 5399 4808 5411 4811
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5399 4780 6009 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7374 4808 7380 4820
rect 6696 4780 7380 4808
rect 6696 4768 6702 4780
rect 7374 4768 7380 4780
rect 7432 4808 7438 4820
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7432 4780 7481 4808
rect 7432 4768 7438 4780
rect 7469 4777 7481 4780
rect 7515 4777 7527 4811
rect 7469 4771 7527 4777
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9766 4808 9772 4820
rect 9539 4780 9772 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 11020 4780 11069 4808
rect 11020 4768 11026 4780
rect 11057 4777 11069 4780
rect 11103 4777 11115 4811
rect 11057 4771 11115 4777
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12710 4808 12716 4820
rect 12207 4780 12716 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14274 4808 14280 4820
rect 14235 4780 14280 4808
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 17862 4808 17868 4820
rect 17819 4780 17868 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 20070 4768 20076 4820
rect 20128 4808 20134 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20128 4780 20637 4808
rect 20128 4768 20134 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 22002 4808 22008 4820
rect 21963 4780 22008 4808
rect 20625 4771 20683 4777
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 22925 4811 22983 4817
rect 22925 4777 22937 4811
rect 22971 4808 22983 4811
rect 23014 4808 23020 4820
rect 22971 4780 23020 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 1854 4700 1860 4752
rect 1912 4740 1918 4752
rect 10042 4740 10048 4752
rect 1912 4712 2084 4740
rect 1912 4700 1918 4712
rect 658 4632 664 4684
rect 716 4672 722 4684
rect 1578 4672 1584 4684
rect 716 4644 1584 4672
rect 716 4632 722 4644
rect 1578 4632 1584 4644
rect 1636 4672 1642 4684
rect 1762 4672 1768 4684
rect 1636 4644 1768 4672
rect 1636 4632 1642 4644
rect 1762 4632 1768 4644
rect 1820 4672 1826 4684
rect 2056 4681 2084 4712
rect 9692 4712 10048 4740
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1820 4644 1961 4672
rect 1820 4632 1826 4644
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 1949 4635 2007 4641
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4672 2099 4675
rect 2406 4672 2412 4684
rect 2087 4644 2412 4672
rect 2087 4641 2099 4644
rect 2041 4635 2099 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4982 4672 4988 4684
rect 4479 4644 4988 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5592 4644 5917 4672
rect 5592 4632 5598 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 8018 4672 8024 4684
rect 7607 4644 8024 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9490 4672 9496 4684
rect 9171 4644 9496 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 9692 4681 9720 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 12434 4740 12440 4752
rect 12400 4712 12440 4740
rect 12400 4700 12406 4712
rect 12434 4700 12440 4712
rect 12492 4749 12498 4752
rect 12492 4743 12556 4749
rect 12492 4709 12510 4743
rect 12544 4740 12556 4743
rect 12544 4712 12585 4740
rect 12544 4709 12556 4712
rect 12492 4703 12556 4709
rect 12492 4700 12498 4703
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 15832 4743 15890 4749
rect 15832 4740 15844 4743
rect 15436 4712 15844 4740
rect 15436 4700 15442 4712
rect 15832 4709 15844 4712
rect 15878 4740 15890 4743
rect 16022 4740 16028 4752
rect 15878 4712 16028 4740
rect 15878 4709 15890 4712
rect 15832 4703 15890 4709
rect 16022 4700 16028 4712
rect 16080 4740 16086 4752
rect 16666 4740 16672 4752
rect 16080 4712 16672 4740
rect 16080 4700 16086 4712
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 19613 4743 19671 4749
rect 19613 4740 19625 4743
rect 19484 4712 19625 4740
rect 19484 4700 19490 4712
rect 19613 4709 19625 4712
rect 19659 4709 19671 4743
rect 19613 4703 19671 4709
rect 21910 4700 21916 4752
rect 21968 4740 21974 4752
rect 22940 4740 22968 4771
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 23474 4768 23480 4820
rect 23532 4808 23538 4820
rect 23658 4808 23664 4820
rect 23532 4780 23664 4808
rect 23532 4768 23538 4780
rect 23658 4768 23664 4780
rect 23716 4768 23722 4820
rect 24854 4768 24860 4820
rect 24912 4808 24918 4820
rect 25041 4811 25099 4817
rect 25041 4808 25053 4811
rect 24912 4780 25053 4808
rect 24912 4768 24918 4780
rect 25041 4777 25053 4780
rect 25087 4777 25099 4811
rect 25041 4771 25099 4777
rect 25501 4811 25559 4817
rect 25501 4777 25513 4811
rect 25547 4808 25559 4811
rect 25682 4808 25688 4820
rect 25547 4780 25688 4808
rect 25547 4777 25559 4780
rect 25501 4771 25559 4777
rect 25682 4768 25688 4780
rect 25740 4768 25746 4820
rect 21968 4712 22968 4740
rect 21968 4700 21974 4712
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9944 4675 10002 4681
rect 9944 4641 9956 4675
rect 9990 4672 10002 4675
rect 10778 4672 10784 4684
rect 9990 4644 10784 4672
rect 9990 4641 10002 4644
rect 9944 4635 10002 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 15562 4672 15568 4684
rect 15523 4644 15568 4672
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 17494 4672 17500 4684
rect 16356 4644 17500 4672
rect 16356 4632 16362 4644
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 18012 4644 18153 4672
rect 18012 4632 18018 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 19334 4672 19340 4684
rect 19295 4644 19340 4672
rect 18141 4635 18199 4641
rect 19334 4632 19340 4644
rect 19392 4672 19398 4684
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 19392 4644 20085 4672
rect 19392 4632 19398 4644
rect 20073 4641 20085 4644
rect 20119 4641 20131 4675
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 20073 4635 20131 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 22833 4675 22891 4681
rect 22833 4641 22845 4675
rect 22879 4672 22891 4675
rect 23198 4672 23204 4684
rect 22879 4644 23204 4672
rect 22879 4641 22891 4644
rect 22833 4635 22891 4641
rect 23198 4632 23204 4644
rect 23256 4632 23262 4684
rect 23474 4632 23480 4684
rect 23532 4672 23538 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23532 4644 24409 4672
rect 23532 4632 23538 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5408 4576 6193 4604
rect 5408 4564 5414 4576
rect 6181 4573 6193 4576
rect 6227 4604 6239 4607
rect 7742 4604 7748 4616
rect 6227 4576 7748 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 12250 4604 12256 4616
rect 12211 4576 12256 4604
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4604 18475 4607
rect 18506 4604 18512 4616
rect 18463 4576 18512 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 18506 4564 18512 4576
rect 18564 4604 18570 4616
rect 19150 4604 19156 4616
rect 18564 4576 19156 4604
rect 18564 4564 18570 4576
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 21174 4564 21180 4616
rect 21232 4604 21238 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21232 4576 21373 4604
rect 21232 4564 21238 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 3605 4539 3663 4545
rect 3605 4536 3617 4539
rect 1964 4508 3617 4536
rect 1964 4480 1992 4508
rect 3605 4505 3617 4508
rect 3651 4505 3663 4539
rect 3605 4499 3663 4505
rect 20806 4496 20812 4548
rect 20864 4536 20870 4548
rect 21468 4536 21496 4567
rect 22370 4536 22376 4548
rect 20864 4508 21496 4536
rect 22283 4508 22376 4536
rect 20864 4496 20870 4508
rect 22370 4496 22376 4508
rect 22428 4536 22434 4548
rect 23032 4536 23060 4567
rect 24118 4564 24124 4616
rect 24176 4604 24182 4616
rect 24489 4607 24547 4613
rect 24489 4604 24501 4607
rect 24176 4576 24501 4604
rect 24176 4564 24182 4576
rect 24489 4573 24501 4576
rect 24535 4573 24547 4607
rect 24489 4567 24547 4573
rect 24578 4564 24584 4616
rect 24636 4604 24642 4616
rect 24854 4604 24860 4616
rect 24636 4576 24860 4604
rect 24636 4564 24642 4576
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 22428 4508 23060 4536
rect 22428 4496 22434 4508
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 1946 4468 1952 4480
rect 1627 4440 1952 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 2590 4468 2596 4480
rect 2551 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3510 4468 3516 4480
rect 3375 4440 3516 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 6178 4468 6184 4480
rect 5583 4440 6184 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6914 4468 6920 4480
rect 6604 4440 6920 4468
rect 6604 4428 6610 4440
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7098 4468 7104 4480
rect 7059 4440 7104 4468
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 8662 4468 8668 4480
rect 8623 4440 8668 4468
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 11790 4468 11796 4480
rect 11471 4440 11796 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 13630 4468 13636 4480
rect 13591 4440 13636 4468
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15105 4471 15163 4477
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 15286 4468 15292 4480
rect 15151 4440 15292 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16540 4440 16957 4468
rect 16540 4428 16546 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 17310 4468 17316 4480
rect 17223 4440 17316 4468
rect 16945 4431 17003 4437
rect 17310 4428 17316 4440
rect 17368 4468 17374 4480
rect 17678 4468 17684 4480
rect 17368 4440 17684 4468
rect 17368 4428 17374 4440
rect 17678 4428 17684 4440
rect 17736 4428 17742 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 18877 4471 18935 4477
rect 18877 4468 18889 4471
rect 18472 4440 18889 4468
rect 18472 4428 18478 4440
rect 18877 4437 18889 4440
rect 18923 4468 18935 4471
rect 19058 4468 19064 4480
rect 18923 4440 19064 4468
rect 18923 4437 18935 4440
rect 18877 4431 18935 4437
rect 19058 4428 19064 4440
rect 19116 4468 19122 4480
rect 19153 4471 19211 4477
rect 19153 4468 19165 4471
rect 19116 4440 19165 4468
rect 19116 4428 19122 4440
rect 19153 4437 19165 4440
rect 19199 4437 19211 4471
rect 19153 4431 19211 4437
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 20901 4471 20959 4477
rect 20901 4468 20913 4471
rect 20772 4440 20913 4468
rect 20772 4428 20778 4440
rect 20901 4437 20913 4440
rect 20947 4437 20959 4471
rect 22462 4468 22468 4480
rect 22423 4440 22468 4468
rect 20901 4431 20959 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 24026 4468 24032 4480
rect 23987 4440 24032 4468
rect 24026 4428 24032 4440
rect 24084 4428 24090 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1486 4264 1492 4276
rect 1447 4236 1492 4264
rect 1486 4224 1492 4236
rect 1544 4224 1550 4276
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 2869 4267 2927 4273
rect 2869 4264 2881 4267
rect 1820 4236 2881 4264
rect 1820 4224 1826 4236
rect 2869 4233 2881 4236
rect 2915 4233 2927 4267
rect 2869 4227 2927 4233
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 4154 4264 4160 4276
rect 3108 4236 4160 4264
rect 3108 4224 3114 4236
rect 4154 4224 4160 4236
rect 4212 4264 4218 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 4212 4236 4629 4264
rect 4212 4224 4218 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 4982 4264 4988 4276
rect 4943 4236 4988 4264
rect 4617 4227 4675 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 6052 4236 6193 4264
rect 6052 4224 6058 4236
rect 6181 4233 6193 4236
rect 6227 4264 6239 4267
rect 6227 4236 7420 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 6825 4199 6883 4205
rect 6825 4196 6837 4199
rect 5592 4168 6837 4196
rect 5592 4156 5598 4168
rect 6825 4165 6837 4168
rect 6871 4165 6883 4199
rect 6825 4159 6883 4165
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2590 4128 2596 4140
rect 2179 4100 2596 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6270 4128 6276 4140
rect 5767 4100 6276 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 7392 4137 7420 4236
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7800 4236 8217 4264
rect 7800 4224 7806 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 9858 4264 9864 4276
rect 9819 4236 9864 4264
rect 8205 4227 8263 4233
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10836 4236 10885 4264
rect 10836 4224 10842 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 10873 4227 10931 4233
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 11020 4236 11253 4264
rect 11020 4224 11026 4236
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 11241 4227 11299 4233
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 15654 4264 15660 4276
rect 15615 4236 15660 4264
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 22741 4267 22799 4273
rect 22741 4233 22753 4267
rect 22787 4264 22799 4267
rect 23014 4264 23020 4276
rect 22787 4236 23020 4264
rect 22787 4233 22799 4236
rect 22741 4227 22799 4233
rect 23014 4224 23020 4236
rect 23072 4224 23078 4276
rect 23474 4264 23480 4276
rect 23435 4236 23480 4264
rect 23474 4224 23480 4236
rect 23532 4224 23538 4276
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24673 4267 24731 4273
rect 24673 4264 24685 4267
rect 24176 4236 24685 4264
rect 24176 4224 24182 4236
rect 24673 4233 24685 4236
rect 24719 4233 24731 4267
rect 24673 4227 24731 4233
rect 10980 4196 11008 4224
rect 10520 4168 11008 4196
rect 10520 4137 10548 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 10505 4091 10563 4097
rect 12912 4100 13001 4128
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 2924 4032 3249 4060
rect 2924 4020 2930 4032
rect 3237 4029 3249 4032
rect 3283 4060 3295 4063
rect 3326 4060 3332 4072
rect 3283 4032 3332 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3326 4020 3332 4032
rect 3384 4060 3390 4072
rect 4062 4060 4068 4072
rect 3384 4032 4068 4060
rect 3384 4020 3390 4032
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 5442 4060 5448 4072
rect 5355 4032 5448 4060
rect 5442 4020 5448 4032
rect 5500 4060 5506 4072
rect 6362 4060 6368 4072
rect 5500 4032 6368 4060
rect 5500 4020 5506 4032
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4060 6610 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6604 4032 7297 4060
rect 6604 4020 6610 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8018 4060 8024 4072
rect 7975 4032 8024 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4060 8631 4063
rect 8662 4060 8668 4072
rect 8619 4032 8668 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 8662 4020 8668 4032
rect 8720 4060 8726 4072
rect 9582 4060 9588 4072
rect 8720 4032 9588 4060
rect 8720 4020 8726 4032
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9692 4032 10241 4060
rect 3510 4001 3516 4004
rect 3504 3992 3516 4001
rect 3471 3964 3516 3992
rect 3504 3955 3516 3964
rect 3510 3952 3516 3955
rect 3568 3952 3574 4004
rect 8849 3995 8907 4001
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 9030 3992 9036 4004
rect 8895 3964 9036 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9692 3992 9720 4032
rect 10229 4029 10241 4032
rect 10275 4060 10287 4063
rect 10778 4060 10784 4072
rect 10275 4032 10784 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4060 12311 4063
rect 12342 4060 12348 4072
rect 12299 4032 12348 4060
rect 12299 4029 12311 4032
rect 12253 4023 12311 4029
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12768 4032 12817 4060
rect 12768 4020 12774 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 9324 3964 9720 3992
rect 9876 3964 10333 3992
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 2464 3896 2513 3924
rect 2464 3884 2470 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 6972 3896 7205 3924
rect 6972 3884 6978 3896
rect 7193 3893 7205 3896
rect 7239 3924 7251 3927
rect 8662 3924 8668 3936
rect 7239 3896 8668 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9324 3933 9352 3964
rect 9876 3936 9904 3964
rect 10321 3961 10333 3964
rect 10367 3992 10379 3995
rect 10686 3992 10692 4004
rect 10367 3964 10692 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 12912 3992 12940 4100
rect 12989 4097 13001 4100
rect 13035 4128 13047 4131
rect 13630 4128 13636 4140
rect 13035 4100 13636 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13630 4088 13636 4100
rect 13688 4128 13694 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13688 4100 13829 4128
rect 13688 4088 13694 4100
rect 13817 4097 13829 4100
rect 13863 4128 13875 4131
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 13863 4100 14565 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 15672 4128 15700 4224
rect 19150 4196 19156 4208
rect 19111 4168 19156 4196
rect 19150 4156 19156 4168
rect 19208 4156 19214 4208
rect 20254 4196 20260 4208
rect 19812 4168 20260 4196
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 15672 4100 16405 4128
rect 14553 4091 14611 4097
rect 16393 4097 16405 4100
rect 16439 4128 16451 4131
rect 16482 4128 16488 4140
rect 16439 4100 16488 4128
rect 16439 4097 16451 4100
rect 16393 4091 16451 4097
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17092 4100 17417 4128
rect 17092 4088 17098 4100
rect 17405 4097 17417 4100
rect 17451 4128 17463 4131
rect 17862 4128 17868 4140
rect 17451 4100 17868 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 19812 4128 19840 4168
rect 20254 4156 20260 4168
rect 20312 4156 20318 4208
rect 19260 4100 19840 4128
rect 19889 4131 19947 4137
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14332 4032 14381 4060
rect 14332 4020 14338 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 15344 4032 16313 4060
rect 15344 4020 15350 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 16816 4032 17785 4060
rect 16816 4020 16822 4032
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 12728 3964 12940 3992
rect 12728 3936 12756 3964
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 13044 3964 13461 3992
rect 13044 3952 13050 3964
rect 13449 3961 13461 3964
rect 13495 3992 13507 3995
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 13495 3964 14473 3992
rect 13495 3961 13507 3964
rect 13449 3955 13507 3961
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 16172 3964 16221 3992
rect 16172 3952 16178 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17037 3995 17095 4001
rect 17037 3992 17049 3995
rect 17000 3964 17049 3992
rect 17000 3952 17006 3964
rect 17037 3961 17049 3964
rect 17083 3961 17095 3995
rect 17788 3992 17816 4023
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18288 4032 18521 4060
rect 18288 4020 18294 4032
rect 18509 4029 18521 4032
rect 18555 4060 18567 4063
rect 18782 4060 18788 4072
rect 18555 4032 18788 4060
rect 18555 4029 18567 4032
rect 18509 4023 18567 4029
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 18417 3995 18475 4001
rect 18417 3992 18429 3995
rect 17788 3964 18429 3992
rect 17037 3955 17095 3961
rect 18417 3961 18429 3964
rect 18463 3992 18475 3995
rect 19260 3992 19288 4100
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20162 4128 20168 4140
rect 19935 4100 20168 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20496 4100 20545 4128
rect 20496 4088 20502 4100
rect 20533 4097 20545 4100
rect 20579 4128 20591 4131
rect 20806 4128 20812 4140
rect 20579 4100 20812 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 20990 4128 20996 4140
rect 20951 4100 20996 4128
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23164 4100 24225 4128
rect 23164 4088 23170 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 24912 4100 25053 4128
rect 24912 4088 24918 4100
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25498 4128 25504 4140
rect 25459 4100 25504 4128
rect 25041 4091 25099 4097
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 26329 4131 26387 4137
rect 26329 4128 26341 4131
rect 25740 4100 26341 4128
rect 25740 4088 25746 4100
rect 26329 4097 26341 4100
rect 26375 4097 26387 4131
rect 26329 4091 26387 4097
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 18463 3964 19288 3992
rect 19444 4032 19625 4060
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 19444 3936 19472 4032
rect 19613 4029 19625 4032
rect 19659 4029 19671 4063
rect 19613 4023 19671 4029
rect 23658 4020 23664 4072
rect 23716 4060 23722 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 23716 4032 24041 4060
rect 23716 4020 23722 4032
rect 24029 4029 24041 4032
rect 24075 4060 24087 4063
rect 24302 4060 24308 4072
rect 24075 4032 24308 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 24302 4020 24308 4032
rect 24360 4020 24366 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25590 4060 25596 4072
rect 25271 4032 25596 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25590 4020 25596 4032
rect 25648 4060 25654 4072
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25648 4032 25973 4060
rect 25648 4020 25654 4032
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 25961 4023 26019 4029
rect 20901 3995 20959 4001
rect 20901 3961 20913 3995
rect 20947 3992 20959 3995
rect 21260 3995 21318 4001
rect 21260 3992 21272 3995
rect 20947 3964 21272 3992
rect 20947 3961 20959 3964
rect 20901 3955 20959 3961
rect 21260 3961 21272 3964
rect 21306 3992 21318 3995
rect 22002 3992 22008 4004
rect 21306 3964 22008 3992
rect 21306 3961 21318 3964
rect 21260 3955 21318 3961
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 23290 3992 23296 4004
rect 22388 3964 23296 3992
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9272 3896 9321 3924
rect 9272 3884 9278 3896
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 9309 3887 9367 3893
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 9858 3924 9864 3936
rect 9815 3896 9864 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12710 3884 12716 3936
rect 12768 3884 12774 3936
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13998 3924 14004 3936
rect 13959 3896 14004 3924
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 19426 3924 19432 3936
rect 19387 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 22388 3933 22416 3964
rect 23290 3952 23296 3964
rect 23348 3952 23354 4004
rect 22373 3927 22431 3933
rect 22373 3893 22385 3927
rect 22419 3893 22431 3927
rect 22373 3887 22431 3893
rect 23109 3927 23167 3933
rect 23109 3893 23121 3927
rect 23155 3924 23167 3927
rect 23198 3924 23204 3936
rect 23155 3896 23204 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 23658 3924 23664 3936
rect 23619 3896 23664 3924
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 24118 3884 24124 3936
rect 24176 3924 24182 3936
rect 24176 3896 24221 3924
rect 24176 3884 24182 3896
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1489 3723 1547 3729
rect 1489 3689 1501 3723
rect 1535 3720 1547 3723
rect 1854 3720 1860 3732
rect 1535 3692 1860 3720
rect 1535 3689 1547 3692
rect 1489 3683 1547 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 2590 3720 2596 3732
rect 2551 3692 2596 3720
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4430 3720 4436 3732
rect 3936 3692 4436 3720
rect 3936 3680 3942 3692
rect 4430 3680 4436 3692
rect 4488 3720 4494 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 4488 3692 4537 3720
rect 4488 3680 4494 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5534 3720 5540 3732
rect 5215 3692 5540 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7742 3720 7748 3732
rect 7147 3692 7748 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 7926 3720 7932 3732
rect 7887 3692 7932 3720
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10962 3720 10968 3732
rect 10744 3692 10968 3720
rect 10744 3680 10750 3692
rect 10962 3680 10968 3692
rect 11020 3720 11026 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 11020 3692 11069 3720
rect 11020 3680 11026 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11514 3720 11520 3732
rect 11475 3692 11520 3720
rect 11057 3683 11115 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12434 3720 12440 3732
rect 12023 3692 12440 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12492 3692 12817 3720
rect 12492 3680 12498 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 13998 3720 14004 3732
rect 12943 3692 14004 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 1949 3655 2007 3661
rect 1949 3652 1961 3655
rect 1728 3624 1961 3652
rect 1728 3612 1734 3624
rect 1949 3621 1961 3624
rect 1995 3652 2007 3655
rect 2498 3652 2504 3664
rect 1995 3624 2504 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 2498 3612 2504 3624
rect 2556 3612 2562 3664
rect 5442 3652 5448 3664
rect 5403 3624 5448 3652
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5994 3661 6000 3664
rect 5988 3652 6000 3661
rect 5955 3624 6000 3652
rect 5988 3615 6000 3624
rect 5994 3612 6000 3615
rect 6052 3612 6058 3664
rect 7374 3652 7380 3664
rect 7335 3624 7380 3652
rect 7374 3612 7380 3624
rect 7432 3612 7438 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 7484 3624 8953 3652
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1854 3584 1860 3596
rect 1452 3556 1860 3584
rect 1452 3544 1458 3556
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 4430 3584 4436 3596
rect 4343 3556 4436 3584
rect 4430 3544 4436 3556
rect 4488 3584 4494 3596
rect 5258 3584 5264 3596
rect 4488 3556 5264 3584
rect 4488 3544 4494 3556
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 6730 3584 6736 3596
rect 5767 3556 6736 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2222 3516 2228 3528
rect 2179 3488 2228 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3467 3488 3893 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3881 3485 3893 3488
rect 3927 3516 3939 3519
rect 3970 3516 3976 3528
rect 3927 3488 3976 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 3970 3476 3976 3488
rect 4028 3516 4034 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4028 3488 4721 3516
rect 4028 3476 4034 3488
rect 4709 3485 4721 3488
rect 4755 3516 4767 3519
rect 5350 3516 5356 3528
rect 4755 3488 5356 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 2958 3448 2964 3460
rect 2871 3420 2964 3448
rect 2958 3408 2964 3420
rect 3016 3448 3022 3460
rect 3510 3448 3516 3460
rect 3016 3420 3516 3448
rect 3016 3408 3022 3420
rect 3510 3408 3516 3420
rect 3568 3408 3574 3460
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4065 3451 4123 3457
rect 4065 3448 4077 3451
rect 3844 3420 4077 3448
rect 3844 3408 3850 3420
rect 4065 3417 4077 3420
rect 4111 3448 4123 3451
rect 4111 3420 5304 3448
rect 4111 3417 4123 3420
rect 4065 3411 4123 3417
rect 5276 3380 5304 3420
rect 7484 3380 7512 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 10042 3652 10048 3664
rect 8941 3615 8999 3621
rect 9692 3624 10048 3652
rect 8294 3584 8300 3596
rect 8255 3556 8300 3584
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 9692 3593 9720 3624
rect 10042 3612 10048 3624
rect 10100 3652 10106 3664
rect 12250 3652 12256 3664
rect 10100 3624 12256 3652
rect 10100 3612 10106 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 12912 3652 12940 3683
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15344 3692 15485 3720
rect 15344 3680 15350 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15838 3720 15844 3732
rect 15799 3692 15844 3720
rect 15473 3683 15531 3689
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16172 3692 16865 3720
rect 16172 3680 16178 3692
rect 16853 3689 16865 3692
rect 16899 3689 16911 3723
rect 16853 3683 16911 3689
rect 18141 3723 18199 3729
rect 18141 3689 18153 3723
rect 18187 3720 18199 3723
rect 18230 3720 18236 3732
rect 18187 3692 18236 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 18598 3720 18604 3732
rect 18555 3692 18604 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19705 3723 19763 3729
rect 19705 3689 19717 3723
rect 19751 3720 19763 3723
rect 19978 3720 19984 3732
rect 19751 3692 19984 3720
rect 19751 3689 19763 3692
rect 19705 3683 19763 3689
rect 19978 3680 19984 3692
rect 20036 3720 20042 3732
rect 20622 3720 20628 3732
rect 20036 3692 20628 3720
rect 20036 3680 20042 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 21174 3720 21180 3732
rect 21135 3692 21180 3720
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 21266 3680 21272 3732
rect 21324 3720 21330 3732
rect 21453 3723 21511 3729
rect 21453 3720 21465 3723
rect 21324 3692 21465 3720
rect 21324 3680 21330 3692
rect 21453 3689 21465 3692
rect 21499 3720 21511 3723
rect 21542 3720 21548 3732
rect 21499 3692 21548 3720
rect 21499 3689 21511 3692
rect 21453 3683 21511 3689
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 24029 3723 24087 3729
rect 24029 3720 24041 3723
rect 21652 3692 24041 3720
rect 13446 3652 13452 3664
rect 12400 3624 12940 3652
rect 13407 3624 13452 3652
rect 12400 3612 12406 3624
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 15105 3655 15163 3661
rect 15105 3621 15117 3655
rect 15151 3652 15163 3655
rect 15378 3652 15384 3664
rect 15151 3624 15384 3652
rect 15151 3621 15163 3624
rect 15105 3615 15163 3621
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 15933 3655 15991 3661
rect 15933 3621 15945 3655
rect 15979 3652 15991 3655
rect 16298 3652 16304 3664
rect 15979 3624 16304 3652
rect 15979 3621 15991 3624
rect 15933 3615 15991 3621
rect 16298 3612 16304 3624
rect 16356 3612 16362 3664
rect 17405 3655 17463 3661
rect 17405 3621 17417 3655
rect 17451 3652 17463 3655
rect 17494 3652 17500 3664
rect 17451 3624 17500 3652
rect 17451 3621 17463 3624
rect 17405 3615 17463 3621
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 18874 3652 18880 3664
rect 18835 3624 18880 3652
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 21192 3652 21220 3680
rect 21652 3652 21680 3692
rect 24029 3689 24041 3692
rect 24075 3689 24087 3723
rect 24029 3683 24087 3689
rect 25501 3723 25559 3729
rect 25501 3689 25513 3723
rect 25547 3720 25559 3723
rect 25590 3720 25596 3732
rect 25547 3692 25596 3720
rect 25547 3689 25559 3692
rect 25501 3683 25559 3689
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 21192 3624 21680 3652
rect 22088 3655 22146 3661
rect 22088 3621 22100 3655
rect 22134 3652 22146 3655
rect 22186 3652 22192 3664
rect 22134 3624 22192 3652
rect 22134 3621 22146 3624
rect 22088 3615 22146 3621
rect 22186 3612 22192 3624
rect 22244 3652 22250 3664
rect 22646 3652 22652 3664
rect 22244 3624 22652 3652
rect 22244 3612 22250 3624
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 23474 3612 23480 3664
rect 23532 3652 23538 3664
rect 24489 3655 24547 3661
rect 24489 3652 24501 3655
rect 23532 3624 24501 3652
rect 23532 3612 23538 3624
rect 24489 3621 24501 3624
rect 24535 3652 24547 3655
rect 25682 3652 25688 3664
rect 24535 3624 25688 3652
rect 24535 3621 24547 3624
rect 24489 3615 24547 3621
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 9950 3593 9956 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 8812 3556 9689 3584
rect 8812 3544 8818 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9944 3547 9956 3593
rect 10008 3584 10014 3596
rect 10008 3556 10044 3584
rect 9950 3544 9956 3547
rect 10008 3544 10014 3556
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14001 3587 14059 3593
rect 14001 3584 14013 3587
rect 13872 3556 14013 3584
rect 13872 3544 13878 3556
rect 14001 3553 14013 3556
rect 14047 3553 14059 3587
rect 17770 3584 17776 3596
rect 14001 3547 14059 3553
rect 14108 3556 17776 3584
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8076 3488 8401 3516
rect 8076 3476 8082 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8536 3488 8581 3516
rect 8536 3476 8542 3488
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12710 3516 12716 3528
rect 11940 3488 12716 3516
rect 11940 3476 11946 3488
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 14108 3516 14136 3556
rect 13688 3488 14136 3516
rect 13688 3476 13694 3488
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 17512 3525 17540 3556
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 19659 3556 20392 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 17497 3519 17555 3525
rect 16080 3488 16125 3516
rect 16080 3476 16086 3488
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 18230 3516 18236 3528
rect 17727 3488 18236 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 19886 3516 19892 3528
rect 19847 3488 19892 3516
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 7834 3448 7840 3460
rect 7747 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3448 7898 3460
rect 8496 3448 8524 3476
rect 7892 3420 8524 3448
rect 12437 3451 12495 3457
rect 7892 3408 7898 3420
rect 12437 3417 12449 3451
rect 12483 3448 12495 3451
rect 12526 3448 12532 3460
rect 12483 3420 12532 3448
rect 12483 3417 12495 3420
rect 12437 3411 12495 3417
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 14737 3451 14795 3457
rect 14737 3417 14749 3451
rect 14783 3448 14795 3451
rect 15286 3448 15292 3460
rect 14783 3420 15292 3448
rect 14783 3417 14795 3420
rect 14737 3411 14795 3417
rect 15286 3408 15292 3420
rect 15344 3408 15350 3460
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 19245 3451 19303 3457
rect 19245 3448 19257 3451
rect 18196 3420 19257 3448
rect 18196 3408 18202 3420
rect 19245 3417 19257 3420
rect 19291 3417 19303 3451
rect 19245 3411 19303 3417
rect 5276 3352 7512 3380
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 8628 3352 9321 3380
rect 8628 3340 8634 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 12894 3380 12900 3392
rect 12391 3352 12900 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 12894 3340 12900 3352
rect 12952 3380 12958 3392
rect 13722 3380 13728 3392
rect 12952 3352 13728 3380
rect 12952 3340 12958 3352
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13906 3380 13912 3392
rect 13867 3352 13912 3380
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 14182 3380 14188 3392
rect 14143 3352 14188 3380
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 16577 3383 16635 3389
rect 16577 3349 16589 3383
rect 16623 3380 16635 3383
rect 16758 3380 16764 3392
rect 16623 3352 16764 3380
rect 16623 3349 16635 3352
rect 16577 3343 16635 3349
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 17034 3380 17040 3392
rect 16995 3352 17040 3380
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 20364 3389 20392 3556
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 21821 3587 21879 3593
rect 21821 3584 21833 3587
rect 21048 3556 21833 3584
rect 21048 3544 21054 3556
rect 21821 3553 21833 3556
rect 21867 3553 21879 3587
rect 21821 3547 21879 3553
rect 23658 3544 23664 3596
rect 23716 3584 23722 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 23716 3556 24409 3584
rect 23716 3544 23722 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24397 3547 24455 3553
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 23106 3408 23112 3460
rect 23164 3448 23170 3460
rect 23201 3451 23259 3457
rect 23201 3448 23213 3451
rect 23164 3420 23213 3448
rect 23164 3408 23170 3420
rect 23201 3417 23213 3420
rect 23247 3448 23259 3451
rect 25041 3451 25099 3457
rect 25041 3448 25053 3451
rect 23247 3420 25053 3448
rect 23247 3417 23259 3420
rect 23201 3411 23259 3417
rect 25041 3417 25053 3420
rect 25087 3417 25099 3451
rect 25041 3411 25099 3417
rect 20349 3383 20407 3389
rect 20349 3349 20361 3383
rect 20395 3380 20407 3383
rect 20530 3380 20536 3392
rect 20395 3352 20536 3380
rect 20395 3349 20407 3352
rect 20349 3343 20407 3349
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 20714 3380 20720 3392
rect 20627 3352 20720 3380
rect 20714 3340 20720 3352
rect 20772 3380 20778 3392
rect 22738 3380 22744 3392
rect 20772 3352 22744 3380
rect 20772 3340 20778 3352
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 23753 3383 23811 3389
rect 23753 3349 23765 3383
rect 23799 3380 23811 3383
rect 24118 3380 24124 3392
rect 23799 3352 24124 3380
rect 23799 3349 23811 3352
rect 23753 3343 23811 3349
rect 24118 3340 24124 3352
rect 24176 3380 24182 3392
rect 24762 3380 24768 3392
rect 24176 3352 24768 3380
rect 24176 3340 24182 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 5258 3176 5264 3188
rect 3108 3148 3153 3176
rect 5219 3148 5264 3176
rect 3108 3136 3114 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 5994 3176 6000 3188
rect 5859 3148 6000 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6178 3176 6184 3188
rect 6139 3148 6184 3176
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 10008 3148 10149 3176
rect 10008 3136 10014 3148
rect 10137 3145 10149 3148
rect 10183 3176 10195 3179
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10183 3148 10425 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10413 3145 10425 3148
rect 10459 3176 10471 3179
rect 10778 3176 10784 3188
rect 10459 3148 10784 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11238 3176 11244 3188
rect 11011 3148 11244 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 3418 3108 3424 3120
rect 3379 3080 3424 3108
rect 3418 3068 3424 3080
rect 3476 3068 3482 3120
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2409 2975 2467 2981
rect 2409 2972 2421 2975
rect 2372 2944 2421 2972
rect 2372 2932 2378 2944
rect 2409 2941 2421 2944
rect 2455 2941 2467 2975
rect 2608 2972 2636 3003
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3384 3012 3617 3040
rect 3384 3000 3390 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 6196 3040 6224 3136
rect 6365 3111 6423 3117
rect 6365 3077 6377 3111
rect 6411 3108 6423 3111
rect 6641 3111 6699 3117
rect 6641 3108 6653 3111
rect 6411 3080 6653 3108
rect 6411 3077 6423 3080
rect 6365 3071 6423 3077
rect 6641 3077 6653 3080
rect 6687 3108 6699 3111
rect 8018 3108 8024 3120
rect 6687 3080 7420 3108
rect 7979 3080 8024 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7392 3049 7420 3080
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 6196 3012 7297 3040
rect 3605 3003 3663 3009
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 7377 3003 7435 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 3050 2972 3056 2984
rect 2608 2944 3056 2972
rect 2409 2935 2467 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 11072 2981 11100 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 11940 3148 11985 3176
rect 11940 3136 11946 3148
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13136 3148 13829 3176
rect 13136 3136 13142 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 15749 3179 15807 3185
rect 15749 3145 15761 3179
rect 15795 3176 15807 3179
rect 15838 3176 15844 3188
rect 15795 3148 15844 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 16850 3176 16856 3188
rect 16163 3148 16856 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16209 3111 16267 3117
rect 16209 3108 16221 3111
rect 15304 3080 16221 3108
rect 11330 3040 11336 3052
rect 11291 3012 11336 3040
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 13872 3012 14105 3040
rect 13872 3000 13878 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 14093 3003 14151 3009
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14516 3012 14565 3040
rect 14516 3000 14522 3012
rect 14553 3009 14565 3012
rect 14599 3040 14611 3043
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14599 3012 15209 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 7156 2944 7205 2972
rect 7156 2932 7162 2944
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12710 2981 12716 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12308 2944 12449 2972
rect 12308 2932 12314 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12704 2972 12716 2981
rect 12671 2944 12716 2972
rect 12437 2935 12495 2941
rect 12704 2935 12716 2944
rect 12710 2932 12716 2935
rect 12768 2932 12774 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14792 2944 15025 2972
rect 14792 2932 14798 2944
rect 15013 2941 15025 2944
rect 15059 2972 15071 2975
rect 15304 2972 15332 3080
rect 16209 3077 16221 3080
rect 16255 3077 16267 3111
rect 16209 3071 16267 3077
rect 16684 3049 16712 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 17770 3176 17776 3188
rect 17359 3148 17776 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 18288 3148 18337 3176
rect 18288 3136 18294 3148
rect 18325 3145 18337 3148
rect 18371 3176 18383 3179
rect 18598 3176 18604 3188
rect 18371 3148 18604 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 20165 3179 20223 3185
rect 20165 3176 20177 3179
rect 19944 3148 20177 3176
rect 19944 3136 19950 3148
rect 20165 3145 20177 3148
rect 20211 3176 20223 3179
rect 22002 3176 22008 3188
rect 20211 3148 22008 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22281 3179 22339 3185
rect 22281 3176 22293 3179
rect 22244 3148 22293 3176
rect 22244 3136 22250 3148
rect 22281 3145 22293 3148
rect 22327 3145 22339 3179
rect 22738 3176 22744 3188
rect 22699 3148 22744 3176
rect 22281 3139 22339 3145
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23658 3176 23664 3188
rect 23155 3148 23664 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 24946 3176 24952 3188
rect 24728 3148 24952 3176
rect 24728 3136 24734 3148
rect 24946 3136 24952 3148
rect 25004 3176 25010 3188
rect 25041 3179 25099 3185
rect 25041 3176 25053 3179
rect 25004 3148 25053 3176
rect 25004 3136 25010 3148
rect 25041 3145 25053 3148
rect 25087 3176 25099 3179
rect 25317 3179 25375 3185
rect 25317 3176 25329 3179
rect 25087 3148 25329 3176
rect 25087 3145 25099 3148
rect 25041 3139 25099 3145
rect 25317 3145 25329 3148
rect 25363 3145 25375 3179
rect 25682 3176 25688 3188
rect 25643 3148 25688 3176
rect 25317 3139 25375 3145
rect 25682 3136 25688 3148
rect 25740 3136 25746 3188
rect 19797 3111 19855 3117
rect 19797 3077 19809 3111
rect 19843 3108 19855 3111
rect 20438 3108 20444 3120
rect 19843 3080 20444 3108
rect 19843 3077 19855 3080
rect 19797 3071 19855 3077
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 25590 3068 25596 3120
rect 25648 3108 25654 3120
rect 26050 3108 26056 3120
rect 25648 3080 26056 3108
rect 25648 3068 25654 3080
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16816 3012 16865 3040
rect 16816 3000 16822 3012
rect 16853 3009 16865 3012
rect 16899 3040 16911 3043
rect 18230 3040 18236 3052
rect 16899 3012 18236 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 20456 3040 20484 3068
rect 20456 3012 20760 3040
rect 15059 2944 15332 2972
rect 18417 2975 18475 2981
rect 15059 2941 15071 2944
rect 15013 2935 15071 2941
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 19058 2972 19064 2984
rect 18463 2944 19064 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 20625 2975 20683 2981
rect 20625 2941 20637 2975
rect 20671 2941 20683 2975
rect 20732 2972 20760 3012
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 23164 3012 23397 3040
rect 23164 3000 23170 3012
rect 23385 3009 23397 3012
rect 23431 3040 23443 3043
rect 23431 3012 23796 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 20898 2981 20904 2984
rect 20881 2975 20904 2981
rect 20881 2972 20893 2975
rect 20732 2944 20893 2972
rect 20625 2935 20683 2941
rect 20881 2941 20893 2944
rect 20956 2972 20962 2984
rect 23661 2975 23719 2981
rect 20956 2944 21029 2972
rect 20881 2935 20904 2941
rect 3872 2907 3930 2913
rect 3872 2873 3884 2907
rect 3918 2904 3930 2907
rect 3970 2904 3976 2916
rect 3918 2876 3976 2904
rect 3918 2873 3930 2876
rect 3872 2867 3930 2873
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 9002 2907 9060 2913
rect 9002 2904 9014 2907
rect 8904 2876 9014 2904
rect 8904 2864 8910 2876
rect 9002 2873 9014 2876
rect 9048 2873 9060 2907
rect 9002 2867 9060 2873
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 15102 2904 15108 2916
rect 13964 2876 15108 2904
rect 13964 2864 13970 2876
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 16574 2904 16580 2916
rect 16535 2876 16580 2904
rect 16574 2864 16580 2876
rect 16632 2864 16638 2916
rect 18684 2907 18742 2913
rect 18684 2873 18696 2907
rect 18730 2904 18742 2907
rect 18874 2904 18880 2916
rect 18730 2876 18880 2904
rect 18730 2873 18742 2876
rect 18684 2867 18742 2873
rect 18874 2864 18880 2876
rect 18932 2864 18938 2916
rect 20640 2904 20668 2935
rect 20898 2932 20904 2935
rect 20956 2932 20962 2944
rect 23661 2941 23673 2975
rect 23707 2941 23719 2975
rect 23768 2972 23796 3012
rect 23917 2975 23975 2981
rect 23917 2972 23929 2975
rect 23768 2944 23929 2972
rect 23661 2935 23719 2941
rect 23917 2941 23929 2944
rect 23963 2941 23975 2975
rect 23917 2935 23975 2941
rect 20990 2904 20996 2916
rect 20640 2876 20996 2904
rect 20990 2864 20996 2876
rect 21048 2864 21054 2916
rect 23676 2904 23704 2935
rect 25590 2904 25596 2916
rect 23676 2876 25596 2904
rect 25590 2864 25596 2876
rect 25648 2864 25654 2916
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 2556 2808 2601 2836
rect 2556 2796 2562 2808
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4985 2839 5043 2845
rect 4985 2836 4997 2839
rect 3568 2808 4997 2836
rect 3568 2796 3574 2808
rect 4985 2805 4997 2808
rect 5031 2836 5043 2839
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 5031 2808 6377 2836
rect 5031 2805 5043 2808
rect 4985 2799 5043 2805
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6365 2799 6423 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12986 2836 12992 2848
rect 12299 2808 12992 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 14642 2836 14648 2848
rect 14603 2808 14648 2836
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17552 2808 17601 2836
rect 17552 2796 17558 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 17589 2799 17647 2805
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 25222 2836 25228 2848
rect 20404 2808 25228 2836
rect 20404 2796 20410 2808
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1394 2632 1400 2644
rect 1355 2604 1400 2632
rect 1394 2592 1400 2604
rect 1452 2592 1458 2644
rect 1854 2632 1860 2644
rect 1815 2604 1860 2632
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2372 2604 2421 2632
rect 2372 2592 2378 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3786 2632 3792 2644
rect 2823 2604 3792 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5350 2632 5356 2644
rect 5215 2604 5356 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 3418 2564 3424 2576
rect 3379 2536 3424 2564
rect 3418 2524 3424 2536
rect 3476 2564 3482 2576
rect 4433 2567 4491 2573
rect 4433 2564 4445 2567
rect 3476 2536 4445 2564
rect 3476 2524 3482 2536
rect 4433 2533 4445 2536
rect 4479 2564 4491 2567
rect 4522 2564 4528 2576
rect 4479 2536 4528 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 2915 2468 4108 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 4080 2369 4108 2468
rect 4522 2428 4528 2440
rect 4483 2400 4528 2428
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5184 2428 5212 2595
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6454 2632 6460 2644
rect 6411 2604 6460 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6380 2496 6408 2595
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 7340 2604 7757 2632
rect 7340 2592 7346 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 7745 2595 7803 2601
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9769 2635 9827 2641
rect 9769 2632 9781 2635
rect 9732 2604 9781 2632
rect 9732 2592 9738 2604
rect 9769 2601 9781 2604
rect 9815 2601 9827 2635
rect 9769 2595 9827 2601
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 11238 2632 11244 2644
rect 10183 2604 11244 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12342 2632 12348 2644
rect 12115 2604 12348 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 15930 2632 15936 2644
rect 14599 2604 15936 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 17773 2635 17831 2641
rect 16632 2604 16677 2632
rect 16632 2592 16638 2604
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 17954 2632 17960 2644
rect 17819 2604 17960 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 17954 2592 17960 2604
rect 18012 2632 18018 2644
rect 18138 2632 18144 2644
rect 18012 2604 18144 2632
rect 18012 2592 18018 2604
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2601 18383 2635
rect 18325 2595 18383 2601
rect 19797 2635 19855 2641
rect 19797 2601 19809 2635
rect 19843 2632 19855 2635
rect 19978 2632 19984 2644
rect 19843 2604 19984 2632
rect 19843 2601 19855 2604
rect 19797 2595 19855 2601
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 12437 2567 12495 2573
rect 9631 2536 10456 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 5767 2468 6408 2496
rect 7653 2499 7711 2505
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8018 2496 8024 2508
rect 7699 2468 8024 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8018 2456 8024 2468
rect 8076 2496 8082 2508
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 8076 2468 8125 2496
rect 8076 2456 8082 2468
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8260 2468 8305 2496
rect 8260 2456 8266 2468
rect 4755 2400 5212 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 6972 2400 7297 2428
rect 6972 2388 6978 2400
rect 7285 2397 7297 2400
rect 7331 2428 7343 2431
rect 8220 2428 8248 2456
rect 7331 2400 8248 2428
rect 8389 2431 8447 2437
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8478 2428 8484 2440
rect 8435 2400 8484 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8478 2388 8484 2400
rect 8536 2428 8542 2440
rect 10428 2437 10456 2536
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12888 2567 12946 2573
rect 12888 2564 12900 2567
rect 12483 2536 12900 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 12888 2533 12900 2536
rect 12934 2564 12946 2567
rect 12986 2564 12992 2576
rect 12934 2536 12992 2564
rect 12934 2533 12946 2536
rect 12888 2527 12946 2533
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 14516 2536 14841 2564
rect 14516 2524 14522 2536
rect 14829 2533 14841 2536
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11514 2496 11520 2508
rect 11471 2468 11520 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8536 2400 9137 2428
rect 8536 2388 8542 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10686 2428 10692 2440
rect 10459 2400 10692 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 4065 2363 4123 2369
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 5537 2363 5595 2369
rect 5537 2360 5549 2363
rect 4111 2332 5549 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 5537 2329 5549 2332
rect 5583 2329 5595 2363
rect 10244 2360 10272 2391
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12618 2428 12624 2440
rect 12308 2400 12624 2428
rect 12308 2388 12314 2400
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 14844 2428 14872 2527
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15841 2567 15899 2573
rect 15841 2564 15853 2567
rect 15344 2536 15853 2564
rect 15344 2524 15350 2536
rect 15841 2533 15853 2536
rect 15887 2564 15899 2567
rect 18340 2564 18368 2595
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20530 2592 20536 2644
rect 20588 2632 20594 2644
rect 21177 2635 21235 2641
rect 21177 2632 21189 2635
rect 20588 2604 21189 2632
rect 20588 2592 20594 2604
rect 21177 2601 21189 2604
rect 21223 2601 21235 2635
rect 21177 2595 21235 2601
rect 21545 2635 21603 2641
rect 21545 2601 21557 2635
rect 21591 2632 21603 2635
rect 22281 2635 22339 2641
rect 22281 2632 22293 2635
rect 21591 2604 22293 2632
rect 21591 2601 21603 2604
rect 21545 2595 21603 2601
rect 22281 2601 22293 2604
rect 22327 2632 22339 2635
rect 22462 2632 22468 2644
rect 22327 2604 22468 2632
rect 22327 2601 22339 2604
rect 22281 2595 22339 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 24026 2632 24032 2644
rect 23987 2604 24032 2632
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 24946 2592 24952 2644
rect 25004 2632 25010 2644
rect 25041 2635 25099 2641
rect 25041 2632 25053 2635
rect 25004 2604 25053 2632
rect 25004 2592 25010 2604
rect 25041 2601 25053 2604
rect 25087 2601 25099 2635
rect 25590 2632 25596 2644
rect 25551 2604 25596 2632
rect 25041 2595 25099 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 20898 2564 20904 2576
rect 15887 2536 18368 2564
rect 20859 2536 20904 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 25501 2567 25559 2573
rect 25501 2533 25513 2567
rect 25547 2564 25559 2567
rect 26050 2564 26056 2576
rect 25547 2536 26056 2564
rect 25547 2533 25559 2536
rect 25501 2527 25559 2533
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 15197 2499 15255 2505
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 16298 2496 16304 2508
rect 15243 2468 16304 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 16298 2456 16304 2468
rect 16356 2456 16362 2508
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16908 2468 17049 2496
rect 16908 2456 16914 2468
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 18046 2496 18052 2508
rect 18007 2468 18052 2496
rect 17037 2459 17095 2465
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 18138 2456 18144 2508
rect 18196 2496 18202 2508
rect 18693 2499 18751 2505
rect 18693 2496 18705 2499
rect 18196 2468 18705 2496
rect 18196 2456 18202 2468
rect 18693 2465 18705 2468
rect 18739 2465 18751 2499
rect 20530 2496 20536 2508
rect 20491 2468 20536 2496
rect 18693 2459 18751 2465
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20916 2496 20944 2524
rect 20916 2468 21772 2496
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 14844 2400 16037 2428
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 18064 2428 18092 2456
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18064 2400 18797 2428
rect 16025 2391 16083 2397
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18923 2400 19349 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 20548 2428 20576 2456
rect 21744 2437 21772 2468
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 23808 2468 24409 2496
rect 23808 2456 23814 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 20548 2400 21649 2428
rect 19337 2391 19395 2397
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 21729 2431 21787 2437
rect 21729 2397 21741 2431
rect 21775 2397 21787 2431
rect 21729 2391 21787 2397
rect 24489 2431 24547 2437
rect 24489 2397 24501 2431
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 24946 2428 24952 2440
rect 24719 2400 24952 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 10870 2360 10876 2372
rect 10244 2332 10876 2360
rect 5537 2323 5595 2329
rect 10870 2320 10876 2332
rect 10928 2320 10934 2372
rect 15470 2360 15476 2372
rect 15431 2332 15476 2360
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 16724 2332 17233 2360
rect 16724 2320 16730 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18892 2360 18920 2391
rect 23474 2360 23480 2372
rect 18288 2332 18920 2360
rect 23435 2332 23480 2360
rect 18288 2320 18294 2332
rect 23474 2320 23480 2332
rect 23532 2360 23538 2372
rect 24504 2360 24532 2391
rect 24946 2388 24952 2400
rect 25004 2388 25010 2440
rect 23532 2332 24532 2360
rect 23532 2320 23538 2332
rect 3786 2292 3792 2304
rect 3747 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2292 3850 2304
rect 4522 2292 4528 2304
rect 3844 2264 4528 2292
rect 3844 2252 3850 2264
rect 4522 2252 4528 2264
rect 4580 2292 4586 2304
rect 4706 2292 4712 2304
rect 4580 2264 4712 2292
rect 4580 2252 4586 2264
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 6178 2292 6184 2304
rect 5951 2264 6184 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 8846 2292 8852 2304
rect 8807 2264 8852 2292
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13998 2292 14004 2304
rect 13959 2264 14004 2292
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 16850 2292 16856 2304
rect 16811 2264 16856 2292
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 20162 2292 20168 2304
rect 20123 2264 20168 2292
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 22554 2292 22560 2304
rect 22515 2264 22560 2292
rect 22554 2252 22560 2264
rect 22612 2252 22618 2304
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 23750 2292 23756 2304
rect 23711 2264 23756 2292
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 12618 2048 12624 2100
rect 12676 2088 12682 2100
rect 17678 2088 17684 2100
rect 12676 2060 17684 2088
rect 12676 2048 12682 2060
rect 17678 2048 17684 2060
rect 17736 2048 17742 2100
rect 3050 1368 3056 1420
rect 3108 1408 3114 1420
rect 8386 1408 8392 1420
rect 3108 1380 8392 1408
rect 3108 1368 3114 1380
rect 8386 1368 8392 1380
rect 8444 1368 8450 1420
rect 4890 552 4896 604
rect 4948 592 4954 604
rect 5258 592 5264 604
rect 4948 564 5264 592
rect 4948 552 4954 564
rect 5258 552 5264 564
rect 5316 552 5322 604
rect 12158 552 12164 604
rect 12216 592 12222 604
rect 12526 592 12532 604
rect 12216 564 12532 592
rect 12216 552 12222 564
rect 12526 552 12532 564
rect 12584 552 12590 604
<< via1 >>
rect 3700 25984 3752 26036
rect 8300 25984 8352 26036
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 24124 25168 24176 25220
rect 24492 25168 24544 25220
rect 4068 25100 4120 25152
rect 5540 25100 5592 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 5540 23808 5592 23860
rect 24216 23808 24268 23860
rect 24124 23604 24176 23656
rect 6828 23468 6880 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24860 23264 24912 23316
rect 24676 23128 24728 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 24860 22720 24912 22772
rect 24952 22559 25004 22568
rect 24952 22525 24961 22559
rect 24961 22525 24995 22559
rect 24995 22525 25004 22559
rect 24952 22516 25004 22525
rect 2044 22423 2096 22432
rect 2044 22389 2053 22423
rect 2053 22389 2087 22423
rect 2087 22389 2096 22423
rect 2044 22380 2096 22389
rect 23480 22423 23532 22432
rect 23480 22389 23489 22423
rect 23489 22389 23523 22423
rect 23523 22389 23532 22423
rect 23480 22380 23532 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 2044 21335 2096 21344
rect 2044 21301 2053 21335
rect 2053 21301 2087 21335
rect 2087 21301 2096 21335
rect 2044 21292 2096 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 2044 21063 2096 21072
rect 2044 21029 2053 21063
rect 2053 21029 2087 21063
rect 2087 21029 2096 21063
rect 2044 21020 2096 21029
rect 2320 20952 2372 21004
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1492 20544 1544 20596
rect 21548 20587 21600 20596
rect 21548 20553 21557 20587
rect 21557 20553 21591 20587
rect 21591 20553 21600 20587
rect 21548 20544 21600 20553
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 19340 20204 19392 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 2412 19864 2464 19916
rect 24216 19864 24268 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19252 1636 19304
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 1492 19116 1544 19168
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 24676 19116 24728 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2688 18955 2740 18964
rect 2688 18921 2697 18955
rect 2697 18921 2731 18955
rect 2731 18921 2740 18955
rect 2688 18912 2740 18921
rect 18236 18955 18288 18964
rect 18236 18921 18245 18955
rect 18245 18921 18279 18955
rect 18279 18921 18288 18955
rect 18236 18912 18288 18921
rect 4344 18887 4396 18896
rect 4344 18853 4353 18887
rect 4353 18853 4387 18887
rect 4387 18853 4396 18887
rect 4344 18844 4396 18853
rect 23940 18844 23992 18896
rect 25320 18844 25372 18896
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 1768 18572 1820 18624
rect 3148 18776 3200 18828
rect 4436 18776 4488 18828
rect 17960 18776 18012 18828
rect 23480 18819 23532 18828
rect 23480 18785 23489 18819
rect 23489 18785 23523 18819
rect 23523 18785 23532 18819
rect 23480 18776 23532 18785
rect 24216 18776 24268 18828
rect 23296 18708 23348 18760
rect 2964 18572 3016 18624
rect 24032 18572 24084 18624
rect 24768 18615 24820 18624
rect 24768 18581 24777 18615
rect 24777 18581 24811 18615
rect 24811 18581 24820 18615
rect 24768 18572 24820 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1400 18368 1452 18420
rect 24124 18368 24176 18420
rect 24584 18207 24636 18216
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 2320 18028 2372 18037
rect 2780 18028 2832 18080
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 3884 18028 3936 18080
rect 4436 18028 4488 18080
rect 17960 18028 18012 18080
rect 23020 18028 23072 18080
rect 24584 18173 24593 18207
rect 24593 18173 24627 18207
rect 24627 18173 24636 18207
rect 24584 18164 24636 18173
rect 23204 18028 23256 18080
rect 23480 18028 23532 18080
rect 24216 18028 24268 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 4160 17824 4212 17876
rect 24676 17824 24728 17876
rect 2320 17756 2372 17808
rect 17868 17756 17920 17808
rect 1492 17688 1544 17740
rect 1768 17688 1820 17740
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 4344 17688 4396 17740
rect 16856 17688 16908 17740
rect 21824 17688 21876 17740
rect 22468 17688 22520 17740
rect 23572 17688 23624 17740
rect 24676 17688 24728 17740
rect 2136 17620 2188 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 2044 17484 2096 17536
rect 2228 17484 2280 17536
rect 3424 17484 3476 17536
rect 3608 17527 3660 17536
rect 3608 17493 3617 17527
rect 3617 17493 3651 17527
rect 3651 17493 3660 17527
rect 3608 17484 3660 17493
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 23480 17484 23532 17536
rect 23664 17527 23716 17536
rect 23664 17493 23673 17527
rect 23673 17493 23707 17527
rect 23707 17493 23716 17527
rect 23664 17484 23716 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 23756 17280 23808 17332
rect 23848 17212 23900 17264
rect 24676 17212 24728 17264
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 2964 17144 3016 17196
rect 13360 17144 13412 17196
rect 3148 17119 3200 17128
rect 3148 17085 3157 17119
rect 3157 17085 3191 17119
rect 3191 17085 3200 17119
rect 3148 17076 3200 17085
rect 3608 17076 3660 17128
rect 4804 17076 4856 17128
rect 13084 17076 13136 17128
rect 2780 17051 2832 17060
rect 2780 17017 2789 17051
rect 2789 17017 2823 17051
rect 2823 17017 2832 17051
rect 2780 17008 2832 17017
rect 13268 17008 13320 17060
rect 18420 17008 18472 17060
rect 22008 17144 22060 17196
rect 20720 17076 20772 17128
rect 24492 17076 24544 17128
rect 22284 17008 22336 17060
rect 22468 17051 22520 17060
rect 22468 17017 22477 17051
rect 22477 17017 22511 17051
rect 22511 17017 22520 17051
rect 22468 17008 22520 17017
rect 23572 17008 23624 17060
rect 24768 17008 24820 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1676 16940 1728 16992
rect 4344 16940 4396 16992
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12900 16940 12952 16992
rect 16856 16940 16908 16992
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 20720 16940 20772 16992
rect 20996 16983 21048 16992
rect 20996 16949 21005 16983
rect 21005 16949 21039 16983
rect 21039 16949 21048 16983
rect 20996 16940 21048 16949
rect 21824 16940 21876 16992
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16736 1636 16788
rect 4068 16736 4120 16788
rect 12256 16736 12308 16788
rect 18420 16736 18472 16788
rect 19984 16736 20036 16788
rect 21916 16736 21968 16788
rect 23940 16736 23992 16788
rect 25504 16779 25556 16788
rect 25504 16745 25513 16779
rect 25513 16745 25547 16779
rect 25547 16745 25556 16779
rect 25504 16736 25556 16745
rect 1676 16600 1728 16652
rect 2504 16600 2556 16652
rect 2780 16600 2832 16652
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 4252 16600 4304 16652
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 5448 16600 5500 16652
rect 13452 16600 13504 16652
rect 14188 16600 14240 16652
rect 17408 16668 17460 16720
rect 21456 16668 21508 16720
rect 22836 16711 22888 16720
rect 22836 16677 22845 16711
rect 22845 16677 22879 16711
rect 22879 16677 22888 16711
rect 22836 16668 22888 16677
rect 24216 16668 24268 16720
rect 17040 16600 17092 16652
rect 4160 16532 4212 16584
rect 2872 16507 2924 16516
rect 2872 16473 2881 16507
rect 2881 16473 2915 16507
rect 2915 16473 2924 16507
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 18604 16532 18656 16584
rect 19708 16643 19760 16652
rect 19708 16609 19717 16643
rect 19717 16609 19751 16643
rect 19751 16609 19760 16643
rect 19708 16600 19760 16609
rect 20076 16532 20128 16584
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 24676 16600 24728 16652
rect 25780 16600 25832 16652
rect 2872 16464 2924 16473
rect 21272 16464 21324 16516
rect 22008 16532 22060 16584
rect 22744 16532 22796 16584
rect 2136 16396 2188 16448
rect 5540 16396 5592 16448
rect 10784 16396 10836 16448
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 20444 16396 20496 16448
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 22468 16439 22520 16448
rect 22468 16405 22477 16439
rect 22477 16405 22511 16439
rect 22511 16405 22520 16439
rect 22468 16396 22520 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1400 16192 1452 16244
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 5540 16192 5592 16244
rect 6368 16192 6420 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 20076 16235 20128 16244
rect 20076 16201 20085 16235
rect 20085 16201 20119 16235
rect 20119 16201 20128 16235
rect 20076 16192 20128 16201
rect 22928 16192 22980 16244
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 3240 16124 3292 16176
rect 22008 16124 22060 16176
rect 1584 16056 1636 16108
rect 2504 16056 2556 16108
rect 2872 16056 2924 16108
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 12532 16056 12584 16108
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 20352 16056 20404 16108
rect 21364 16056 21416 16108
rect 22744 16124 22796 16176
rect 23940 16056 23992 16108
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 2964 15988 3016 16040
rect 4160 16031 4212 16040
rect 4160 15997 4169 16031
rect 4169 15997 4203 16031
rect 4203 15997 4212 16031
rect 4160 15988 4212 15997
rect 12072 15988 12124 16040
rect 1768 15852 1820 15904
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 3332 15852 3384 15904
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 11704 15852 11756 15904
rect 12164 15920 12216 15972
rect 13360 15920 13412 15972
rect 20444 16031 20496 16040
rect 20444 15997 20453 16031
rect 20453 15997 20487 16031
rect 20487 15997 20496 16031
rect 20444 15988 20496 15997
rect 22008 16031 22060 16040
rect 22008 15997 22017 16031
rect 22017 15997 22051 16031
rect 22051 15997 22060 16031
rect 22008 15988 22060 15997
rect 22836 15988 22888 16040
rect 14096 15920 14148 15972
rect 14832 15920 14884 15972
rect 17960 15920 18012 15972
rect 19708 15963 19760 15972
rect 19708 15929 19717 15963
rect 19717 15929 19751 15963
rect 19751 15929 19760 15963
rect 19708 15920 19760 15929
rect 21732 15920 21784 15972
rect 23480 15963 23532 15972
rect 23480 15929 23489 15963
rect 23489 15929 23523 15963
rect 23523 15929 23532 15963
rect 23480 15920 23532 15929
rect 24124 15920 24176 15972
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 12808 15852 12860 15904
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 13452 15852 13504 15861
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 14280 15852 14332 15904
rect 15936 15852 15988 15904
rect 16304 15852 16356 15904
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 18052 15895 18104 15904
rect 18052 15861 18061 15895
rect 18061 15861 18095 15895
rect 18095 15861 18104 15895
rect 18052 15852 18104 15861
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 18696 15852 18748 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 21640 15895 21692 15904
rect 21640 15861 21649 15895
rect 21649 15861 21683 15895
rect 21683 15861 21692 15895
rect 21640 15852 21692 15861
rect 23572 15852 23624 15904
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 3056 15648 3108 15700
rect 3884 15648 3936 15700
rect 5172 15648 5224 15700
rect 6368 15691 6420 15700
rect 6368 15657 6377 15691
rect 6377 15657 6411 15691
rect 6411 15657 6420 15691
rect 6368 15648 6420 15657
rect 6828 15648 6880 15700
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 13360 15648 13412 15700
rect 14556 15648 14608 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 20444 15648 20496 15700
rect 22468 15648 22520 15700
rect 2320 15580 2372 15632
rect 5448 15580 5500 15632
rect 2136 15555 2188 15564
rect 2136 15521 2145 15555
rect 2145 15521 2179 15555
rect 2179 15521 2188 15555
rect 2136 15512 2188 15521
rect 3148 15512 3200 15564
rect 3700 15512 3752 15564
rect 6000 15512 6052 15564
rect 7656 15512 7708 15564
rect 11796 15555 11848 15564
rect 11796 15521 11830 15555
rect 11830 15521 11848 15555
rect 11796 15512 11848 15521
rect 12440 15580 12492 15632
rect 17960 15580 18012 15632
rect 13636 15512 13688 15564
rect 1952 15444 2004 15496
rect 2504 15444 2556 15496
rect 4252 15444 4304 15496
rect 4804 15444 4856 15496
rect 10048 15444 10100 15496
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 1768 15376 1820 15428
rect 5540 15419 5592 15428
rect 5540 15385 5549 15419
rect 5549 15385 5583 15419
rect 5583 15385 5592 15419
rect 5540 15376 5592 15385
rect 12808 15376 12860 15428
rect 13728 15376 13780 15428
rect 17500 15444 17552 15496
rect 18236 15444 18288 15496
rect 19616 15555 19668 15564
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 19524 15444 19576 15496
rect 22192 15580 22244 15632
rect 22560 15580 22612 15632
rect 22744 15623 22796 15632
rect 22744 15589 22753 15623
rect 22753 15589 22787 15623
rect 22787 15589 22796 15623
rect 22744 15580 22796 15589
rect 24676 15623 24728 15632
rect 24676 15589 24685 15623
rect 24685 15589 24719 15623
rect 24719 15589 24728 15623
rect 24676 15580 24728 15589
rect 24952 15580 25004 15632
rect 23664 15512 23716 15564
rect 25044 15512 25096 15564
rect 20444 15444 20496 15496
rect 22100 15444 22152 15496
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 23572 15444 23624 15496
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 20536 15376 20588 15428
rect 1308 15308 1360 15360
rect 2320 15308 2372 15360
rect 2504 15308 2556 15360
rect 2780 15308 2832 15360
rect 2964 15308 3016 15360
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 4988 15308 5040 15360
rect 8116 15308 8168 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 13176 15308 13228 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15292 15351 15344 15360
rect 15292 15317 15301 15351
rect 15301 15317 15335 15351
rect 15335 15317 15344 15351
rect 15292 15308 15344 15317
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 16580 15308 16632 15360
rect 17408 15308 17460 15360
rect 18880 15308 18932 15360
rect 20444 15308 20496 15360
rect 21272 15308 21324 15360
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 21732 15351 21784 15360
rect 21732 15317 21741 15351
rect 21741 15317 21775 15351
rect 21775 15317 21784 15351
rect 21732 15308 21784 15317
rect 22468 15308 22520 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 6828 15104 6880 15156
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 10140 15104 10192 15156
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 13820 15104 13872 15156
rect 17868 15104 17920 15156
rect 21364 15104 21416 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 22376 15104 22428 15156
rect 12440 15036 12492 15088
rect 13636 15036 13688 15088
rect 14188 15079 14240 15088
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 19340 15036 19392 15088
rect 24768 15036 24820 15088
rect 3608 15011 3660 15020
rect 3608 14977 3617 15011
rect 3617 14977 3651 15011
rect 3651 14977 3660 15011
rect 3608 14968 3660 14977
rect 4804 14968 4856 15020
rect 6920 14968 6972 15020
rect 11060 14968 11112 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 4068 14900 4120 14952
rect 4344 14900 4396 14952
rect 4988 14943 5040 14952
rect 4988 14909 4997 14943
rect 4997 14909 5031 14943
rect 5031 14909 5040 14943
rect 4988 14900 5040 14909
rect 6000 14900 6052 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8024 14900 8076 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 14740 14968 14792 15020
rect 16764 15011 16816 15020
rect 16764 14977 16773 15011
rect 16773 14977 16807 15011
rect 16807 14977 16816 15011
rect 16764 14968 16816 14977
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 23388 14968 23440 15020
rect 23848 14968 23900 15020
rect 13176 14900 13228 14952
rect 15844 14900 15896 14952
rect 16948 14900 17000 14952
rect 18788 14900 18840 14952
rect 2136 14764 2188 14816
rect 2412 14807 2464 14816
rect 2412 14773 2421 14807
rect 2421 14773 2455 14807
rect 2455 14773 2464 14807
rect 2412 14764 2464 14773
rect 2872 14764 2924 14816
rect 3884 14764 3936 14816
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 4804 14764 4856 14816
rect 12808 14832 12860 14884
rect 14648 14832 14700 14884
rect 18604 14832 18656 14884
rect 20536 14900 20588 14952
rect 21916 14900 21968 14952
rect 22284 14943 22336 14952
rect 22284 14909 22293 14943
rect 22293 14909 22327 14943
rect 22327 14909 22336 14943
rect 22284 14900 22336 14909
rect 23664 14900 23716 14952
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 19616 14832 19668 14884
rect 20076 14832 20128 14884
rect 21548 14832 21600 14884
rect 22100 14832 22152 14884
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 12992 14764 13044 14816
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 18328 14764 18380 14816
rect 18972 14764 19024 14816
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20444 14764 20496 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2688 14560 2740 14612
rect 3424 14560 3476 14612
rect 4528 14560 4580 14612
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 7932 14560 7984 14612
rect 11796 14560 11848 14612
rect 14740 14603 14792 14612
rect 14740 14569 14749 14603
rect 14749 14569 14783 14603
rect 14783 14569 14792 14603
rect 14740 14560 14792 14569
rect 18236 14560 18288 14612
rect 20536 14560 20588 14612
rect 20720 14560 20772 14612
rect 22284 14560 22336 14612
rect 23572 14560 23624 14612
rect 2688 14424 2740 14476
rect 4620 14424 4672 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 4528 14356 4580 14408
rect 6644 14492 6696 14544
rect 12992 14492 13044 14544
rect 5448 14424 5500 14476
rect 6184 14424 6236 14476
rect 8208 14424 8260 14476
rect 10876 14424 10928 14476
rect 6092 14356 6144 14408
rect 13636 14424 13688 14476
rect 14004 14424 14056 14476
rect 16028 14424 16080 14476
rect 4160 14288 4212 14340
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 3608 14220 3660 14272
rect 3700 14220 3752 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 6460 14220 6512 14272
rect 7840 14220 7892 14272
rect 8116 14220 8168 14272
rect 9128 14220 9180 14272
rect 14740 14356 14792 14408
rect 16120 14356 16172 14408
rect 10968 14220 11020 14272
rect 11520 14220 11572 14272
rect 12440 14288 12492 14340
rect 15016 14331 15068 14340
rect 15016 14297 15025 14331
rect 15025 14297 15059 14331
rect 15059 14297 15068 14331
rect 15016 14288 15068 14297
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 15660 14220 15712 14272
rect 15936 14220 15988 14272
rect 16396 14220 16448 14272
rect 16764 14492 16816 14544
rect 17224 14467 17276 14476
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17224 14424 17276 14433
rect 16948 14356 17000 14408
rect 21364 14492 21416 14544
rect 22100 14492 22152 14544
rect 22652 14492 22704 14544
rect 23204 14492 23256 14544
rect 18880 14467 18932 14476
rect 18880 14433 18914 14467
rect 18914 14433 18932 14467
rect 18880 14424 18932 14433
rect 19432 14424 19484 14476
rect 18236 14356 18288 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 20720 14356 20772 14408
rect 23940 14424 23992 14476
rect 23020 14356 23072 14408
rect 18328 14331 18380 14340
rect 18328 14297 18337 14331
rect 18337 14297 18371 14331
rect 18371 14297 18380 14331
rect 18328 14288 18380 14297
rect 22376 14288 22428 14340
rect 17592 14220 17644 14272
rect 20076 14220 20128 14272
rect 21916 14220 21968 14272
rect 23388 14220 23440 14272
rect 25044 14263 25096 14272
rect 25044 14229 25053 14263
rect 25053 14229 25087 14263
rect 25087 14229 25096 14263
rect 25044 14220 25096 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3056 14016 3108 14068
rect 6092 14016 6144 14068
rect 6828 14016 6880 14068
rect 7932 14016 7984 14068
rect 8300 14016 8352 14068
rect 9036 14016 9088 14068
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12808 14016 12860 14068
rect 12992 14016 13044 14068
rect 14740 14016 14792 14068
rect 15476 14059 15528 14068
rect 15476 14025 15485 14059
rect 15485 14025 15519 14059
rect 15519 14025 15528 14059
rect 21364 14059 21416 14068
rect 15476 14016 15528 14025
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 8760 13880 8812 13932
rect 6184 13855 6236 13864
rect 1676 13744 1728 13796
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 6644 13812 6696 13864
rect 7840 13812 7892 13864
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 4896 13744 4948 13796
rect 7196 13744 7248 13796
rect 9128 13812 9180 13864
rect 11060 13880 11112 13932
rect 15568 13948 15620 14000
rect 15752 13948 15804 14000
rect 21364 14025 21373 14059
rect 21373 14025 21407 14059
rect 21407 14025 21416 14059
rect 21364 14016 21416 14025
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 22376 14016 22428 14068
rect 14188 13880 14240 13932
rect 16672 13948 16724 14000
rect 19432 13991 19484 14000
rect 19432 13957 19441 13991
rect 19441 13957 19475 13991
rect 19475 13957 19484 13991
rect 19432 13948 19484 13957
rect 23204 13948 23256 14000
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 23388 13880 23440 13932
rect 24032 13880 24084 13932
rect 12532 13812 12584 13864
rect 13452 13812 13504 13864
rect 15108 13812 15160 13864
rect 16948 13812 17000 13864
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 18144 13812 18196 13864
rect 13544 13744 13596 13796
rect 2228 13676 2280 13728
rect 5540 13676 5592 13728
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13912 13676 13964 13728
rect 14464 13719 14516 13728
rect 14464 13685 14473 13719
rect 14473 13685 14507 13719
rect 14507 13685 14516 13719
rect 14464 13676 14516 13685
rect 20996 13744 21048 13796
rect 21364 13744 21416 13796
rect 24124 13744 24176 13796
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 18144 13676 18196 13728
rect 20260 13719 20312 13728
rect 20260 13685 20269 13719
rect 20269 13685 20303 13719
rect 20303 13685 20312 13719
rect 20260 13676 20312 13685
rect 20536 13676 20588 13728
rect 21732 13676 21784 13728
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 25780 13676 25832 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 3148 13472 3200 13524
rect 4068 13472 4120 13524
rect 5448 13472 5500 13524
rect 6092 13472 6144 13524
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 9036 13515 9088 13524
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9036 13472 9088 13481
rect 2228 13404 2280 13456
rect 7748 13404 7800 13456
rect 12164 13404 12216 13456
rect 12624 13404 12676 13456
rect 12808 13472 12860 13524
rect 12992 13472 13044 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 18880 13472 18932 13524
rect 19248 13472 19300 13524
rect 20260 13472 20312 13524
rect 20444 13472 20496 13524
rect 20628 13472 20680 13524
rect 21364 13515 21416 13524
rect 21364 13481 21373 13515
rect 21373 13481 21407 13515
rect 21407 13481 21416 13515
rect 21364 13472 21416 13481
rect 21640 13472 21692 13524
rect 22652 13472 22704 13524
rect 24032 13472 24084 13524
rect 25872 13472 25924 13524
rect 14464 13404 14516 13456
rect 14740 13404 14792 13456
rect 19340 13447 19392 13456
rect 1860 13336 1912 13388
rect 4620 13336 4672 13388
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 5448 13336 5500 13388
rect 7472 13336 7524 13388
rect 8116 13336 8168 13388
rect 8760 13336 8812 13388
rect 9680 13336 9732 13388
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 13912 13336 13964 13388
rect 10140 13268 10192 13320
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10876 13268 10928 13320
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 15568 13336 15620 13388
rect 15936 13336 15988 13388
rect 16488 13336 16540 13388
rect 19340 13413 19349 13447
rect 19349 13413 19383 13447
rect 19383 13413 19392 13447
rect 19340 13404 19392 13413
rect 23388 13447 23440 13456
rect 23388 13413 23422 13447
rect 23422 13413 23440 13447
rect 23388 13404 23440 13413
rect 21548 13336 21600 13388
rect 25320 13379 25372 13388
rect 25320 13345 25329 13379
rect 25329 13345 25363 13379
rect 25363 13345 25372 13379
rect 25320 13336 25372 13345
rect 14464 13268 14516 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16580 13268 16632 13320
rect 20076 13268 20128 13320
rect 20628 13268 20680 13320
rect 21088 13268 21140 13320
rect 21916 13311 21968 13320
rect 21916 13277 21925 13311
rect 21925 13277 21959 13311
rect 21959 13277 21968 13311
rect 21916 13268 21968 13277
rect 1216 13132 1268 13184
rect 2044 13132 2096 13184
rect 3240 13132 3292 13184
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 19892 13200 19944 13252
rect 13176 13132 13228 13184
rect 16212 13132 16264 13184
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18144 13132 18196 13141
rect 18972 13175 19024 13184
rect 18972 13141 18981 13175
rect 18981 13141 19015 13175
rect 19015 13141 19024 13175
rect 18972 13132 19024 13141
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20536 13132 20588 13184
rect 21732 13132 21784 13184
rect 22284 13200 22336 13252
rect 23020 13200 23072 13252
rect 25780 13200 25832 13252
rect 24124 13132 24176 13184
rect 24952 13132 25004 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2688 12928 2740 12980
rect 3424 12928 3476 12980
rect 5356 12928 5408 12980
rect 7196 12971 7248 12980
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 10416 12928 10468 12980
rect 12532 12928 12584 12980
rect 13544 12928 13596 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 16672 12928 16724 12980
rect 18512 12928 18564 12980
rect 20628 12971 20680 12980
rect 20628 12937 20637 12971
rect 20637 12937 20671 12971
rect 20671 12937 20680 12971
rect 20628 12928 20680 12937
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21548 12928 21600 12980
rect 23388 12928 23440 12980
rect 25320 12971 25372 12980
rect 25320 12937 25329 12971
rect 25329 12937 25363 12971
rect 25363 12937 25372 12971
rect 25320 12928 25372 12937
rect 2044 12860 2096 12912
rect 2228 12860 2280 12912
rect 5632 12860 5684 12912
rect 6920 12860 6972 12912
rect 16212 12860 16264 12912
rect 16396 12860 16448 12912
rect 1676 12792 1728 12844
rect 3424 12792 3476 12844
rect 3608 12792 3660 12844
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 3240 12724 3292 12776
rect 5356 12792 5408 12844
rect 5540 12792 5592 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 8392 12792 8444 12844
rect 13728 12792 13780 12844
rect 18144 12792 18196 12844
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 19064 12860 19116 12912
rect 20076 12792 20128 12844
rect 22652 12835 22704 12844
rect 22652 12801 22661 12835
rect 22661 12801 22695 12835
rect 22695 12801 22704 12835
rect 22652 12792 22704 12801
rect 24124 12792 24176 12844
rect 24860 12792 24912 12844
rect 4988 12724 5040 12776
rect 8944 12724 8996 12776
rect 9864 12724 9916 12776
rect 10876 12724 10928 12776
rect 14004 12724 14056 12776
rect 14188 12767 14240 12776
rect 14188 12733 14222 12767
rect 14222 12733 14240 12767
rect 14188 12724 14240 12733
rect 18696 12724 18748 12776
rect 21916 12767 21968 12776
rect 21916 12733 21925 12767
rect 21925 12733 21959 12767
rect 21959 12733 21968 12767
rect 21916 12724 21968 12733
rect 23388 12724 23440 12776
rect 24676 12724 24728 12776
rect 2780 12656 2832 12708
rect 5080 12699 5132 12708
rect 5080 12665 5089 12699
rect 5089 12665 5123 12699
rect 5123 12665 5132 12699
rect 5080 12656 5132 12665
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 2320 12588 2372 12597
rect 3240 12588 3292 12640
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 3976 12588 4028 12597
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 6920 12588 6972 12640
rect 9128 12699 9180 12708
rect 9128 12665 9137 12699
rect 9137 12665 9171 12699
rect 9171 12665 9180 12699
rect 9128 12656 9180 12665
rect 10784 12656 10836 12708
rect 18512 12699 18564 12708
rect 11060 12588 11112 12640
rect 11980 12588 12032 12640
rect 12164 12588 12216 12640
rect 14464 12588 14516 12640
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 16396 12588 16448 12597
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 16948 12588 17000 12640
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 20168 12656 20220 12708
rect 20628 12588 20680 12640
rect 22008 12631 22060 12640
rect 22008 12597 22017 12631
rect 22017 12597 22051 12631
rect 22051 12597 22060 12631
rect 22008 12588 22060 12597
rect 22192 12588 22244 12640
rect 23664 12588 23716 12640
rect 24032 12631 24084 12640
rect 24032 12597 24041 12631
rect 24041 12597 24075 12631
rect 24075 12597 24084 12631
rect 24032 12588 24084 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1400 12384 1452 12436
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 8392 12427 8444 12436
rect 8392 12393 8401 12427
rect 8401 12393 8435 12427
rect 8435 12393 8444 12427
rect 8392 12384 8444 12393
rect 8944 12427 8996 12436
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 2044 12316 2096 12368
rect 2504 12248 2556 12300
rect 2872 12248 2924 12300
rect 4620 12316 4672 12368
rect 4344 12291 4396 12300
rect 4344 12257 4378 12291
rect 4378 12257 4396 12291
rect 6092 12291 6144 12300
rect 4344 12248 4396 12257
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 7564 12316 7616 12368
rect 11336 12316 11388 12368
rect 13360 12384 13412 12436
rect 14740 12384 14792 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 15752 12384 15804 12436
rect 16948 12384 17000 12436
rect 19248 12384 19300 12436
rect 19340 12384 19392 12436
rect 20076 12427 20128 12436
rect 20076 12393 20085 12427
rect 20085 12393 20119 12427
rect 20119 12393 20128 12427
rect 20076 12384 20128 12393
rect 20168 12384 20220 12436
rect 21180 12384 21232 12436
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 22192 12384 22244 12436
rect 22284 12384 22336 12436
rect 23388 12384 23440 12436
rect 7288 12291 7340 12300
rect 7288 12257 7322 12291
rect 7322 12257 7340 12291
rect 7288 12248 7340 12257
rect 9404 12248 9456 12300
rect 9772 12248 9824 12300
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 9956 12180 10008 12232
rect 11060 12248 11112 12300
rect 14004 12316 14056 12368
rect 16764 12316 16816 12368
rect 22560 12316 22612 12368
rect 13176 12291 13228 12300
rect 13176 12257 13210 12291
rect 13210 12257 13228 12291
rect 13176 12248 13228 12257
rect 14740 12248 14792 12300
rect 19340 12291 19392 12300
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 20076 12248 20128 12300
rect 20444 12248 20496 12300
rect 20904 12291 20956 12300
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 12072 12180 12124 12232
rect 16580 12180 16632 12232
rect 18236 12180 18288 12232
rect 18512 12180 18564 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22376 12248 22428 12300
rect 23020 12248 23072 12300
rect 19524 12180 19576 12189
rect 20996 12180 21048 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 22560 12180 22612 12232
rect 2228 12112 2280 12164
rect 17776 12112 17828 12164
rect 22652 12112 22704 12164
rect 22836 12180 22888 12232
rect 24952 12316 25004 12368
rect 24124 12291 24176 12300
rect 24124 12257 24158 12291
rect 24158 12257 24176 12291
rect 24124 12248 24176 12257
rect 2136 12044 2188 12096
rect 2412 12044 2464 12096
rect 3976 12044 4028 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 14188 12044 14240 12096
rect 15568 12044 15620 12096
rect 16580 12044 16632 12096
rect 18604 12044 18656 12096
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 20720 12044 20772 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22836 12044 22888 12096
rect 25228 12087 25280 12096
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 25228 12044 25280 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2320 11840 2372 11892
rect 4528 11840 4580 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 9772 11840 9824 11892
rect 9956 11883 10008 11892
rect 9956 11849 9965 11883
rect 9965 11849 9999 11883
rect 9999 11849 10008 11883
rect 9956 11840 10008 11849
rect 10140 11840 10192 11892
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 12808 11840 12860 11892
rect 13176 11840 13228 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 16212 11840 16264 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17592 11840 17644 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 19432 11840 19484 11892
rect 22652 11840 22704 11892
rect 24860 11840 24912 11892
rect 2044 11772 2096 11824
rect 4068 11772 4120 11824
rect 4344 11772 4396 11824
rect 4712 11772 4764 11824
rect 4896 11772 4948 11824
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 3976 11747 4028 11756
rect 2320 11704 2372 11713
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 5172 11704 5224 11756
rect 7748 11815 7800 11824
rect 7748 11781 7757 11815
rect 7757 11781 7791 11815
rect 7791 11781 7800 11815
rect 7748 11772 7800 11781
rect 6828 11747 6880 11756
rect 3884 11636 3936 11688
rect 4344 11636 4396 11688
rect 4528 11636 4580 11688
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 8208 11704 8260 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 9496 11704 9548 11756
rect 11244 11772 11296 11824
rect 12440 11815 12492 11824
rect 12440 11781 12449 11815
rect 12449 11781 12483 11815
rect 12483 11781 12492 11815
rect 12440 11772 12492 11781
rect 19984 11772 20036 11824
rect 20444 11772 20496 11824
rect 25320 11815 25372 11824
rect 25320 11781 25329 11815
rect 25329 11781 25363 11815
rect 25363 11781 25372 11815
rect 25320 11772 25372 11781
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 9036 11636 9088 11688
rect 5448 11568 5500 11620
rect 6184 11568 6236 11620
rect 11060 11704 11112 11756
rect 12532 11704 12584 11756
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 23388 11704 23440 11756
rect 12624 11636 12676 11688
rect 13268 11636 13320 11688
rect 14004 11636 14056 11688
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 18328 11636 18380 11688
rect 18420 11636 18472 11688
rect 20536 11636 20588 11688
rect 25228 11636 25280 11688
rect 15292 11568 15344 11620
rect 1584 11500 1636 11552
rect 2044 11500 2096 11552
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4896 11500 4948 11552
rect 5080 11500 5132 11552
rect 7564 11500 7616 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 9956 11500 10008 11552
rect 10140 11500 10192 11552
rect 10784 11500 10836 11552
rect 12808 11500 12860 11552
rect 13268 11500 13320 11552
rect 20444 11500 20496 11552
rect 21088 11568 21140 11620
rect 24308 11568 24360 11620
rect 21272 11500 21324 11552
rect 22560 11500 22612 11552
rect 23020 11500 23072 11552
rect 25688 11543 25740 11552
rect 25688 11509 25697 11543
rect 25697 11509 25731 11543
rect 25731 11509 25740 11543
rect 25688 11500 25740 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1492 11296 1544 11348
rect 2688 11296 2740 11348
rect 3148 11296 3200 11348
rect 3884 11296 3936 11348
rect 4436 11296 4488 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 8484 11296 8536 11348
rect 10692 11296 10744 11348
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 13268 11339 13320 11348
rect 1584 11271 1636 11280
rect 1584 11237 1593 11271
rect 1593 11237 1627 11271
rect 1627 11237 1636 11271
rect 1584 11228 1636 11237
rect 2320 11228 2372 11280
rect 4160 11228 4212 11280
rect 4896 11228 4948 11280
rect 6644 11228 6696 11280
rect 8208 11228 8260 11280
rect 9956 11228 10008 11280
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 1216 11160 1268 11212
rect 1492 11160 1544 11212
rect 2412 11160 2464 11212
rect 3884 11203 3936 11212
rect 3884 11169 3893 11203
rect 3893 11169 3927 11203
rect 3927 11169 3936 11203
rect 3884 11160 3936 11169
rect 2228 11092 2280 11144
rect 1860 11024 1912 11076
rect 4528 11067 4580 11076
rect 4528 11033 4537 11067
rect 4537 11033 4571 11067
rect 4571 11033 4580 11067
rect 9404 11160 9456 11212
rect 9864 11160 9916 11212
rect 12624 11228 12676 11280
rect 14004 11228 14056 11280
rect 15292 11296 15344 11348
rect 16948 11296 17000 11348
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 18328 11339 18380 11348
rect 18328 11305 18337 11339
rect 18337 11305 18371 11339
rect 18371 11305 18380 11339
rect 18328 11296 18380 11305
rect 18788 11296 18840 11348
rect 19340 11296 19392 11348
rect 20260 11296 20312 11348
rect 20904 11296 20956 11348
rect 21732 11296 21784 11348
rect 22100 11296 22152 11348
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 23480 11296 23532 11348
rect 15752 11228 15804 11280
rect 20996 11228 21048 11280
rect 10968 11203 11020 11212
rect 10968 11169 11002 11203
rect 11002 11169 11020 11203
rect 10968 11160 11020 11169
rect 13268 11160 13320 11212
rect 13360 11160 13412 11212
rect 13820 11203 13872 11212
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 16120 11160 16172 11212
rect 17592 11160 17644 11212
rect 18328 11160 18380 11212
rect 18696 11160 18748 11212
rect 19524 11160 19576 11212
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 22468 11228 22520 11280
rect 22192 11203 22244 11212
rect 19708 11160 19760 11169
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 22652 11160 22704 11212
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5540 11092 5592 11144
rect 4528 11024 4580 11033
rect 5080 11024 5132 11076
rect 6460 11092 6512 11144
rect 7380 11092 7432 11144
rect 7656 11092 7708 11144
rect 8116 11092 8168 11144
rect 6828 11024 6880 11076
rect 13728 11092 13780 11144
rect 10140 11024 10192 11076
rect 11704 11024 11756 11076
rect 4436 10956 4488 11008
rect 7840 10956 7892 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 9680 10956 9732 11008
rect 12072 10956 12124 11008
rect 12808 10956 12860 11008
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 14372 11092 14424 11144
rect 16580 11092 16632 11144
rect 15476 11024 15528 11076
rect 19432 11024 19484 11076
rect 20444 11092 20496 11144
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 24032 11296 24084 11348
rect 24124 11296 24176 11348
rect 25412 11296 25464 11348
rect 24952 11271 25004 11280
rect 24952 11237 24961 11271
rect 24961 11237 24995 11271
rect 24995 11237 25004 11271
rect 25688 11271 25740 11280
rect 24952 11228 25004 11237
rect 25688 11237 25697 11271
rect 25697 11237 25731 11271
rect 25731 11237 25740 11271
rect 25688 11228 25740 11237
rect 25596 11160 25648 11212
rect 22468 11092 22520 11101
rect 23940 11092 23992 11144
rect 24308 11092 24360 11144
rect 21824 11067 21876 11076
rect 21824 11033 21833 11067
rect 21833 11033 21867 11067
rect 21867 11033 21876 11067
rect 21824 11024 21876 11033
rect 23756 11024 23808 11076
rect 14372 10956 14424 11008
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 16948 10956 17000 11008
rect 20352 10956 20404 11008
rect 25044 10956 25096 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2228 10752 2280 10804
rect 4068 10795 4120 10804
rect 4068 10761 4077 10795
rect 4077 10761 4111 10795
rect 4111 10761 4120 10795
rect 4068 10752 4120 10761
rect 4896 10752 4948 10804
rect 5172 10752 5224 10804
rect 5448 10752 5500 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9312 10752 9364 10804
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 15384 10752 15436 10804
rect 16488 10752 16540 10804
rect 17224 10752 17276 10804
rect 19432 10752 19484 10804
rect 19524 10752 19576 10804
rect 21088 10795 21140 10804
rect 3976 10684 4028 10736
rect 6644 10727 6696 10736
rect 6644 10693 6653 10727
rect 6653 10693 6687 10727
rect 6687 10693 6696 10727
rect 6644 10684 6696 10693
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 4436 10616 4488 10668
rect 4620 10548 4672 10600
rect 5356 10548 5408 10600
rect 7380 10548 7432 10600
rect 8116 10548 8168 10600
rect 8208 10548 8260 10600
rect 10232 10616 10284 10668
rect 10784 10684 10836 10736
rect 11612 10684 11664 10736
rect 17500 10684 17552 10736
rect 21088 10761 21097 10795
rect 21097 10761 21131 10795
rect 21131 10761 21140 10795
rect 21088 10752 21140 10761
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 12532 10616 12584 10668
rect 13452 10616 13504 10668
rect 14004 10616 14056 10668
rect 15568 10616 15620 10668
rect 17316 10616 17368 10668
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 10048 10548 10100 10600
rect 14832 10548 14884 10600
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 16948 10548 17000 10600
rect 18052 10548 18104 10600
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 19064 10548 19116 10600
rect 20536 10548 20588 10600
rect 22468 10616 22520 10668
rect 23572 10616 23624 10668
rect 2688 10480 2740 10532
rect 3424 10480 3476 10532
rect 6920 10480 6972 10532
rect 11152 10480 11204 10532
rect 15292 10480 15344 10532
rect 17408 10480 17460 10532
rect 19984 10523 20036 10532
rect 19984 10489 20018 10523
rect 20018 10489 20036 10523
rect 19984 10480 20036 10489
rect 24952 10548 25004 10600
rect 6460 10412 6512 10464
rect 7840 10412 7892 10464
rect 10048 10412 10100 10464
rect 10692 10412 10744 10464
rect 11060 10412 11112 10464
rect 11980 10412 12032 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13360 10412 13412 10464
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 15844 10412 15896 10464
rect 17132 10412 17184 10464
rect 17592 10412 17644 10464
rect 17868 10412 17920 10464
rect 21732 10412 21784 10464
rect 22836 10480 22888 10532
rect 23572 10480 23624 10532
rect 24216 10523 24268 10532
rect 24216 10489 24250 10523
rect 24250 10489 24268 10523
rect 24216 10480 24268 10489
rect 21916 10412 21968 10464
rect 22652 10412 22704 10464
rect 25320 10455 25372 10464
rect 25320 10421 25329 10455
rect 25329 10421 25363 10455
rect 25363 10421 25372 10455
rect 25320 10412 25372 10421
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2688 10208 2740 10260
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 4896 10208 4948 10260
rect 6920 10208 6972 10260
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 9036 10251 9088 10260
rect 7104 10208 7156 10217
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 10784 10208 10836 10260
rect 14372 10208 14424 10260
rect 15660 10208 15712 10260
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 18512 10208 18564 10260
rect 19248 10208 19300 10260
rect 20168 10208 20220 10260
rect 22008 10208 22060 10260
rect 22192 10208 22244 10260
rect 22652 10208 22704 10260
rect 23296 10208 23348 10260
rect 23940 10251 23992 10260
rect 23940 10217 23949 10251
rect 23949 10217 23983 10251
rect 23983 10217 23992 10251
rect 23940 10208 23992 10217
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 24308 10208 24360 10260
rect 25228 10208 25280 10260
rect 25780 10251 25832 10260
rect 25780 10217 25789 10251
rect 25789 10217 25823 10251
rect 25823 10217 25832 10251
rect 25780 10208 25832 10217
rect 1860 10140 1912 10192
rect 2780 10140 2832 10192
rect 5448 10140 5500 10192
rect 10048 10140 10100 10192
rect 14464 10140 14516 10192
rect 2964 10072 3016 10124
rect 3516 10072 3568 10124
rect 4436 10072 4488 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 7656 10115 7708 10124
rect 7656 10081 7690 10115
rect 7690 10081 7708 10115
rect 7656 10072 7708 10081
rect 9956 10072 10008 10124
rect 10876 10115 10928 10124
rect 10876 10081 10910 10115
rect 10910 10081 10928 10115
rect 10876 10072 10928 10081
rect 12072 10072 12124 10124
rect 17316 10140 17368 10192
rect 17500 10140 17552 10192
rect 17776 10140 17828 10192
rect 18972 10140 19024 10192
rect 22928 10140 22980 10192
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 20352 10072 20404 10124
rect 21180 10072 21232 10124
rect 21364 10072 21416 10124
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 12624 10004 12676 10056
rect 8760 9979 8812 9988
rect 8760 9945 8769 9979
rect 8769 9945 8803 9979
rect 8803 9945 8812 9979
rect 8760 9936 8812 9945
rect 9680 9936 9732 9988
rect 2320 9868 2372 9920
rect 3148 9868 3200 9920
rect 4804 9868 4856 9920
rect 8576 9868 8628 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 10048 9868 10100 9920
rect 12348 9936 12400 9988
rect 11980 9911 12032 9920
rect 11980 9877 11989 9911
rect 11989 9877 12023 9911
rect 12023 9877 12032 9911
rect 11980 9868 12032 9877
rect 12164 9868 12216 9920
rect 12532 9868 12584 9920
rect 15844 10004 15896 10056
rect 19524 10004 19576 10056
rect 19984 10004 20036 10056
rect 21272 10004 21324 10056
rect 22468 10072 22520 10124
rect 15292 9936 15344 9988
rect 14188 9868 14240 9920
rect 15384 9868 15436 9920
rect 15936 9868 15988 9920
rect 16120 9868 16172 9920
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 20260 9911 20312 9920
rect 20260 9877 20269 9911
rect 20269 9877 20303 9911
rect 20303 9877 20312 9911
rect 20260 9868 20312 9877
rect 21640 9868 21692 9920
rect 22836 9911 22888 9920
rect 22836 9877 22845 9911
rect 22845 9877 22879 9911
rect 22879 9877 22888 9911
rect 22836 9868 22888 9877
rect 23940 10072 23992 10124
rect 24860 10072 24912 10124
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 24216 9868 24268 9920
rect 24768 9868 24820 9920
rect 25596 9868 25648 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 5448 9664 5500 9716
rect 1952 9596 2004 9648
rect 4528 9596 4580 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 3884 9528 3936 9580
rect 7288 9664 7340 9716
rect 12072 9664 12124 9716
rect 12624 9664 12676 9716
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 20168 9664 20220 9716
rect 23940 9664 23992 9716
rect 24032 9664 24084 9716
rect 24676 9664 24728 9716
rect 25228 9664 25280 9716
rect 25780 9664 25832 9716
rect 10876 9596 10928 9648
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 12164 9596 12216 9648
rect 12808 9596 12860 9648
rect 13176 9596 13228 9648
rect 14464 9639 14516 9648
rect 14464 9605 14473 9639
rect 14473 9605 14507 9639
rect 14507 9605 14516 9639
rect 14464 9596 14516 9605
rect 19432 9596 19484 9648
rect 24952 9596 25004 9648
rect 2964 9460 3016 9512
rect 10692 9460 10744 9512
rect 12072 9528 12124 9580
rect 12348 9460 12400 9512
rect 12440 9460 12492 9512
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 17960 9528 18012 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 22836 9528 22888 9580
rect 24860 9528 24912 9580
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 4896 9392 4948 9444
rect 6368 9392 6420 9444
rect 8668 9392 8720 9444
rect 12164 9435 12216 9444
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 16212 9460 16264 9512
rect 19340 9460 19392 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 22100 9460 22152 9512
rect 23388 9460 23440 9512
rect 25596 9460 25648 9512
rect 16396 9392 16448 9444
rect 20260 9392 20312 9444
rect 23296 9392 23348 9444
rect 23940 9392 23992 9444
rect 2872 9324 2924 9376
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 3424 9324 3476 9376
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 5448 9324 5500 9376
rect 7656 9324 7708 9376
rect 9404 9324 9456 9376
rect 10784 9324 10836 9376
rect 11060 9324 11112 9376
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 14832 9324 14884 9376
rect 17316 9324 17368 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 19340 9324 19392 9376
rect 19524 9324 19576 9376
rect 20352 9324 20404 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21364 9324 21416 9376
rect 22008 9367 22060 9376
rect 22008 9333 22017 9367
rect 22017 9333 22051 9367
rect 22051 9333 22060 9367
rect 22008 9324 22060 9333
rect 22468 9367 22520 9376
rect 22468 9333 22477 9367
rect 22477 9333 22511 9367
rect 22511 9333 22520 9367
rect 22468 9324 22520 9333
rect 22560 9324 22612 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2136 9120 2188 9172
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 4988 9120 5040 9172
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 9220 9120 9272 9172
rect 10692 9120 10744 9172
rect 11796 9120 11848 9172
rect 13820 9120 13872 9172
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 16856 9163 16908 9172
rect 15752 9120 15804 9129
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 17868 9120 17920 9172
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 19156 9120 19208 9172
rect 20628 9163 20680 9172
rect 20628 9129 20637 9163
rect 20637 9129 20671 9163
rect 20671 9129 20680 9163
rect 20628 9120 20680 9129
rect 20904 9120 20956 9172
rect 22928 9163 22980 9172
rect 22928 9129 22937 9163
rect 22937 9129 22971 9163
rect 22971 9129 22980 9163
rect 22928 9120 22980 9129
rect 23848 9120 23900 9172
rect 24860 9163 24912 9172
rect 2504 9052 2556 9104
rect 2044 8984 2096 9036
rect 3148 8984 3200 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 2688 8848 2740 8900
rect 4712 9052 4764 9104
rect 10876 9052 10928 9104
rect 12992 9052 13044 9104
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 6828 8984 6880 9036
rect 7380 8984 7432 9036
rect 7840 8984 7892 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9956 8984 10008 9036
rect 3976 8916 4028 8968
rect 5540 8916 5592 8968
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 17684 9052 17736 9104
rect 20168 9052 20220 9104
rect 21732 9095 21784 9104
rect 21732 9061 21741 9095
rect 21741 9061 21775 9095
rect 21775 9061 21784 9095
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 25136 9120 25188 9172
rect 25596 9163 25648 9172
rect 25596 9129 25605 9163
rect 25605 9129 25639 9163
rect 25639 9129 25648 9163
rect 25596 9120 25648 9129
rect 21732 9052 21784 9061
rect 13268 8984 13320 9036
rect 13452 8984 13504 9036
rect 19432 8984 19484 9036
rect 7104 8891 7156 8900
rect 7104 8857 7113 8891
rect 7113 8857 7147 8891
rect 7147 8857 7156 8891
rect 7104 8848 7156 8857
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 17316 8916 17368 8968
rect 19984 8984 20036 9036
rect 23480 8984 23532 9036
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 21456 8916 21508 8968
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 13268 8848 13320 8900
rect 14372 8848 14424 8900
rect 22836 8916 22888 8968
rect 25688 9052 25740 9104
rect 25044 9027 25096 9036
rect 25044 8993 25053 9027
rect 25053 8993 25087 9027
rect 25087 8993 25096 9027
rect 25044 8984 25096 8993
rect 25872 8916 25924 8968
rect 24216 8848 24268 8900
rect 24308 8848 24360 8900
rect 24860 8848 24912 8900
rect 3884 8780 3936 8832
rect 4804 8780 4856 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 5448 8780 5500 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 12164 8780 12216 8832
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 19524 8780 19576 8832
rect 20720 8780 20772 8832
rect 22836 8780 22888 8832
rect 23388 8780 23440 8832
rect 23848 8780 23900 8832
rect 24032 8780 24084 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2872 8576 2924 8628
rect 2964 8576 3016 8628
rect 4620 8576 4672 8628
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 4068 8508 4120 8560
rect 4528 8508 4580 8560
rect 5356 8440 5408 8492
rect 7104 8440 7156 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 10876 8576 10928 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12072 8576 12124 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 15844 8576 15896 8628
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 17868 8576 17920 8628
rect 19892 8576 19944 8628
rect 20168 8619 20220 8628
rect 20168 8585 20177 8619
rect 20177 8585 20211 8619
rect 20211 8585 20220 8619
rect 20168 8576 20220 8585
rect 21732 8576 21784 8628
rect 22100 8576 22152 8628
rect 23940 8576 23992 8628
rect 25688 8619 25740 8628
rect 25688 8585 25697 8619
rect 25697 8585 25731 8619
rect 25731 8585 25740 8619
rect 25688 8576 25740 8585
rect 9772 8508 9824 8560
rect 1676 8372 1728 8424
rect 2136 8415 2188 8424
rect 2136 8381 2170 8415
rect 2170 8381 2188 8415
rect 2136 8372 2188 8381
rect 4712 8372 4764 8424
rect 9220 8372 9272 8424
rect 3148 8304 3200 8356
rect 4620 8304 4672 8356
rect 8852 8304 8904 8356
rect 11980 8440 12032 8492
rect 10232 8372 10284 8424
rect 10784 8372 10836 8424
rect 10968 8304 11020 8356
rect 12164 8372 12216 8424
rect 16396 8440 16448 8492
rect 16580 8440 16632 8492
rect 14372 8372 14424 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 12808 8304 12860 8356
rect 13084 8304 13136 8356
rect 13728 8304 13780 8356
rect 13912 8304 13964 8356
rect 18236 8347 18288 8356
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 7840 8236 7892 8288
rect 9220 8236 9272 8288
rect 12440 8236 12492 8288
rect 13636 8236 13688 8288
rect 13820 8236 13872 8288
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 18236 8313 18245 8347
rect 18245 8313 18279 8347
rect 18279 8313 18288 8347
rect 19064 8347 19116 8356
rect 18236 8304 18288 8313
rect 19064 8313 19076 8347
rect 19076 8313 19116 8347
rect 19064 8304 19116 8313
rect 17868 8236 17920 8288
rect 19156 8236 19208 8288
rect 19524 8372 19576 8424
rect 21088 8372 21140 8424
rect 23296 8440 23348 8492
rect 25044 8440 25096 8492
rect 23480 8415 23532 8424
rect 23480 8381 23489 8415
rect 23489 8381 23523 8415
rect 23523 8381 23532 8415
rect 23480 8372 23532 8381
rect 20352 8236 20404 8288
rect 20904 8304 20956 8356
rect 22468 8304 22520 8356
rect 22836 8236 22888 8288
rect 23296 8236 23348 8288
rect 24216 8304 24268 8356
rect 24032 8236 24084 8288
rect 25688 8236 25740 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2136 8032 2188 8084
rect 3976 8032 4028 8084
rect 4252 8032 4304 8084
rect 4896 8032 4948 8084
rect 5356 8032 5408 8084
rect 7380 8032 7432 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10968 8032 11020 8084
rect 12532 8032 12584 8084
rect 12992 8032 13044 8084
rect 13268 8032 13320 8084
rect 2044 7964 2096 8016
rect 3332 7964 3384 8016
rect 5172 7964 5224 8016
rect 5632 7964 5684 8016
rect 7932 7964 7984 8016
rect 9588 7964 9640 8016
rect 13636 8007 13688 8016
rect 3516 7939 3568 7948
rect 2228 7828 2280 7880
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 2412 7803 2464 7812
rect 2412 7769 2421 7803
rect 2421 7769 2455 7803
rect 2455 7769 2464 7803
rect 2412 7760 2464 7769
rect 2504 7760 2556 7812
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 6184 7896 6236 7948
rect 6920 7896 6972 7948
rect 10324 7896 10376 7948
rect 11796 7896 11848 7948
rect 3976 7828 4028 7880
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9956 7828 10008 7880
rect 13636 7973 13645 8007
rect 13645 7973 13679 8007
rect 13679 7973 13688 8007
rect 13636 7964 13688 7973
rect 13452 7896 13504 7948
rect 14372 8032 14424 8084
rect 15660 8032 15712 8084
rect 16764 8032 16816 8084
rect 18880 8032 18932 8084
rect 20168 8032 20220 8084
rect 20352 8032 20404 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 22744 8032 22796 8084
rect 24676 8075 24728 8084
rect 24676 8041 24685 8075
rect 24685 8041 24719 8075
rect 24719 8041 24728 8075
rect 24676 8032 24728 8041
rect 25688 8032 25740 8084
rect 15752 8007 15804 8016
rect 15752 7973 15761 8007
rect 15761 7973 15795 8007
rect 15795 7973 15804 8007
rect 15752 7964 15804 7973
rect 16580 8007 16632 8016
rect 16580 7973 16614 8007
rect 16614 7973 16632 8007
rect 16580 7964 16632 7973
rect 19432 7964 19484 8016
rect 23112 7964 23164 8016
rect 13268 7828 13320 7880
rect 14832 7896 14884 7948
rect 16856 7896 16908 7948
rect 17776 7896 17828 7948
rect 18328 7896 18380 7948
rect 19064 7896 19116 7948
rect 8668 7760 8720 7812
rect 10140 7760 10192 7812
rect 13452 7760 13504 7812
rect 1584 7692 1636 7744
rect 3056 7692 3108 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6552 7692 6604 7744
rect 7012 7692 7064 7744
rect 7196 7692 7248 7744
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 12440 7692 12492 7744
rect 15844 7828 15896 7880
rect 16028 7828 16080 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20904 7896 20956 7948
rect 23204 7896 23256 7948
rect 25504 7896 25556 7948
rect 21916 7828 21968 7880
rect 19248 7760 19300 7812
rect 20352 7803 20404 7812
rect 20352 7769 20361 7803
rect 20361 7769 20395 7803
rect 20395 7769 20404 7803
rect 20352 7760 20404 7769
rect 23664 7828 23716 7880
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 14832 7692 14884 7744
rect 18236 7692 18288 7744
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 23296 7692 23348 7744
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2872 7488 2924 7540
rect 3056 7488 3108 7540
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 4988 7488 5040 7540
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 2504 7420 2556 7472
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 5264 7352 5316 7404
rect 5540 7352 5592 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 7840 7352 7892 7404
rect 2872 7284 2924 7336
rect 8576 7488 8628 7540
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 10324 7531 10376 7540
rect 8668 7488 8720 7497
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 11060 7488 11112 7540
rect 10140 7420 10192 7472
rect 12164 7420 12216 7472
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 11704 7352 11756 7404
rect 12532 7488 12584 7540
rect 16212 7488 16264 7540
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18880 7488 18932 7540
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 19984 7488 20036 7540
rect 21916 7531 21968 7540
rect 21916 7497 21925 7531
rect 21925 7497 21959 7531
rect 21959 7497 21968 7531
rect 21916 7488 21968 7497
rect 23388 7488 23440 7540
rect 23940 7488 23992 7540
rect 24032 7488 24084 7540
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 16764 7420 16816 7472
rect 16212 7352 16264 7404
rect 18236 7352 18288 7404
rect 18880 7352 18932 7404
rect 20168 7352 20220 7404
rect 24216 7420 24268 7472
rect 24676 7352 24728 7404
rect 9220 7284 9272 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 13636 7284 13688 7336
rect 13820 7327 13872 7336
rect 13820 7293 13854 7327
rect 13854 7293 13872 7327
rect 13820 7284 13872 7293
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 18052 7284 18104 7336
rect 20628 7284 20680 7336
rect 4344 7216 4396 7268
rect 6000 7216 6052 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 2136 7148 2188 7200
rect 3332 7148 3384 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 6184 7148 6236 7200
rect 6920 7148 6972 7200
rect 7840 7148 7892 7200
rect 9496 7148 9548 7200
rect 9588 7148 9640 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 10876 7148 10928 7200
rect 13912 7216 13964 7268
rect 16672 7216 16724 7268
rect 17776 7216 17828 7268
rect 23296 7216 23348 7268
rect 24860 7216 24912 7268
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 12624 7191 12676 7200
rect 12624 7157 12633 7191
rect 12633 7157 12667 7191
rect 12667 7157 12676 7191
rect 12624 7148 12676 7157
rect 12808 7148 12860 7200
rect 13452 7148 13504 7200
rect 14372 7148 14424 7200
rect 15568 7148 15620 7200
rect 16028 7148 16080 7200
rect 16488 7148 16540 7200
rect 18328 7148 18380 7200
rect 20352 7148 20404 7200
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 22100 7148 22152 7200
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 26148 7216 26200 7268
rect 25504 7148 25556 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3424 6944 3476 6996
rect 5080 6987 5132 6996
rect 5080 6953 5089 6987
rect 5089 6953 5123 6987
rect 5123 6953 5132 6987
rect 5080 6944 5132 6953
rect 5816 6944 5868 6996
rect 6000 6944 6052 6996
rect 1492 6876 1544 6928
rect 2688 6876 2740 6928
rect 5540 6876 5592 6928
rect 8208 6944 8260 6996
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 12440 6944 12492 6996
rect 13268 6987 13320 6996
rect 13268 6953 13277 6987
rect 13277 6953 13311 6987
rect 13311 6953 13320 6987
rect 13268 6944 13320 6953
rect 16672 6987 16724 6996
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5356 6808 5408 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2596 6740 2648 6792
rect 4160 6740 4212 6792
rect 5264 6740 5316 6792
rect 1768 6672 1820 6724
rect 6184 6808 6236 6860
rect 6460 6808 6512 6860
rect 6644 6808 6696 6860
rect 9864 6876 9916 6928
rect 14096 6876 14148 6928
rect 14740 6876 14792 6928
rect 16672 6953 16681 6987
rect 16681 6953 16715 6987
rect 16715 6953 16724 6987
rect 16672 6944 16724 6953
rect 17040 6987 17092 6996
rect 17040 6953 17049 6987
rect 17049 6953 17083 6987
rect 17083 6953 17092 6987
rect 17040 6944 17092 6953
rect 19524 6944 19576 6996
rect 20628 6944 20680 6996
rect 22284 6944 22336 6996
rect 17224 6876 17276 6928
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 8576 6808 8628 6860
rect 9588 6808 9640 6860
rect 9772 6808 9824 6860
rect 10232 6851 10284 6860
rect 10232 6817 10255 6851
rect 10255 6817 10284 6851
rect 10232 6808 10284 6817
rect 11428 6808 11480 6860
rect 11704 6808 11756 6860
rect 11888 6808 11940 6860
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 16580 6808 16632 6860
rect 18236 6876 18288 6928
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 19340 6808 19392 6860
rect 20444 6808 20496 6860
rect 20996 6808 21048 6860
rect 21548 6808 21600 6860
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 8208 6740 8260 6792
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 12072 6740 12124 6792
rect 13820 6740 13872 6792
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 11060 6672 11112 6724
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 14188 6672 14240 6724
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 18236 6783 18288 6792
rect 17224 6740 17276 6749
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 20076 6740 20128 6792
rect 22100 6808 22152 6860
rect 23204 6808 23256 6860
rect 23388 6851 23440 6860
rect 23388 6817 23422 6851
rect 23422 6817 23440 6851
rect 23388 6808 23440 6817
rect 25320 6851 25372 6860
rect 25320 6817 25329 6851
rect 25329 6817 25363 6851
rect 25363 6817 25372 6851
rect 25320 6808 25372 6817
rect 17500 6672 17552 6724
rect 19248 6715 19300 6724
rect 19248 6681 19257 6715
rect 19257 6681 19291 6715
rect 19291 6681 19300 6715
rect 19248 6672 19300 6681
rect 24124 6672 24176 6724
rect 3424 6604 3476 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 7104 6604 7156 6656
rect 7380 6604 7432 6656
rect 7932 6604 7984 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 10876 6604 10928 6656
rect 11796 6604 11848 6656
rect 14832 6604 14884 6656
rect 17316 6604 17368 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 21272 6604 21324 6656
rect 22100 6604 22152 6656
rect 24216 6604 24268 6656
rect 24676 6604 24728 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 25228 6604 25280 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2320 6400 2372 6452
rect 5448 6400 5500 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 8300 6400 8352 6452
rect 8576 6443 8628 6452
rect 8576 6409 8585 6443
rect 8585 6409 8619 6443
rect 8619 6409 8628 6443
rect 8576 6400 8628 6409
rect 8852 6443 8904 6452
rect 8852 6409 8861 6443
rect 8861 6409 8895 6443
rect 8895 6409 8904 6443
rect 8852 6400 8904 6409
rect 10232 6400 10284 6452
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 12348 6400 12400 6452
rect 13176 6400 13228 6452
rect 14556 6400 14608 6452
rect 17224 6400 17276 6452
rect 19340 6400 19392 6452
rect 19524 6400 19576 6452
rect 20812 6443 20864 6452
rect 20812 6409 20821 6443
rect 20821 6409 20855 6443
rect 20855 6409 20864 6443
rect 20812 6400 20864 6409
rect 21548 6400 21600 6452
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 25688 6400 25740 6452
rect 5356 6332 5408 6384
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 15292 6332 15344 6384
rect 17500 6375 17552 6384
rect 17500 6341 17509 6375
rect 17509 6341 17543 6375
rect 17543 6341 17552 6375
rect 17500 6332 17552 6341
rect 20628 6332 20680 6384
rect 3516 6196 3568 6248
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5080 6196 5132 6205
rect 5264 6196 5316 6248
rect 2504 6128 2556 6180
rect 5448 6128 5500 6180
rect 6092 6196 6144 6248
rect 6736 6196 6788 6248
rect 7104 6196 7156 6248
rect 9036 6239 9088 6248
rect 9036 6205 9052 6239
rect 9052 6205 9086 6239
rect 9086 6205 9088 6239
rect 9036 6196 9088 6205
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 21272 6307 21324 6316
rect 21272 6273 21281 6307
rect 21281 6273 21315 6307
rect 21315 6273 21324 6307
rect 21272 6264 21324 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 24124 6307 24176 6316
rect 22192 6264 22244 6273
rect 9588 6196 9640 6248
rect 11152 6196 11204 6248
rect 12532 6196 12584 6248
rect 15568 6196 15620 6248
rect 17960 6196 18012 6248
rect 18420 6196 18472 6248
rect 20904 6196 20956 6248
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 25412 6307 25464 6316
rect 25412 6273 25421 6307
rect 25421 6273 25455 6307
rect 25455 6273 25464 6307
rect 25412 6264 25464 6273
rect 24032 6239 24084 6248
rect 24032 6205 24041 6239
rect 24041 6205 24075 6239
rect 24075 6205 24084 6239
rect 24032 6196 24084 6205
rect 25044 6196 25096 6248
rect 10048 6128 10100 6180
rect 2596 6060 2648 6112
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 3148 6060 3200 6112
rect 5080 6060 5132 6112
rect 6644 6060 6696 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 11888 6060 11940 6112
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 13636 6128 13688 6180
rect 15660 6171 15712 6180
rect 15660 6137 15669 6171
rect 15669 6137 15703 6171
rect 15703 6137 15712 6171
rect 15660 6128 15712 6137
rect 18512 6128 18564 6180
rect 19432 6128 19484 6180
rect 26516 6128 26568 6180
rect 13728 6060 13780 6112
rect 13820 6060 13872 6112
rect 20076 6060 20128 6112
rect 22560 6103 22612 6112
rect 22560 6069 22569 6103
rect 22569 6069 22603 6103
rect 22603 6069 22612 6103
rect 22560 6060 22612 6069
rect 23388 6060 23440 6112
rect 24676 6060 24728 6112
rect 25964 6103 26016 6112
rect 25964 6069 25973 6103
rect 25973 6069 26007 6103
rect 26007 6069 26016 6103
rect 25964 6060 26016 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2872 5856 2924 5908
rect 3884 5856 3936 5908
rect 4804 5856 4856 5908
rect 7196 5856 7248 5908
rect 7380 5856 7432 5908
rect 8208 5856 8260 5908
rect 3332 5831 3384 5840
rect 3332 5797 3341 5831
rect 3341 5797 3375 5831
rect 3375 5797 3384 5831
rect 3332 5788 3384 5797
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 1952 5763 2004 5772
rect 1952 5729 1986 5763
rect 1986 5729 2004 5763
rect 1952 5720 2004 5729
rect 3424 5720 3476 5772
rect 5080 5788 5132 5840
rect 8392 5788 8444 5840
rect 4160 5720 4212 5772
rect 6276 5720 6328 5772
rect 8208 5720 8260 5772
rect 9036 5856 9088 5908
rect 9496 5856 9548 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 12992 5856 13044 5908
rect 13636 5899 13688 5908
rect 11520 5720 11572 5772
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14648 5856 14700 5908
rect 15016 5856 15068 5908
rect 15292 5856 15344 5908
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 21272 5856 21324 5908
rect 22468 5856 22520 5908
rect 24124 5856 24176 5908
rect 25136 5856 25188 5908
rect 25688 5856 25740 5908
rect 14372 5788 14424 5840
rect 20536 5788 20588 5840
rect 23664 5788 23716 5840
rect 24860 5788 24912 5840
rect 13636 5720 13688 5772
rect 18420 5720 18472 5772
rect 18604 5763 18656 5772
rect 18604 5729 18638 5763
rect 18638 5729 18656 5763
rect 18604 5720 18656 5729
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 22376 5720 22428 5772
rect 22744 5720 22796 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 26148 5720 26200 5772
rect 5080 5652 5132 5704
rect 2780 5516 2832 5568
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 6184 5516 6236 5568
rect 9772 5652 9824 5704
rect 10784 5652 10836 5704
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 14188 5695 14240 5704
rect 14188 5661 14197 5695
rect 14197 5661 14231 5695
rect 14231 5661 14240 5695
rect 14188 5652 14240 5661
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 21364 5695 21416 5704
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 11060 5584 11112 5636
rect 12900 5584 12952 5636
rect 6736 5516 6788 5568
rect 7104 5516 7156 5568
rect 11152 5516 11204 5568
rect 11796 5516 11848 5568
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 23572 5652 23624 5704
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 24952 5652 25004 5704
rect 25412 5584 25464 5636
rect 15568 5516 15620 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 18512 5516 18564 5568
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 23388 5516 23440 5568
rect 23664 5559 23716 5568
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2596 5312 2648 5364
rect 4160 5244 4212 5296
rect 1676 5176 1728 5228
rect 6000 5312 6052 5364
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 7196 5312 7248 5364
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 10784 5355 10836 5364
rect 10784 5321 10793 5355
rect 10793 5321 10827 5355
rect 10827 5321 10836 5355
rect 10784 5312 10836 5321
rect 11980 5312 12032 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 13820 5312 13872 5364
rect 14372 5312 14424 5364
rect 15844 5312 15896 5364
rect 16672 5312 16724 5364
rect 18604 5312 18656 5364
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 21364 5312 21416 5364
rect 22744 5312 22796 5364
rect 23112 5312 23164 5364
rect 24952 5312 25004 5364
rect 25412 5312 25464 5364
rect 25780 5312 25832 5364
rect 6184 5244 6236 5296
rect 6460 5244 6512 5296
rect 2872 5108 2924 5160
rect 7564 5176 7616 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 10140 5244 10192 5296
rect 15292 5244 15344 5296
rect 12256 5176 12308 5228
rect 13636 5176 13688 5228
rect 14188 5176 14240 5228
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 17592 5244 17644 5296
rect 2596 5083 2648 5092
rect 2596 5049 2630 5083
rect 2630 5049 2648 5083
rect 2596 5040 2648 5049
rect 4068 5040 4120 5092
rect 10968 5108 11020 5160
rect 16396 5108 16448 5160
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 22928 5176 22980 5228
rect 5080 5040 5132 5092
rect 9864 5040 9916 5092
rect 11060 5040 11112 5092
rect 11888 5040 11940 5092
rect 13268 5083 13320 5092
rect 13268 5049 13277 5083
rect 13277 5049 13311 5083
rect 13311 5049 13320 5083
rect 13268 5040 13320 5049
rect 17776 5083 17828 5092
rect 17776 5049 17785 5083
rect 17785 5049 17819 5083
rect 17819 5049 17828 5083
rect 17776 5040 17828 5049
rect 19156 5040 19208 5092
rect 20076 5108 20128 5160
rect 21916 5151 21968 5160
rect 21916 5117 21925 5151
rect 21925 5117 21959 5151
rect 21959 5117 21968 5151
rect 21916 5108 21968 5117
rect 23296 5108 23348 5160
rect 23664 5244 23716 5296
rect 25688 5108 25740 5160
rect 1952 4972 2004 5024
rect 2228 4972 2280 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 9588 4972 9640 5024
rect 10968 4972 11020 5024
rect 12072 4972 12124 5024
rect 16120 4972 16172 5024
rect 16396 4972 16448 5024
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 22744 4972 22796 5024
rect 24768 4972 24820 5024
rect 25412 4972 25464 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 5172 4768 5224 4820
rect 6644 4768 6696 4820
rect 7380 4768 7432 4820
rect 9772 4768 9824 4820
rect 10968 4768 11020 4820
rect 12716 4768 12768 4820
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 17868 4768 17920 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 20076 4768 20128 4820
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 1860 4700 1912 4752
rect 664 4632 716 4684
rect 1584 4632 1636 4684
rect 1768 4632 1820 4684
rect 2412 4632 2464 4684
rect 4988 4632 5040 4684
rect 5540 4632 5592 4684
rect 8024 4632 8076 4684
rect 9496 4632 9548 4684
rect 10048 4700 10100 4752
rect 12348 4700 12400 4752
rect 12440 4700 12492 4752
rect 15384 4700 15436 4752
rect 16028 4700 16080 4752
rect 16672 4700 16724 4752
rect 19432 4700 19484 4752
rect 21916 4700 21968 4752
rect 23020 4768 23072 4820
rect 23480 4768 23532 4820
rect 23664 4811 23716 4820
rect 23664 4777 23673 4811
rect 23673 4777 23707 4811
rect 23707 4777 23716 4811
rect 23664 4768 23716 4777
rect 24860 4768 24912 4820
rect 25688 4768 25740 4820
rect 10784 4632 10836 4684
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 16304 4632 16356 4684
rect 17500 4632 17552 4684
rect 17960 4632 18012 4684
rect 19340 4675 19392 4684
rect 19340 4641 19349 4675
rect 19349 4641 19383 4675
rect 19383 4641 19392 4675
rect 19340 4632 19392 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 23204 4632 23256 4684
rect 23480 4632 23532 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 5356 4564 5408 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 18512 4564 18564 4616
rect 19156 4564 19208 4616
rect 21180 4564 21232 4616
rect 20812 4496 20864 4548
rect 22376 4539 22428 4548
rect 22376 4505 22385 4539
rect 22385 4505 22419 4539
rect 22419 4505 22428 4539
rect 24124 4564 24176 4616
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 24860 4564 24912 4616
rect 22376 4496 22428 4505
rect 1952 4428 2004 4480
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 3516 4428 3568 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 6184 4428 6236 4480
rect 6552 4428 6604 4480
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 8668 4471 8720 4480
rect 8668 4437 8677 4471
rect 8677 4437 8711 4471
rect 8711 4437 8720 4471
rect 8668 4428 8720 4437
rect 11796 4471 11848 4480
rect 11796 4437 11805 4471
rect 11805 4437 11839 4471
rect 11839 4437 11848 4471
rect 11796 4428 11848 4437
rect 13636 4471 13688 4480
rect 13636 4437 13645 4471
rect 13645 4437 13679 4471
rect 13679 4437 13688 4471
rect 13636 4428 13688 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15292 4428 15344 4480
rect 16488 4428 16540 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17684 4471 17736 4480
rect 17316 4428 17368 4437
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 18420 4428 18472 4480
rect 19064 4428 19116 4480
rect 20720 4428 20772 4480
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 24032 4471 24084 4480
rect 24032 4437 24041 4471
rect 24041 4437 24075 4471
rect 24075 4437 24084 4471
rect 24032 4428 24084 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1492 4267 1544 4276
rect 1492 4233 1501 4267
rect 1501 4233 1535 4267
rect 1535 4233 1544 4267
rect 1492 4224 1544 4233
rect 1768 4224 1820 4276
rect 3056 4224 3108 4276
rect 4160 4224 4212 4276
rect 4988 4267 5040 4276
rect 4988 4233 4997 4267
rect 4997 4233 5031 4267
rect 5031 4233 5040 4267
rect 4988 4224 5040 4233
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 6000 4224 6052 4276
rect 5540 4156 5592 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2596 4088 2648 4140
rect 6276 4088 6328 4140
rect 7748 4224 7800 4276
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 10784 4224 10836 4276
rect 10968 4224 11020 4276
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 15660 4267 15712 4276
rect 15660 4233 15669 4267
rect 15669 4233 15703 4267
rect 15703 4233 15712 4267
rect 15660 4224 15712 4233
rect 23020 4224 23072 4276
rect 23480 4267 23532 4276
rect 23480 4233 23489 4267
rect 23489 4233 23523 4267
rect 23523 4233 23532 4267
rect 23480 4224 23532 4233
rect 24124 4224 24176 4276
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 2872 4020 2924 4072
rect 3332 4020 3384 4072
rect 4068 4020 4120 4072
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 6368 4020 6420 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8024 4020 8076 4072
rect 8668 4020 8720 4072
rect 9588 4020 9640 4072
rect 3516 3995 3568 4004
rect 3516 3961 3550 3995
rect 3550 3961 3568 3995
rect 3516 3952 3568 3961
rect 9036 3952 9088 4004
rect 10784 4020 10836 4072
rect 12348 4020 12400 4072
rect 12716 4020 12768 4072
rect 2412 3884 2464 3936
rect 6920 3884 6972 3936
rect 8668 3884 8720 3936
rect 9220 3884 9272 3936
rect 10692 3952 10744 4004
rect 13636 4088 13688 4140
rect 19156 4199 19208 4208
rect 19156 4165 19165 4199
rect 19165 4165 19199 4199
rect 19199 4165 19208 4199
rect 19156 4156 19208 4165
rect 16488 4088 16540 4140
rect 17040 4088 17092 4140
rect 17868 4088 17920 4140
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 20260 4156 20312 4208
rect 14280 4020 14332 4072
rect 15292 4020 15344 4072
rect 16764 4020 16816 4072
rect 12992 3952 13044 4004
rect 16120 3952 16172 4004
rect 16948 3952 17000 4004
rect 18236 4020 18288 4072
rect 18788 4020 18840 4072
rect 20168 4088 20220 4140
rect 20444 4088 20496 4140
rect 20812 4088 20864 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 23112 4088 23164 4140
rect 24860 4088 24912 4140
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 25688 4088 25740 4140
rect 23664 4020 23716 4072
rect 24308 4020 24360 4072
rect 25596 4020 25648 4072
rect 22008 3952 22060 4004
rect 9864 3884 9916 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12716 3884 12768 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 23296 3952 23348 4004
rect 23204 3884 23256 3936
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1860 3680 1912 3732
rect 2596 3723 2648 3732
rect 2596 3689 2605 3723
rect 2605 3689 2639 3723
rect 2639 3689 2648 3723
rect 2596 3680 2648 3689
rect 3884 3680 3936 3732
rect 4436 3680 4488 3732
rect 5540 3680 5592 3732
rect 7748 3680 7800 3732
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 10692 3680 10744 3732
rect 10968 3680 11020 3732
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 12440 3680 12492 3732
rect 1676 3612 1728 3664
rect 2504 3612 2556 3664
rect 5448 3655 5500 3664
rect 5448 3621 5457 3655
rect 5457 3621 5491 3655
rect 5491 3621 5500 3655
rect 5448 3612 5500 3621
rect 6000 3655 6052 3664
rect 6000 3621 6034 3655
rect 6034 3621 6052 3655
rect 6000 3612 6052 3621
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 1400 3544 1452 3596
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5264 3544 5316 3596
rect 6736 3544 6788 3596
rect 2228 3476 2280 3528
rect 3976 3476 4028 3528
rect 5356 3476 5408 3528
rect 2964 3451 3016 3460
rect 2964 3417 2973 3451
rect 2973 3417 3007 3451
rect 3007 3417 3016 3451
rect 2964 3408 3016 3417
rect 3516 3408 3568 3460
rect 3792 3408 3844 3460
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8760 3544 8812 3596
rect 10048 3612 10100 3664
rect 12256 3612 12308 3664
rect 12348 3612 12400 3664
rect 14004 3680 14056 3732
rect 15292 3680 15344 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 16120 3680 16172 3732
rect 18236 3680 18288 3732
rect 18604 3680 18656 3732
rect 19984 3680 20036 3732
rect 20628 3680 20680 3732
rect 21180 3723 21232 3732
rect 21180 3689 21189 3723
rect 21189 3689 21223 3723
rect 21223 3689 21232 3723
rect 21180 3680 21232 3689
rect 21272 3680 21324 3732
rect 21548 3680 21600 3732
rect 13452 3655 13504 3664
rect 13452 3621 13461 3655
rect 13461 3621 13495 3655
rect 13495 3621 13504 3655
rect 13452 3612 13504 3621
rect 15384 3612 15436 3664
rect 16304 3612 16356 3664
rect 17500 3612 17552 3664
rect 18880 3655 18932 3664
rect 18880 3621 18889 3655
rect 18889 3621 18923 3655
rect 18923 3621 18932 3655
rect 18880 3612 18932 3621
rect 25596 3680 25648 3732
rect 22192 3612 22244 3664
rect 22652 3612 22704 3664
rect 23480 3612 23532 3664
rect 25688 3612 25740 3664
rect 9956 3587 10008 3596
rect 9956 3553 9990 3587
rect 9990 3553 10008 3587
rect 9956 3544 10008 3553
rect 13820 3544 13872 3596
rect 8024 3476 8076 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 11888 3476 11940 3528
rect 12716 3476 12768 3528
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 13636 3476 13688 3528
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 17776 3544 17828 3596
rect 16028 3476 16080 3485
rect 18236 3476 18288 3528
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 7840 3451 7892 3460
rect 7840 3417 7849 3451
rect 7849 3417 7883 3451
rect 7883 3417 7892 3451
rect 7840 3408 7892 3417
rect 12532 3408 12584 3460
rect 15292 3408 15344 3460
rect 18144 3408 18196 3460
rect 8576 3340 8628 3392
rect 12900 3340 12952 3392
rect 13728 3340 13780 3392
rect 13912 3383 13964 3392
rect 13912 3349 13921 3383
rect 13921 3349 13955 3383
rect 13955 3349 13964 3383
rect 13912 3340 13964 3349
rect 14188 3383 14240 3392
rect 14188 3349 14197 3383
rect 14197 3349 14231 3383
rect 14231 3349 14240 3383
rect 14188 3340 14240 3349
rect 16764 3340 16816 3392
rect 17040 3383 17092 3392
rect 17040 3349 17049 3383
rect 17049 3349 17083 3383
rect 17083 3349 17092 3383
rect 17040 3340 17092 3349
rect 20996 3544 21048 3596
rect 23664 3544 23716 3596
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 23112 3408 23164 3460
rect 20536 3340 20588 3392
rect 20720 3383 20772 3392
rect 20720 3349 20729 3383
rect 20729 3349 20763 3383
rect 20763 3349 20772 3383
rect 20720 3340 20772 3349
rect 22744 3340 22796 3392
rect 24124 3340 24176 3392
rect 24768 3340 24820 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 5264 3179 5316 3188
rect 3056 3136 3108 3145
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6000 3136 6052 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 9956 3136 10008 3188
rect 10784 3136 10836 3188
rect 3424 3111 3476 3120
rect 3424 3077 3433 3111
rect 3433 3077 3467 3111
rect 3467 3077 3476 3111
rect 3424 3068 3476 3077
rect 2320 2932 2372 2984
rect 3332 3000 3384 3052
rect 8024 3111 8076 3120
rect 8024 3077 8033 3111
rect 8033 3077 8067 3111
rect 8067 3077 8076 3111
rect 8024 3068 8076 3077
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 3056 2932 3108 2984
rect 7104 2932 7156 2984
rect 11244 3136 11296 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 13084 3136 13136 3188
rect 15844 3136 15896 3188
rect 11336 3043 11388 3052
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 13820 3000 13872 3052
rect 14464 3000 14516 3052
rect 12256 2932 12308 2984
rect 12716 2975 12768 2984
rect 12716 2941 12750 2975
rect 12750 2941 12768 2975
rect 12716 2932 12768 2941
rect 14740 2932 14792 2984
rect 16856 3136 16908 3188
rect 17776 3136 17828 3188
rect 18236 3136 18288 3188
rect 18604 3136 18656 3188
rect 19892 3136 19944 3188
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 22192 3136 22244 3188
rect 22744 3179 22796 3188
rect 22744 3145 22753 3179
rect 22753 3145 22787 3179
rect 22787 3145 22796 3179
rect 22744 3136 22796 3145
rect 23664 3136 23716 3188
rect 24676 3136 24728 3188
rect 24952 3136 25004 3188
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 20444 3111 20496 3120
rect 20444 3077 20453 3111
rect 20453 3077 20487 3111
rect 20487 3077 20496 3111
rect 20444 3068 20496 3077
rect 25596 3068 25648 3120
rect 26056 3111 26108 3120
rect 26056 3077 26065 3111
rect 26065 3077 26099 3111
rect 26099 3077 26108 3111
rect 26056 3068 26108 3077
rect 16764 3000 16816 3052
rect 18236 3000 18288 3052
rect 19064 2932 19116 2984
rect 23112 3000 23164 3052
rect 20904 2975 20956 2984
rect 20904 2941 20927 2975
rect 20927 2941 20956 2975
rect 3976 2864 4028 2916
rect 8852 2864 8904 2916
rect 13912 2864 13964 2916
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 16580 2907 16632 2916
rect 16580 2873 16589 2907
rect 16589 2873 16623 2907
rect 16623 2873 16632 2907
rect 16580 2864 16632 2873
rect 18880 2864 18932 2916
rect 20904 2932 20956 2941
rect 20996 2864 21048 2916
rect 25596 2864 25648 2916
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 3516 2796 3568 2848
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 12992 2796 13044 2848
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 17500 2796 17552 2848
rect 20352 2796 20404 2848
rect 25228 2796 25280 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1400 2635 1452 2644
rect 1400 2601 1409 2635
rect 1409 2601 1443 2635
rect 1443 2601 1452 2635
rect 1400 2592 1452 2601
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 2320 2592 2372 2644
rect 3792 2592 3844 2644
rect 3424 2567 3476 2576
rect 3424 2533 3433 2567
rect 3433 2533 3467 2567
rect 3467 2533 3476 2567
rect 3424 2524 3476 2533
rect 4528 2524 4580 2576
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 5356 2592 5408 2644
rect 6460 2592 6512 2644
rect 6828 2592 6880 2644
rect 7288 2592 7340 2644
rect 9680 2592 9732 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 12348 2592 12400 2644
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 17960 2592 18012 2644
rect 18144 2592 18196 2644
rect 8024 2456 8076 2508
rect 8208 2499 8260 2508
rect 8208 2465 8217 2499
rect 8217 2465 8251 2499
rect 8251 2465 8260 2499
rect 8208 2456 8260 2465
rect 6920 2388 6972 2440
rect 8484 2388 8536 2440
rect 12992 2524 13044 2576
rect 14464 2524 14516 2576
rect 11520 2456 11572 2508
rect 10692 2388 10744 2440
rect 12256 2388 12308 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 15292 2524 15344 2576
rect 19984 2592 20036 2644
rect 20536 2592 20588 2644
rect 22468 2592 22520 2644
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 24952 2592 25004 2644
rect 25596 2635 25648 2644
rect 25596 2601 25605 2635
rect 25605 2601 25639 2635
rect 25639 2601 25648 2635
rect 25596 2592 25648 2601
rect 20904 2567 20956 2576
rect 20904 2533 20913 2567
rect 20913 2533 20947 2567
rect 20947 2533 20956 2567
rect 20904 2524 20956 2533
rect 26056 2524 26108 2576
rect 16304 2456 16356 2508
rect 16856 2456 16908 2508
rect 18052 2499 18104 2508
rect 18052 2465 18061 2499
rect 18061 2465 18095 2499
rect 18095 2465 18104 2499
rect 18052 2456 18104 2465
rect 18144 2456 18196 2508
rect 20536 2499 20588 2508
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 23756 2456 23808 2508
rect 10876 2363 10928 2372
rect 10876 2329 10885 2363
rect 10885 2329 10919 2363
rect 10919 2329 10928 2363
rect 10876 2320 10928 2329
rect 15476 2363 15528 2372
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 16672 2320 16724 2372
rect 18236 2320 18288 2372
rect 23480 2363 23532 2372
rect 23480 2329 23489 2363
rect 23489 2329 23523 2363
rect 23523 2329 23532 2363
rect 24952 2388 25004 2440
rect 23480 2320 23532 2329
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 4528 2252 4580 2304
rect 4712 2252 4764 2304
rect 6184 2252 6236 2304
rect 8852 2295 8904 2304
rect 8852 2261 8861 2295
rect 8861 2261 8895 2295
rect 8895 2261 8904 2295
rect 8852 2252 8904 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 14004 2295 14056 2304
rect 14004 2261 14013 2295
rect 14013 2261 14047 2295
rect 14047 2261 14056 2295
rect 14004 2252 14056 2261
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 22560 2295 22612 2304
rect 22560 2261 22569 2295
rect 22569 2261 22603 2295
rect 22603 2261 22612 2295
rect 22560 2252 22612 2261
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 12624 2048 12676 2100
rect 17684 2048 17736 2100
rect 3056 1368 3108 1420
rect 8392 1368 8444 1420
rect 4896 552 4948 604
rect 5264 552 5316 604
rect 12164 552 12216 604
rect 12532 552 12584 604
<< metal2 >>
rect 3422 27704 3478 27713
rect 3422 27639 3478 27648
rect 2686 26616 2742 26625
rect 2686 26551 2742 26560
rect 1582 24304 1638 24313
rect 1582 24239 1638 24248
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1504 21690 1532 23151
rect 1596 22778 1624 24239
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 2594 22536 2650 22545
rect 2594 22471 2650 22480
rect 2044 22432 2096 22438
rect 2042 22400 2044 22409
rect 2096 22400 2098 22409
rect 2042 22335 2098 22344
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1490 21448 1546 21457
rect 1490 21383 1546 21392
rect 1504 20602 1532 21383
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 2056 21078 2084 21286
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 1582 20904 1638 20913
rect 1582 20839 1638 20848
rect 1492 20596 1544 20602
rect 1492 20538 1544 20544
rect 1490 20360 1546 20369
rect 1490 20295 1546 20304
rect 1398 19680 1454 19689
rect 1398 19615 1454 19624
rect 1412 18426 1440 19615
rect 1504 19174 1532 20295
rect 1596 20058 1624 20839
rect 2332 20262 2360 20946
rect 2044 20256 2096 20262
rect 2042 20224 2044 20233
rect 2320 20256 2372 20262
rect 2096 20224 2098 20233
rect 2320 20198 2372 20204
rect 2042 20159 2098 20168
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1596 18986 1624 19246
rect 1504 18958 1624 18986
rect 2332 18986 2360 20198
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2424 19174 2452 19858
rect 2412 19168 2464 19174
rect 2410 19136 2412 19145
rect 2464 19136 2466 19145
rect 2410 19071 2466 19080
rect 2332 18958 2452 18986
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1504 18306 1532 18958
rect 1584 18624 1636 18630
rect 1582 18592 1584 18601
rect 1768 18624 1820 18630
rect 1636 18592 1638 18601
rect 1768 18566 1820 18572
rect 1582 18527 1638 18536
rect 1412 18278 1532 18306
rect 1412 16402 1440 18278
rect 1780 17746 1808 18566
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1492 17740 1544 17746
rect 1492 17682 1544 17688
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1320 16374 1440 16402
rect 1320 15366 1348 16374
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 1412 14498 1440 16186
rect 1320 14470 1440 14498
rect 1216 13184 1268 13190
rect 1216 13126 1268 13132
rect 1228 11218 1256 13126
rect 1320 12322 1348 14470
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 12442 1440 14350
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1320 12294 1440 12322
rect 1216 11212 1268 11218
rect 1216 11154 1268 11160
rect 1412 9081 1440 12294
rect 1504 11354 1532 17682
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1596 16794 1624 16934
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1596 16114 1624 16730
rect 1688 16658 1716 16934
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1688 13954 1716 16594
rect 1768 15904 1820 15910
rect 1820 15852 1900 15858
rect 1768 15846 1900 15852
rect 1780 15830 1900 15846
rect 1872 15473 1900 15830
rect 1964 15688 1992 18022
rect 2332 17814 2360 18022
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 17202 2084 17478
rect 2148 17202 2176 17614
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2044 16584 2096 16590
rect 2042 16552 2044 16561
rect 2148 16572 2176 17138
rect 2096 16552 2176 16572
rect 2098 16544 2176 16552
rect 2042 16487 2098 16496
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 1964 15660 2084 15688
rect 1952 15496 2004 15502
rect 1858 15464 1914 15473
rect 1768 15428 1820 15434
rect 1952 15438 2004 15444
rect 1858 15399 1914 15408
rect 1768 15370 1820 15376
rect 1780 14958 1808 15370
rect 1872 15026 1900 15399
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1964 14278 1992 15438
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1596 13926 1716 13954
rect 1596 11558 1624 13926
rect 1860 13864 1912 13870
rect 1964 13841 1992 14214
rect 1860 13806 1912 13812
rect 1950 13832 2006 13841
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1688 13530 1716 13738
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1688 12850 1716 13466
rect 1872 13394 1900 13806
rect 1950 13767 2006 13776
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1766 11656 1822 11665
rect 1766 11591 1822 11600
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1582 11384 1638 11393
rect 1492 11348 1544 11354
rect 1582 11319 1638 11328
rect 1492 11290 1544 11296
rect 1596 11286 1624 11319
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1504 7585 1532 11154
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 664 4684 716 4690
rect 664 4626 716 4632
rect 676 3233 704 4626
rect 1412 3602 1440 7142
rect 1492 6928 1544 6934
rect 1492 6870 1544 6876
rect 1504 4282 1532 6870
rect 1596 4690 1624 7686
rect 1688 5778 1716 8366
rect 1780 6730 1808 11591
rect 1872 11082 1900 13330
rect 1950 13288 2006 13297
rect 1950 13223 2006 13232
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10674 1900 11018
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 10198 1900 10610
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1964 9654 1992 13223
rect 2056 13190 2084 15660
rect 2148 15570 2176 16390
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 2056 12374 2084 12854
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11830 2084 12310
rect 2148 12102 2176 14758
rect 2240 14113 2268 17478
rect 2320 15632 2372 15638
rect 2424 15609 2452 18958
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2516 16250 2544 16594
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2320 15574 2372 15580
rect 2410 15600 2466 15609
rect 2332 15450 2360 15574
rect 2410 15535 2466 15544
rect 2516 15502 2544 16050
rect 2504 15496 2556 15502
rect 2332 15422 2452 15450
rect 2504 15438 2556 15444
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2226 14104 2282 14113
rect 2226 14039 2282 14048
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2240 13462 2268 13670
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2240 12918 2268 13398
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2332 12753 2360 15302
rect 2424 14822 2452 15422
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2318 12744 2374 12753
rect 2318 12679 2374 12688
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2240 12209 2268 12582
rect 2332 12481 2360 12582
rect 2318 12472 2374 12481
rect 2318 12407 2374 12416
rect 2226 12200 2282 12209
rect 2226 12135 2228 12144
rect 2280 12135 2282 12144
rect 2228 12106 2280 12112
rect 2136 12096 2188 12102
rect 2240 12075 2268 12106
rect 2136 12038 2188 12044
rect 2226 11928 2282 11937
rect 2332 11898 2360 12407
rect 2424 12186 2452 14758
rect 2516 12306 2544 15302
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2424 12158 2544 12186
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2226 11863 2282 11872
rect 2320 11892 2372 11898
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 2240 11762 2268 11863
rect 2320 11834 2372 11840
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2134 11520 2190 11529
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 2056 9466 2084 11494
rect 2134 11455 2190 11464
rect 2148 9586 2176 11455
rect 2240 11393 2268 11698
rect 2226 11384 2282 11393
rect 2226 11319 2282 11328
rect 2332 11286 2360 11698
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2424 11218 2452 12038
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10810 2268 11086
rect 2410 10976 2466 10985
rect 2410 10911 2466 10920
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1872 9438 2084 9466
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1688 5234 1716 5714
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1872 4758 1900 9438
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9042 2084 9318
rect 2148 9178 2176 9522
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2148 8430 2176 9114
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 8090 2176 8366
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1964 5030 1992 5714
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1860 4752 1912 4758
rect 1860 4694 1912 4700
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1674 4312 1730 4321
rect 1492 4276 1544 4282
rect 1780 4282 1808 4626
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1674 4247 1730 4256
rect 1768 4276 1820 4282
rect 1492 4218 1544 4224
rect 1582 3768 1638 3777
rect 1504 3726 1582 3754
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 662 3224 718 3233
rect 662 3159 718 3168
rect 846 3224 902 3233
rect 846 3159 902 3168
rect 294 1728 350 1737
rect 294 1663 350 1672
rect 308 480 336 1663
rect 860 480 888 3159
rect 1398 2680 1454 2689
rect 1398 2615 1400 2624
rect 1452 2615 1454 2624
rect 1400 2586 1452 2592
rect 1504 1850 1532 3726
rect 1582 3703 1638 3712
rect 1688 3670 1716 4247
rect 1768 4218 1820 4224
rect 1858 4176 1914 4185
rect 1964 4146 1992 4422
rect 1858 4111 1914 4120
rect 1952 4140 2004 4146
rect 1872 4078 1900 4111
rect 1952 4082 2004 4088
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1872 3738 1900 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1688 3194 1716 3606
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1872 2650 1900 3538
rect 2056 3194 2084 7958
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 6798 2176 7142
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6633 2176 6734
rect 2134 6624 2190 6633
rect 2134 6559 2190 6568
rect 2240 5273 2268 7822
rect 2332 6458 2360 9862
rect 2424 9178 2452 10911
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2516 9110 2544 12158
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2410 7848 2466 7857
rect 2410 7783 2412 7792
rect 2464 7783 2466 7792
rect 2504 7812 2556 7818
rect 2412 7754 2464 7760
rect 2504 7754 2556 7760
rect 2516 7478 2544 7754
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2608 6882 2636 22471
rect 2700 18970 2728 26551
rect 3436 24562 3464 27639
rect 3514 27520 3570 28000
rect 10506 27520 10562 28000
rect 17498 27520 17554 28000
rect 24214 27704 24270 27713
rect 24214 27639 24270 27648
rect 3528 24721 3556 27520
rect 4066 27160 4122 27169
rect 4122 27118 4200 27146
rect 4066 27095 4122 27104
rect 3698 26072 3754 26081
rect 3698 26007 3700 26016
rect 3752 26007 3754 26016
rect 3700 25978 3752 25984
rect 4066 25392 4122 25401
rect 4066 25327 4122 25336
rect 4080 25158 4108 25327
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 3514 24712 3570 24721
rect 3514 24647 3570 24656
rect 3436 24534 3556 24562
rect 2778 23760 2834 23769
rect 2778 23695 2834 23704
rect 2792 23089 2820 23695
rect 2778 23080 2834 23089
rect 2778 23015 2834 23024
rect 2870 19000 2926 19009
rect 2688 18964 2740 18970
rect 2870 18935 2926 18944
rect 2688 18906 2740 18912
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2700 17082 2728 17682
rect 2792 17513 2820 18022
rect 2884 17882 2912 18935
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 2976 17202 3004 18566
rect 3160 18086 3188 18770
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3148 17128 3200 17134
rect 2778 17096 2834 17105
rect 2700 17054 2778 17082
rect 3148 17070 3200 17076
rect 2778 17031 2780 17040
rect 2832 17031 2834 17040
rect 2780 17002 2832 17008
rect 2792 16971 2820 17002
rect 3160 16697 3188 17070
rect 2686 16688 2742 16697
rect 3146 16688 3202 16697
rect 2686 16623 2742 16632
rect 2780 16652 2832 16658
rect 2700 14618 2728 16623
rect 3146 16623 3202 16632
rect 2780 16594 2832 16600
rect 2792 15706 2820 16594
rect 2870 16552 2926 16561
rect 2870 16487 2872 16496
rect 2924 16487 2926 16496
rect 2872 16458 2924 16464
rect 2884 16114 2912 16458
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2870 15736 2926 15745
rect 2780 15700 2832 15706
rect 2870 15671 2926 15680
rect 2780 15642 2832 15648
rect 2792 15366 2820 15642
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2884 14906 2912 15671
rect 2976 15366 3004 15982
rect 3056 15904 3108 15910
rect 3252 15892 3280 16118
rect 3332 15904 3384 15910
rect 3252 15864 3332 15892
rect 3056 15846 3108 15852
rect 3332 15846 3384 15852
rect 3068 15706 3096 15846
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2792 14878 2912 14906
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2700 12986 2728 14418
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2792 12714 2820 14878
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2884 12594 2912 14758
rect 2976 13025 3004 15302
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 14074 3096 14350
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3054 13832 3110 13841
rect 3054 13767 3110 13776
rect 2962 13016 3018 13025
rect 2962 12951 3018 12960
rect 2792 12566 2912 12594
rect 2792 11370 2820 12566
rect 3068 12458 3096 13767
rect 3160 13530 3188 15506
rect 3238 14920 3294 14929
rect 3238 14855 3294 14864
rect 3252 13977 3280 14855
rect 3238 13968 3294 13977
rect 3238 13903 3294 13912
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 12782 3280 13126
rect 3240 12776 3292 12782
rect 3146 12744 3202 12753
rect 3240 12718 3292 12724
rect 3146 12679 3202 12688
rect 2976 12430 3096 12458
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 11558 2912 12242
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2700 11354 2820 11370
rect 2688 11348 2820 11354
rect 2740 11342 2820 11348
rect 2688 11290 2740 11296
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 10266 2728 10474
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2792 10198 2820 11342
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2884 9874 2912 11494
rect 2976 10130 3004 12430
rect 3054 12064 3110 12073
rect 3054 11999 3110 12008
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2792 9846 2912 9874
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 6934 2728 8842
rect 2516 6854 2636 6882
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2516 6186 2544 6854
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2608 6118 2636 6734
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5370 2636 6054
rect 2792 5794 2820 9846
rect 2976 9518 3004 10066
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2872 9376 2924 9382
rect 2870 9344 2872 9353
rect 2924 9344 2926 9353
rect 2870 9279 2926 9288
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2976 8634 3004 9454
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 7546 2912 7822
rect 3068 7750 3096 11999
rect 3160 11354 3188 12679
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3146 10160 3202 10169
rect 3146 10095 3202 10104
rect 3160 9926 3188 10095
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3160 9382 3188 9415
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3160 8362 3188 8978
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7546 3096 7686
rect 2872 7540 2924 7546
rect 3056 7540 3108 7546
rect 2924 7500 3004 7528
rect 2872 7482 2924 7488
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2884 6118 2912 7278
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5914 2912 6054
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2700 5766 2820 5794
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2226 5264 2282 5273
rect 2700 5250 2728 5766
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2226 5199 2282 5208
rect 2516 5222 2728 5250
rect 2228 5024 2280 5030
rect 2134 4992 2190 5001
rect 2228 4966 2280 4972
rect 2134 4927 2190 4936
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2148 2530 2176 4927
rect 2240 4622 2268 4966
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2318 4584 2374 4593
rect 2240 3534 2268 4558
rect 2318 4519 2374 4528
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 2650 2268 3470
rect 2332 2990 2360 4519
rect 2424 3942 2452 4626
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 2650 2360 2926
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 1412 1822 1532 1850
rect 1964 2502 2176 2530
rect 1412 480 1440 1822
rect 1964 480 1992 2502
rect 2424 2009 2452 3878
rect 2516 3670 2544 5222
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2608 4808 2636 5034
rect 2792 4808 2820 5510
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2608 4780 2820 4808
rect 2608 4486 2636 4780
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2608 4146 2636 4422
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 3738 2636 4082
rect 2884 4078 2912 5102
rect 2872 4072 2924 4078
rect 2976 4049 3004 7500
rect 3056 7482 3108 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 5574 3096 7346
rect 3160 6118 3188 8298
rect 3148 6112 3200 6118
rect 3252 6089 3280 12582
rect 3344 9897 3372 15846
rect 3436 14618 3464 17478
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3436 12986 3464 14554
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 10538 3464 12786
rect 3528 11937 3556 24534
rect 3974 21992 4030 22001
rect 3974 21927 4030 21936
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17134 3648 17478
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3896 15706 3924 18022
rect 3988 16561 4016 21927
rect 4172 17882 4200 27118
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5552 23866 5580 25094
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 7838 24848 7894 24857
rect 7838 24783 7894 24792
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 4710 22400 4766 22409
rect 4710 22335 4766 22344
rect 4342 19136 4398 19145
rect 4342 19071 4398 19080
rect 4356 18902 4384 19071
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4448 18086 4476 18770
rect 4436 18080 4488 18086
rect 4250 18048 4306 18057
rect 4436 18022 4488 18028
rect 4250 17983 4306 17992
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3974 16552 4030 16561
rect 3974 16487 4030 16496
rect 4080 16289 4108 16730
rect 4264 16658 4292 17983
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4356 16998 4384 17682
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4066 16280 4122 16289
rect 4066 16215 4122 16224
rect 4172 16046 4200 16526
rect 4160 16040 4212 16046
rect 4158 16008 4160 16017
rect 4212 16008 4214 16017
rect 4158 15943 4214 15952
rect 4356 15881 4384 16934
rect 4342 15872 4398 15881
rect 4342 15807 4398 15816
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3620 14278 3648 14962
rect 3712 14278 3740 15506
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 14958 4108 15302
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3620 12850 3648 14214
rect 3712 13297 3740 14214
rect 3896 13841 3924 14758
rect 3974 14648 4030 14657
rect 3974 14583 4030 14592
rect 3988 13977 4016 14583
rect 3974 13968 4030 13977
rect 3974 13903 4030 13912
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3882 13696 3938 13705
rect 3882 13631 3938 13640
rect 3698 13288 3754 13297
rect 3698 13223 3754 13232
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3606 12744 3662 12753
rect 3606 12679 3662 12688
rect 3514 11928 3570 11937
rect 3514 11863 3570 11872
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3528 10130 3556 11863
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3330 9888 3386 9897
rect 3330 9823 3386 9832
rect 3528 9636 3556 10066
rect 3330 9616 3386 9625
rect 3330 9551 3386 9560
rect 3436 9608 3556 9636
rect 3344 8022 3372 9551
rect 3436 9382 3464 9608
rect 3620 9489 3648 12679
rect 3790 11792 3846 11801
rect 3790 11727 3846 11736
rect 3804 10713 3832 11727
rect 3896 11694 3924 13631
rect 4080 13530 4108 14894
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4172 12968 4200 14282
rect 4264 14278 4292 15438
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4080 12940 4200 12968
rect 4080 12850 4108 12940
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12640 4028 12646
rect 3974 12608 3976 12617
rect 4028 12608 4030 12617
rect 3974 12543 4030 12552
rect 4172 12345 4200 12940
rect 4158 12336 4214 12345
rect 4158 12271 4214 12280
rect 4264 12220 4292 14214
rect 4356 12753 4384 14894
rect 4342 12744 4398 12753
rect 4342 12679 4398 12688
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4172 12192 4292 12220
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11762 4016 12038
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 11393 3924 11494
rect 3882 11384 3938 11393
rect 4080 11336 4108 11766
rect 4172 11540 4200 12192
rect 4356 11830 4384 12242
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4172 11512 4292 11540
rect 3882 11319 3884 11328
rect 3936 11319 3938 11328
rect 3884 11290 3936 11296
rect 3988 11308 4108 11336
rect 3882 11248 3938 11257
rect 3882 11183 3884 11192
rect 3936 11183 3938 11192
rect 3884 11154 3936 11160
rect 3988 10742 4016 11308
rect 4160 11280 4212 11286
rect 4080 11240 4160 11268
rect 4080 10810 4108 11240
rect 4160 11222 4212 11228
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3976 10736 4028 10742
rect 3790 10704 3846 10713
rect 3976 10678 4028 10684
rect 3790 10639 3846 10648
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3804 9625 3832 10231
rect 3790 9616 3846 9625
rect 3790 9551 3846 9560
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3148 6054 3200 6060
rect 3238 6080 3294 6089
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2872 4014 2924 4020
rect 2962 4040 3018 4049
rect 2962 3975 3018 3984
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2504 2848 2556 2854
rect 2502 2816 2504 2825
rect 2556 2816 2558 2825
rect 2502 2751 2558 2760
rect 2410 2000 2466 2009
rect 2410 1935 2466 1944
rect 2608 1442 2636 3023
rect 2516 1414 2636 1442
rect 2516 480 2544 1414
rect 2884 921 2912 3567
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2976 2446 3004 3402
rect 3068 3194 3096 4218
rect 3160 3641 3188 6054
rect 3238 6015 3294 6024
rect 3344 5953 3372 7142
rect 3436 7002 3464 9318
rect 3620 9217 3648 9318
rect 3606 9208 3662 9217
rect 3606 9143 3662 9152
rect 3804 8265 3832 9415
rect 3896 8838 3924 9522
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3790 8256 3846 8265
rect 3790 8191 3846 8200
rect 3514 7984 3570 7993
rect 3514 7919 3516 7928
rect 3568 7919 3570 7928
rect 3516 7890 3568 7896
rect 3424 6996 3476 7002
rect 3476 6956 3556 6984
rect 3424 6938 3476 6944
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6322 3464 6598
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 6089 3464 6258
rect 3528 6254 3556 6956
rect 3896 6662 3924 8774
rect 3988 8090 4016 8910
rect 4080 8650 4108 10367
rect 4080 8622 4200 8650
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3988 7585 4016 7822
rect 3974 7576 4030 7585
rect 3974 7511 3976 7520
rect 4028 7511 4030 7520
rect 3976 7482 4028 7488
rect 4080 6984 4108 8502
rect 4172 7970 4200 8622
rect 4264 8090 4292 11512
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4172 7942 4292 7970
rect 3988 6956 4200 6984
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3422 6080 3478 6089
rect 3422 6015 3478 6024
rect 3330 5944 3386 5953
rect 3330 5879 3386 5888
rect 3344 5846 3372 5879
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3436 5778 3464 6015
rect 3896 5914 3924 6598
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3606 5808 3662 5817
rect 3424 5772 3476 5778
rect 3988 5794 4016 6956
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 4172 6798 4200 6956
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4264 6610 4292 7942
rect 4356 7274 4384 11630
rect 4448 11354 4476 18022
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4632 16833 4660 16934
rect 4618 16824 4674 16833
rect 4618 16759 4674 16768
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15337 4568 15846
rect 4526 15328 4582 15337
rect 4526 15263 4582 15272
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14618 4568 14758
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4632 14482 4660 16594
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 11898 4568 14350
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12374 4660 13330
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4540 11694 4568 11727
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4632 11200 4660 12310
rect 4724 11937 4752 22335
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5354 20224 5410 20233
rect 5354 20159 5410 20168
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 5262 17096 5318 17105
rect 4816 16114 4844 17070
rect 5262 17031 5318 17040
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4816 15026 4844 15438
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5000 14958 5028 15302
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4710 11928 4766 11937
rect 4710 11863 4766 11872
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4448 11172 4660 11200
rect 4448 11014 4476 11172
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4448 10674 4476 10950
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4448 10130 4476 10610
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4540 9654 4568 11018
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 10266 4660 10542
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4618 9888 4674 9897
rect 4618 9823 4674 9832
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4526 9072 4582 9081
rect 4526 9007 4528 9016
rect 4580 9007 4582 9016
rect 4528 8978 4580 8984
rect 4540 8566 4568 8978
rect 4632 8634 4660 9823
rect 4724 9110 4752 11766
rect 4816 10985 4844 14758
rect 4894 14104 4950 14113
rect 4894 14039 4950 14048
rect 4908 13954 4936 14039
rect 4908 13926 5028 13954
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4908 13394 4936 13738
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5000 13274 5028 13926
rect 5184 13410 5212 15642
rect 4908 13246 5028 13274
rect 5092 13382 5212 13410
rect 4908 11830 4936 13246
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11286 4936 11494
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4802 10976 4858 10985
rect 4802 10911 4858 10920
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 10266 4936 10746
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4540 8072 4568 8502
rect 4632 8362 4660 8570
rect 4724 8430 4752 9046
rect 4816 8838 4844 9862
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4448 8044 4568 8072
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 3606 5743 3662 5752
rect 3712 5766 4016 5794
rect 4080 6582 4292 6610
rect 3424 5714 3476 5720
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3146 3632 3202 3641
rect 3146 3567 3202 3576
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3068 2990 3096 3130
rect 3344 3058 3372 4014
rect 3528 4010 3556 4422
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3422 3496 3478 3505
rect 3528 3466 3556 3946
rect 3422 3431 3478 3440
rect 3516 3460 3568 3466
rect 3436 3126 3464 3431
rect 3516 3402 3568 3408
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3528 2854 3556 3402
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3424 2576 3476 2582
rect 3422 2544 3424 2553
rect 3476 2544 3478 2553
rect 3422 2479 3478 2488
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3056 1420 3108 1426
rect 3056 1362 3108 1368
rect 2870 912 2926 921
rect 2870 847 2926 856
rect 3068 480 3096 1362
rect 3620 480 3648 5743
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 3712 377 3740 5766
rect 4080 5658 4108 6582
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3988 5630 4108 5658
rect 3988 4865 4016 5630
rect 4172 5302 4200 5714
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3974 4856 4030 4865
rect 3974 4791 4030 4800
rect 4080 4078 4108 5034
rect 4172 4282 4200 5238
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4264 4185 4292 4422
rect 4250 4176 4306 4185
rect 4250 4111 4306 4120
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4448 3738 4476 8044
rect 4632 7970 4660 8298
rect 4540 7942 4660 7970
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 3896 3505 3924 3674
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 3976 3528 4028 3534
rect 3882 3496 3938 3505
rect 3792 3460 3844 3466
rect 3976 3470 4028 3476
rect 3882 3431 3938 3440
rect 3792 3402 3844 3408
rect 3804 2650 3832 3402
rect 3988 2922 4016 3470
rect 4158 2952 4214 2961
rect 3976 2916 4028 2922
rect 4158 2887 4214 2896
rect 3976 2858 4028 2864
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3804 1465 3832 2246
rect 3790 1456 3846 1465
rect 3790 1391 3846 1400
rect 4172 480 4200 2887
rect 4448 2689 4476 3538
rect 4434 2680 4490 2689
rect 4434 2615 4490 2624
rect 4540 2582 4568 7942
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4540 2310 4568 2382
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 3698 368 3754 377
rect 3698 303 3754 312
rect 4158 0 4214 480
rect 4632 105 4660 4422
rect 4724 2310 4752 8366
rect 4816 8265 4844 8774
rect 4908 8634 4936 9386
rect 5000 9178 5028 12718
rect 5092 12714 5120 13382
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 11762 5212 12582
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11082 5120 11494
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4894 8528 4950 8537
rect 4894 8463 4950 8472
rect 4802 8256 4858 8265
rect 4802 8191 4858 8200
rect 4908 8090 4936 8463
rect 4896 8084 4948 8090
rect 4948 8044 5028 8072
rect 4896 8026 4948 8032
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 5914 4844 7822
rect 5000 7546 5028 8044
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5092 7002 5120 11018
rect 5184 10810 5212 11086
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5276 8922 5304 17031
rect 5368 12986 5396 20159
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6840 19394 6868 23462
rect 6840 19366 6960 19394
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 15910 5488 16594
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 16250 5580 16390
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15638 5488 15846
rect 6380 15706 6408 16186
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5538 15464 5594 15473
rect 5538 15399 5540 15408
rect 5592 15399 5594 15408
rect 5540 15370 5592 15376
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 14958 6040 15506
rect 6840 15162 6868 15642
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6932 15026 6960 19366
rect 7102 16552 7158 16561
rect 7102 16487 7158 16496
rect 7116 15706 7144 16487
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7010 15600 7066 15609
rect 7010 15535 7066 15544
rect 7656 15564 7708 15570
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 14385 5488 14418
rect 5446 14376 5502 14385
rect 5446 14311 5502 14320
rect 5460 13530 5488 14311
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 10606 5396 12786
rect 5460 12102 5488 13330
rect 5552 12850 5580 13670
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5644 12646 5672 12854
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11665 6040 14894
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6104 14074 6132 14350
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6104 13530 6132 14010
rect 6196 13870 6224 14418
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6196 13433 6224 13806
rect 6182 13424 6238 13433
rect 6182 13359 6238 13368
rect 6472 12617 6500 14214
rect 6656 13870 6684 14486
rect 6734 14240 6790 14249
rect 6734 14175 6790 14184
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6458 12608 6514 12617
rect 6458 12543 6514 12552
rect 6472 12442 6500 12543
rect 6564 12481 6592 13126
rect 6656 13025 6684 13806
rect 6642 13016 6698 13025
rect 6642 12951 6698 12960
rect 6550 12472 6606 12481
rect 6460 12436 6512 12442
rect 6550 12407 6606 12416
rect 6460 12378 6512 12384
rect 6090 12336 6146 12345
rect 6090 12271 6092 12280
rect 6144 12271 6146 12280
rect 6092 12242 6144 12248
rect 5998 11656 6054 11665
rect 5448 11620 5500 11626
rect 5998 11591 6054 11600
rect 6184 11620 6236 11626
rect 5448 11562 5500 11568
rect 6184 11562 6236 11568
rect 5460 10810 5488 11562
rect 6196 11354 6224 11562
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5184 8894 5304 8922
rect 5184 8022 5212 8894
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8294 5304 8774
rect 5368 8498 5396 10542
rect 5460 10198 5488 10746
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5460 9722 5488 10134
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8838 5488 9318
rect 5552 8974 5580 11086
rect 6182 10976 6238 10985
rect 5622 10908 5918 10928
rect 6182 10911 6238 10920
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6196 10441 6224 10911
rect 6366 10568 6422 10577
rect 6366 10503 6422 10512
rect 6182 10432 6238 10441
rect 6182 10367 6238 10376
rect 6380 9897 6408 10503
rect 6472 10470 6500 11086
rect 6656 10742 6684 11222
rect 6644 10736 6696 10742
rect 6642 10704 6644 10713
rect 6696 10704 6698 10713
rect 6642 10639 6698 10648
rect 6460 10464 6512 10470
rect 6458 10432 6460 10441
rect 6512 10432 6514 10441
rect 6458 10367 6514 10376
rect 6458 10296 6514 10305
rect 6458 10231 6514 10240
rect 6366 9888 6422 9897
rect 5622 9820 5918 9840
rect 6366 9823 6422 9832
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 8974 6408 9386
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5276 7410 5304 8230
rect 5368 8090 5396 8434
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4986 6624 5042 6633
rect 4986 6559 5042 6568
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5000 4826 5028 6559
rect 5080 6248 5132 6254
rect 5078 6216 5080 6225
rect 5132 6216 5134 6225
rect 5078 6151 5134 6160
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5846 5120 6054
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5092 5710 5120 5782
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5098 5120 5646
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5184 4826 5212 7142
rect 5368 6866 5396 8026
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 6254 5304 6734
rect 5368 6390 5396 6802
rect 5460 6458 5488 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6366 8392 6422 8401
rect 6366 8327 6422 8336
rect 5630 8120 5686 8129
rect 5630 8055 5686 8064
rect 5644 8022 5672 8055
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5644 7732 5672 7958
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 5552 7704 5672 7732
rect 6092 7744 6144 7750
rect 5998 7712 6054 7721
rect 5552 7410 5580 7704
rect 5622 7644 5918 7664
rect 6092 7686 6144 7692
rect 5998 7647 6054 7656
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 7002 5856 7346
rect 6012 7274 6040 7647
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6104 7177 6132 7686
rect 6196 7206 6224 7890
rect 6184 7200 6236 7206
rect 6090 7168 6146 7177
rect 6184 7142 6236 7148
rect 6090 7103 6146 7112
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 6384 5408 6390
rect 5552 6338 5580 6870
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5356 6326 5408 6332
rect 5460 6310 5580 6338
rect 5630 6352 5686 6361
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5460 6186 5488 6310
rect 5630 6287 5632 6296
rect 5684 6287 5686 6296
rect 5632 6258 5684 6264
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5681 5488 6122
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5370 6040 6938
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5000 4321 5028 4626
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4986 4312 5042 4321
rect 5368 4282 5396 4558
rect 4986 4247 4988 4256
rect 5040 4247 5042 4256
rect 5356 4276 5408 4282
rect 4988 4218 5040 4224
rect 5356 4218 5408 4224
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4816 1034 4844 3975
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 3194 5304 3538
rect 5368 3534 5396 4218
rect 5552 4214 5580 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4282 6040 5306
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5460 3670 5488 4014
rect 5552 3738 5580 4150
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 6012 3670 6040 4218
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4894 2680 4950 2689
rect 5368 2650 5396 3470
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 3194 6040 3606
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 4894 2615 4950 2624
rect 5356 2644 5408 2650
rect 4724 1006 4844 1034
rect 4724 480 4752 1006
rect 4908 610 4936 2615
rect 5356 2586 5408 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 1306 6132 6190
rect 6196 5574 6224 6802
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6288 6458 6316 6695
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6196 5302 6224 5510
rect 6288 5370 6316 5714
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6274 5128 6330 5137
rect 6274 5063 6330 5072
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 3194 6224 4422
rect 6288 4146 6316 5063
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6380 4078 6408 8327
rect 6472 6866 6500 10231
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6472 3924 6500 5238
rect 6564 4486 6592 7686
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6254 6776 14175
rect 6840 14074 6868 14894
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6920 12912 6972 12918
rect 6918 12880 6920 12889
rect 6972 12880 6974 12889
rect 6828 12844 6880 12850
rect 6918 12815 6974 12824
rect 6828 12786 6880 12792
rect 6840 12753 6868 12786
rect 6826 12744 6882 12753
rect 6826 12679 6882 12688
rect 6920 12640 6972 12646
rect 6840 12600 6920 12628
rect 6840 11762 6868 12600
rect 6920 12582 6972 12588
rect 6920 12232 6972 12238
rect 6918 12200 6920 12209
rect 6972 12200 6974 12209
rect 6918 12135 6974 12144
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6840 9178 6868 11018
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 10266 6960 10474
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8514 6868 8978
rect 7024 8634 7052 15535
rect 7656 15506 7708 15512
rect 7668 14822 7696 15506
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 12986 7236 13738
rect 7472 13388 7524 13394
rect 7524 13348 7604 13376
rect 7472 13330 7524 13336
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7576 12374 7604 13348
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7288 12300 7340 12306
rect 7340 12260 7420 12288
rect 7288 12242 7340 12248
rect 7392 11694 7420 12260
rect 7380 11688 7432 11694
rect 7378 11656 7380 11665
rect 7432 11656 7434 11665
rect 7378 11591 7434 11600
rect 7102 11248 7158 11257
rect 7102 11183 7158 11192
rect 7116 10266 7144 11183
rect 7392 11150 7420 11591
rect 7576 11558 7604 12310
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9722 7328 10066
rect 7392 10062 7420 10542
rect 7380 10056 7432 10062
rect 7378 10024 7380 10033
rect 7432 10024 7434 10033
rect 7378 9959 7434 9968
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7300 9625 7328 9658
rect 7286 9616 7342 9625
rect 7286 9551 7342 9560
rect 7392 9042 7420 9959
rect 7576 9586 7604 11494
rect 7668 11150 7696 14758
rect 7852 14618 7880 24783
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7944 14618 7972 15098
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13870 7880 14214
rect 7944 14074 7972 14554
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 12850 7788 13398
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7760 11830 7788 12786
rect 7852 11898 7880 13806
rect 8036 13705 8064 14894
rect 8128 14278 8156 15302
rect 8312 15162 8340 25978
rect 10520 25786 10548 27520
rect 10520 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 9310 23080 9366 23089
rect 9310 23015 9366 23024
rect 8758 20360 8814 20369
rect 8758 20295 8814 20304
rect 8482 16008 8538 16017
rect 8482 15943 8538 15952
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8022 13696 8078 13705
rect 8022 13631 8078 13640
rect 8128 13394 8156 14214
rect 8220 13870 8248 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8208 13864 8260 13870
rect 8206 13832 8208 13841
rect 8260 13832 8262 13841
rect 8206 13767 8262 13776
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 8206 11792 8262 11801
rect 8206 11727 8208 11736
rect 8260 11727 8262 11736
rect 8208 11698 8260 11704
rect 8220 11286 8248 11698
rect 8208 11280 8260 11286
rect 8114 11248 8170 11257
rect 8208 11222 8260 11228
rect 8114 11183 8170 11192
rect 8128 11150 8156 11183
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 8116 11144 8168 11150
rect 8312 11098 8340 14010
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8404 12442 8432 12786
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8404 11762 8432 12378
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8496 11354 8524 15943
rect 8574 14376 8630 14385
rect 8574 14311 8630 14320
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8116 11086 8168 11092
rect 8220 11070 8340 11098
rect 7840 11008 7892 11014
rect 8220 10962 8248 11070
rect 7840 10950 7892 10956
rect 7852 10470 7880 10950
rect 8128 10934 8248 10962
rect 8128 10606 8156 10934
rect 8496 10810 8524 11290
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7668 9382 7696 10066
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6840 8486 7052 8514
rect 7116 8498 7144 8842
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7546 6960 7890
rect 7024 7750 7052 8486
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 8090 7420 8230
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6656 4826 6684 6054
rect 6840 5953 6868 6054
rect 6826 5944 6882 5953
rect 6826 5879 6882 5888
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6552 4072 6604 4078
rect 6550 4040 6552 4049
rect 6604 4040 6606 4049
rect 6550 3975 6606 3984
rect 6380 3896 6500 3924
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6196 2009 6224 2246
rect 6182 2000 6238 2009
rect 6182 1935 6238 1944
rect 5828 1278 6132 1306
rect 4896 604 4948 610
rect 4896 546 4948 552
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5276 480 5304 546
rect 5828 480 5856 1278
rect 6380 480 6408 3896
rect 6748 3602 6776 5510
rect 6932 4865 6960 7142
rect 7104 6792 7156 6798
rect 7102 6760 7104 6769
rect 7156 6760 7158 6769
rect 7102 6695 7158 6704
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 6254 7144 6598
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7208 6202 7236 7686
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6322 7420 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7208 6174 7328 6202
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7102 5944 7158 5953
rect 7208 5914 7236 6054
rect 7102 5879 7158 5888
rect 7196 5908 7248 5914
rect 7116 5574 7144 5879
rect 7196 5850 7248 5856
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7208 5370 7236 5850
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6918 4856 6974 4865
rect 6918 4791 6974 4800
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6932 3942 6960 4422
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7116 2990 7144 4422
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6828 2848 6880 2854
rect 6826 2816 6828 2825
rect 6880 2816 6882 2825
rect 6826 2751 6882 2760
rect 6458 2680 6514 2689
rect 7116 2666 7144 2926
rect 6840 2650 7144 2666
rect 7300 2650 7328 6174
rect 7392 6089 7420 6258
rect 7378 6080 7434 6089
rect 7378 6015 7434 6024
rect 7392 5914 7420 6015
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7392 3670 7420 4762
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7484 2802 7512 8599
rect 7668 8498 7696 9318
rect 7852 9042 7880 10406
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7852 8294 7880 8978
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 7410 7880 8230
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 7206 7880 7346
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7760 5234 7788 5335
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7576 3346 7604 5170
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4729 7696 4966
rect 7654 4720 7710 4729
rect 7654 4655 7710 4664
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 4282 7788 4558
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7760 3738 7788 4218
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3466 7880 7142
rect 7944 6662 7972 7958
rect 8220 7002 8248 10542
rect 8588 9926 8616 14311
rect 8772 13938 8800 20295
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13530 8800 13874
rect 9048 13530 9076 14010
rect 9140 13870 9168 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8772 12986 8800 13330
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12442 8984 12718
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9036 11688 9088 11694
rect 8758 11656 8814 11665
rect 9036 11630 9088 11636
rect 8758 11591 8814 11600
rect 8772 9994 8800 11591
rect 8942 11248 8998 11257
rect 8942 11183 8998 11192
rect 8956 10810 8984 11183
rect 9048 11014 9076 11630
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9048 10266 9076 10950
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8390 9616 8446 9625
rect 8390 9551 8446 9560
rect 8298 8528 8354 8537
rect 8298 8463 8354 8472
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8208 6792 8260 6798
rect 8312 6780 8340 8463
rect 8404 6866 8432 9551
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8680 8838 8708 9386
rect 8758 8936 8814 8945
rect 8758 8871 8814 8880
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8482 8256 8538 8265
rect 8482 8191 8538 8200
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8260 6752 8340 6780
rect 8208 6734 8260 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7944 3738 7972 6598
rect 8220 6225 8248 6598
rect 8312 6458 8340 6752
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8206 6216 8262 6225
rect 8206 6151 8262 6160
rect 8220 5914 8248 6151
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8312 5794 8340 6394
rect 8404 5846 8432 6802
rect 8220 5778 8340 5794
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8208 5772 8340 5778
rect 8260 5766 8340 5772
rect 8208 5714 8260 5720
rect 8312 5370 8340 5766
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8298 5264 8354 5273
rect 8298 5199 8354 5208
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4078 8064 4626
rect 8116 4616 8168 4622
rect 8114 4584 8116 4593
rect 8168 4584 8170 4593
rect 8114 4519 8170 4528
rect 8024 4072 8076 4078
rect 8022 4040 8024 4049
rect 8076 4040 8078 4049
rect 8022 3975 8078 3984
rect 8312 3913 8340 5199
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 8496 3754 8524 8191
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 7546 8616 7822
rect 8680 7818 8708 8774
rect 8772 8634 8800 8871
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8680 7546 8708 7754
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6497 8616 6802
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8574 6488 8630 6497
rect 8574 6423 8576 6432
rect 8628 6423 8630 6432
rect 8576 6394 8628 6400
rect 8680 6225 8708 6598
rect 8864 6458 8892 8298
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 9036 6248 9088 6254
rect 8666 6216 8722 6225
rect 9036 6190 9088 6196
rect 8666 6151 8722 6160
rect 9048 5914 9076 6190
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4078 8708 4422
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8404 3726 8524 3754
rect 8298 3632 8354 3641
rect 8298 3567 8300 3576
rect 8352 3567 8354 3576
rect 8300 3538 8352 3544
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7576 3318 7880 3346
rect 7484 2774 7595 2802
rect 7567 2666 7595 2774
rect 6458 2615 6460 2624
rect 6512 2615 6514 2624
rect 6828 2644 7144 2650
rect 6460 2586 6512 2592
rect 6880 2638 7144 2644
rect 7288 2644 7340 2650
rect 6828 2586 6880 2592
rect 7567 2638 7604 2666
rect 7288 2586 7340 2592
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6932 480 6960 2382
rect 7576 480 7604 2638
rect 7852 1442 7880 3318
rect 8036 3126 8064 3470
rect 8312 3194 8340 3538
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8024 3120 8076 3126
rect 8022 3088 8024 3097
rect 8076 3088 8078 3097
rect 8022 3023 8078 3032
rect 8206 2544 8262 2553
rect 8024 2508 8076 2514
rect 8206 2479 8208 2488
rect 8024 2450 8076 2456
rect 8260 2479 8262 2488
rect 8208 2450 8260 2456
rect 8036 1601 8064 2450
rect 8022 1592 8078 1601
rect 8022 1527 8078 1536
rect 7852 1414 8156 1442
rect 8404 1426 8432 3726
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8496 2446 8524 3470
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 2825 8616 3334
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8128 480 8156 1414
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8680 480 8708 3878
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3058 8800 3538
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8864 2310 8892 2858
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 1873 8892 2246
rect 8850 1864 8906 1873
rect 8850 1799 8906 1808
rect 9048 1737 9076 3946
rect 9140 2689 9168 12650
rect 9232 9178 9260 14758
rect 9324 10810 9352 23015
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 20505 10824 25758
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 12346 24712 12402 24721
rect 12346 24647 12402 24656
rect 10782 20496 10838 20505
rect 10782 20431 10838 20440
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 11886 17776 11942 17785
rect 11886 17711 11942 17720
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10138 16144 10194 16153
rect 10138 16079 10194 16088
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 12306 9444 15846
rect 10048 15496 10100 15502
rect 9494 15464 9550 15473
rect 10048 15438 10100 15444
rect 9494 15399 9550 15408
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9508 12186 9536 15399
rect 9770 13696 9826 13705
rect 9770 13631 9826 13640
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9586 13016 9642 13025
rect 9586 12951 9642 12960
rect 9600 12322 9628 12951
rect 9692 12442 9720 13330
rect 9784 13161 9812 13631
rect 9954 13288 10010 13297
rect 9954 13223 10010 13232
rect 9864 13184 9916 13190
rect 9770 13152 9826 13161
rect 9864 13126 9916 13132
rect 9770 13087 9826 13096
rect 9876 12782 9904 13126
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9600 12294 9720 12322
rect 9416 12158 9536 12186
rect 9416 11642 9444 12158
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11762 9536 12038
rect 9692 11778 9720 12294
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11898 9812 12242
rect 9968 12238 9996 13223
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11898 9996 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9496 11756 9548 11762
rect 9692 11750 9812 11778
rect 9496 11698 9548 11704
rect 9416 11614 9536 11642
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11218 9444 11494
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9508 10010 9536 11614
rect 9586 11384 9642 11393
rect 9586 11319 9642 11328
rect 9324 9982 9536 10010
rect 9324 9353 9352 9982
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9382 9444 9862
rect 9404 9376 9456 9382
rect 9310 9344 9366 9353
rect 9404 9318 9456 9324
rect 9310 9279 9366 9288
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9232 8430 9260 9114
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9232 7342 9260 8026
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3233 9260 3878
rect 9218 3224 9274 3233
rect 9218 3159 9274 3168
rect 9324 3108 9352 9279
rect 9416 8838 9444 9318
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 6361 9444 8774
rect 9600 8022 9628 11319
rect 9680 11008 9732 11014
rect 9678 10976 9680 10985
rect 9732 10976 9734 10985
rect 9678 10911 9734 10920
rect 9678 10704 9734 10713
rect 9678 10639 9734 10648
rect 9692 9994 9720 10639
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9678 9072 9734 9081
rect 9678 9007 9680 9016
rect 9732 9007 9734 9016
rect 9680 8978 9732 8984
rect 9784 8786 9812 11750
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11286 9996 11494
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 11064 9904 11154
rect 9876 11036 9996 11064
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 9692 8758 9812 8786
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9402 6352 9458 6361
rect 9402 6287 9458 6296
rect 9416 5953 9444 6287
rect 9402 5944 9458 5953
rect 9508 5914 9536 7142
rect 9600 6866 9628 7142
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 6769 9628 6802
rect 9586 6760 9642 6769
rect 9586 6695 9642 6704
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9402 5879 9458 5888
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9508 4690 9536 5850
rect 9600 5030 9628 6190
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9692 4706 9720 8758
rect 9876 8673 9904 10911
rect 9968 10130 9996 11036
rect 10060 10810 10088 15438
rect 10152 15162 10180 16079
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15162 10824 16390
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 11072 15026 11100 15302
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10152 11898 10180 13262
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11082 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 13767
rect 10888 13734 10916 14418
rect 11532 14278 11560 15438
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13326 10916 13670
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10876 13184 10928 13190
rect 10980 13172 11008 14214
rect 11716 13954 11744 15846
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 15162 11836 15506
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 14618 11836 15098
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11808 14074 11836 14554
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11060 13932 11112 13938
rect 11716 13926 11836 13954
rect 11060 13874 11112 13880
rect 10928 13144 11008 13172
rect 10876 13126 10928 13132
rect 10888 12782 10916 13126
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10796 12238 10824 12650
rect 11072 12646 11100 13874
rect 11702 12880 11758 12889
rect 11702 12815 11758 12824
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12306 11100 12582
rect 11716 12481 11744 12815
rect 11702 12472 11758 12481
rect 11702 12407 11704 12416
rect 11756 12407 11758 12416
rect 11704 12378 11756 12384
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11610 12336 11666 12345
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 11072 11762 11100 12242
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11830 11284 12038
rect 11348 11898 11376 12310
rect 11610 12271 11666 12280
rect 11336 11892 11388 11898
rect 11388 11852 11560 11880
rect 11336 11834 11388 11840
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10874 11520 10930 11529
rect 10796 11393 10824 11494
rect 10874 11455 10930 11464
rect 10782 11384 10838 11393
rect 10692 11348 10744 11354
rect 10782 11319 10838 11328
rect 10692 11290 10744 11296
rect 10322 11112 10378 11121
rect 10140 11076 10192 11082
rect 10322 11047 10378 11056
rect 10140 11018 10192 11024
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10060 10606 10088 10746
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10048 10464 10100 10470
rect 10046 10432 10048 10441
rect 10100 10432 10102 10441
rect 10046 10367 10102 10376
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 10060 10198 10088 10231
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 9042 9996 10066
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9862 8664 9918 8673
rect 9862 8599 9918 8608
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 8401 9812 8502
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9784 6866 9812 7346
rect 9876 6934 9904 8055
rect 9956 7880 10008 7886
rect 10060 7868 10088 9862
rect 10152 9761 10180 11018
rect 10336 10810 10364 11047
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10784 10736 10836 10742
rect 10230 10704 10286 10713
rect 10784 10678 10836 10684
rect 10230 10639 10232 10648
rect 10284 10639 10286 10648
rect 10232 10610 10284 10616
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10138 9752 10194 9761
rect 10138 9687 10194 9696
rect 10704 9518 10732 10406
rect 10796 10266 10824 10678
rect 10888 10282 10916 11455
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10980 10962 11008 11154
rect 10980 10934 11100 10962
rect 11072 10470 11100 10934
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11060 10464 11112 10470
rect 11164 10441 11192 10474
rect 11060 10406 11112 10412
rect 11150 10432 11206 10441
rect 11150 10367 11206 10376
rect 11426 10432 11482 10441
rect 11426 10367 11482 10376
rect 11150 10296 11206 10305
rect 10784 10260 10836 10266
rect 10888 10254 11008 10282
rect 10784 10202 10836 10208
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10796 9466 10824 10202
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9654 10916 10066
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9178 10732 9454
rect 10796 9438 10916 9466
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8430 10272 8774
rect 10796 8430 10824 9318
rect 10888 9110 10916 9438
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10888 8634 10916 9046
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 8537 11008 10254
rect 11150 10231 11206 10240
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10966 8528 11022 8537
rect 10966 8463 11022 8472
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10138 8256 10194 8265
rect 10690 8256 10746 8265
rect 10138 8191 10194 8200
rect 10008 7840 10088 7868
rect 9956 7822 10008 7828
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9968 6798 9996 7822
rect 10152 7818 10180 8191
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10048 7744 10100 7750
rect 10336 7721 10364 7890
rect 10048 7686 10100 7692
rect 10138 7712 10194 7721
rect 10060 7585 10088 7686
rect 10138 7647 10194 7656
rect 10322 7712 10378 7721
rect 10322 7647 10378 7656
rect 10046 7576 10102 7585
rect 10046 7511 10102 7520
rect 10152 7478 10180 7647
rect 10336 7546 10364 7647
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10704 7313 10732 8191
rect 10980 8090 11008 8298
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10690 7304 10746 7313
rect 10690 7239 10746 7248
rect 10888 7206 10916 7686
rect 11072 7546 11100 9318
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 9956 6792 10008 6798
rect 10008 6752 10088 6780
rect 9956 6734 10008 6740
rect 10060 6186 10088 6752
rect 10244 6458 10272 6802
rect 10232 6452 10284 6458
rect 10152 6412 10232 6440
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9954 5672 10010 5681
rect 9784 5370 9812 5646
rect 9954 5607 9956 5616
rect 10008 5607 10010 5616
rect 9956 5578 10008 5584
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 4826 9812 5306
rect 9954 5264 10010 5273
rect 9954 5199 10010 5208
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9496 4684 9548 4690
rect 9692 4678 9812 4706
rect 9496 4626 9548 4632
rect 9588 4072 9640 4078
rect 9640 4032 9720 4060
rect 9588 4014 9640 4020
rect 9232 3080 9352 3108
rect 9126 2680 9182 2689
rect 9126 2615 9182 2624
rect 9034 1728 9090 1737
rect 9034 1663 9090 1672
rect 9232 480 9260 3080
rect 9692 2650 9720 4032
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 480 9812 4678
rect 9876 4282 9904 5034
rect 9968 5001 9996 5199
rect 9954 4992 10010 5001
rect 9954 4927 10010 4936
rect 10060 4758 10088 6122
rect 10152 5302 10180 6412
rect 10232 6394 10284 6400
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5296 10192 5302
rect 10704 5273 10732 7142
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10876 6656 10928 6662
rect 10796 6604 10876 6610
rect 10796 6598 10928 6604
rect 10796 6582 10916 6598
rect 10796 5710 10824 6582
rect 11072 6361 11100 6666
rect 11164 6458 11192 10231
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11072 6066 11100 6287
rect 11164 6254 11192 6394
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11072 6038 11192 6066
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5370 10824 5646
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10140 5238 10192 5244
rect 10690 5264 10746 5273
rect 11072 5250 11100 5578
rect 11164 5574 11192 6038
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10690 5199 10746 5208
rect 10980 5222 11100 5250
rect 10980 5166 11008 5222
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10980 4826 11008 4966
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3777 9904 3878
rect 9862 3768 9918 3777
rect 9862 3703 9918 3712
rect 10060 3670 10088 4694
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4282 10824 4626
rect 10980 4282 11008 4762
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10796 4162 10824 4218
rect 10796 4134 11008 4162
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10704 3913 10732 3946
rect 10690 3904 10746 3913
rect 10289 3836 10585 3856
rect 10690 3839 10746 3848
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3777 10824 4014
rect 10782 3768 10838 3777
rect 10692 3732 10744 3738
rect 10980 3738 11008 4134
rect 10782 3703 10838 3712
rect 10968 3732 11020 3738
rect 10692 3674 10744 3680
rect 10968 3674 11020 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9968 3194 9996 3538
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2446 10732 3674
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10692 2440 10744 2446
rect 10322 2408 10378 2417
rect 10692 2382 10744 2388
rect 10322 2343 10378 2352
rect 10336 480 10364 2343
rect 10796 2281 10824 3130
rect 10874 2408 10930 2417
rect 10874 2343 10876 2352
rect 10928 2343 10930 2352
rect 10876 2314 10928 2320
rect 10782 2272 10838 2281
rect 10782 2207 10838 2216
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 10888 480 10916 1527
rect 11072 1465 11100 5034
rect 11256 3194 11284 8327
rect 11440 6866 11468 10367
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11334 6352 11390 6361
rect 11334 6287 11390 6296
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11348 3058 11376 6287
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5953 11468 6054
rect 11426 5944 11482 5953
rect 11426 5879 11482 5888
rect 11532 5778 11560 11852
rect 11624 10742 11652 12271
rect 11716 11898 11744 12378
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11716 10169 11744 11018
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 11808 9466 11836 13926
rect 11624 9438 11836 9466
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11624 5001 11652 9438
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 9178 11836 9318
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11900 8634 11928 17711
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16046 12112 16390
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12176 15978 12204 16934
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12268 15910 12296 16730
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 12646 12204 13398
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11992 10554 12020 12582
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11354 12112 12174
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10810 12112 10950
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11992 10526 12112 10554
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 9926 12020 10406
rect 12084 10130 12112 10526
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11992 8498 12020 9862
rect 12084 9722 12112 10066
rect 12162 10024 12218 10033
rect 12162 9959 12218 9968
rect 12176 9926 12204 9959
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9761 12204 9862
rect 12162 9752 12218 9761
rect 12072 9716 12124 9722
rect 12162 9687 12218 9696
rect 12072 9658 12124 9664
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 8838 12112 9522
rect 12176 9489 12204 9590
rect 12162 9480 12218 9489
rect 12162 9415 12164 9424
rect 12216 9415 12218 9424
rect 12164 9386 12216 9392
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12084 8634 12112 8774
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12176 8430 12204 8774
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12268 8072 12296 15846
rect 12360 10146 12388 24647
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 17038 20496 17094 20505
rect 17038 20431 17094 20440
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 16946 19272 17002 19281
rect 16946 19207 17002 19216
rect 15566 18864 15622 18873
rect 15566 18799 15622 18808
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 12622 18320 12678 18329
rect 12622 18255 12678 18264
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16114 12572 16390
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15745 12480 15846
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12452 15094 12480 15574
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14346 12480 14894
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13870 12572 14214
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12636 13462 12664 18255
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17134 13124 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12624 13456 12676 13462
rect 12530 13424 12586 13433
rect 12624 13398 12676 13404
rect 12530 13359 12532 13368
rect 12584 13359 12586 13368
rect 12532 13330 12584 13336
rect 12544 12986 12572 13330
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11824 12492 11830
rect 12438 11792 12440 11801
rect 12492 11792 12494 11801
rect 12544 11762 12572 12038
rect 12438 11727 12494 11736
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12544 11665 12572 11698
rect 12624 11688 12676 11694
rect 12530 11656 12586 11665
rect 12624 11630 12676 11636
rect 12530 11591 12586 11600
rect 12636 11286 12664 11630
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 11121 12664 11222
rect 12622 11112 12678 11121
rect 12622 11047 12678 11056
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12360 10118 12480 10146
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12360 9518 12388 9930
rect 12452 9518 12480 10118
rect 12544 9926 12572 10610
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12084 8044 12296 8072
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7002 11744 7346
rect 11808 7206 11836 7890
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11610 4992 11666 5001
rect 11610 4927 11666 4936
rect 11716 4842 11744 6802
rect 11808 6662 11836 7142
rect 11978 7032 12034 7041
rect 11978 6967 12034 6976
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11900 6118 11928 6802
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11992 5914 12020 6967
rect 12084 6882 12112 8044
rect 12452 7970 12480 8230
rect 12544 8090 12572 9862
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12622 9480 12678 9489
rect 12622 9415 12678 9424
rect 12636 8634 12664 9415
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12176 7942 12480 7970
rect 12176 7857 12204 7942
rect 12162 7848 12218 7857
rect 12162 7783 12218 7792
rect 12164 7472 12216 7478
rect 12162 7440 12164 7449
rect 12216 7440 12218 7449
rect 12162 7375 12218 7384
rect 12360 6984 12388 7942
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7342 12480 7686
rect 12544 7546 12572 8026
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12440 7336 12492 7342
rect 12438 7304 12440 7313
rect 12492 7304 12494 7313
rect 12438 7239 12494 7248
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12440 6996 12492 7002
rect 12360 6956 12440 6984
rect 12084 6854 12296 6882
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12162 6760 12218 6769
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11440 4814 11744 4842
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11242 2680 11298 2689
rect 11242 2615 11244 2624
rect 11296 2615 11298 2624
rect 11244 2586 11296 2592
rect 11058 1456 11114 1465
rect 11058 1391 11114 1400
rect 11440 480 11468 4814
rect 11808 4486 11836 5510
rect 11900 5098 11928 5714
rect 11992 5370 12020 5850
rect 12084 5710 12112 6734
rect 12162 6695 12164 6704
rect 12216 6695 12218 6704
rect 12164 6666 12216 6672
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5817 12204 6054
rect 12162 5808 12218 5817
rect 12162 5743 12218 5752
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 12084 5030 12112 5646
rect 12268 5234 12296 6854
rect 12360 6458 12388 6956
rect 12440 6938 12492 6944
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12438 4992 12494 5001
rect 12438 4927 12494 4936
rect 12452 4758 12480 4927
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12256 4616 12308 4622
rect 11978 4584 12034 4593
rect 12256 4558 12308 4564
rect 11978 4519 12034 4528
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11808 4321 11836 4422
rect 11794 4312 11850 4321
rect 11794 4247 11850 4256
rect 11518 4176 11574 4185
rect 11518 4111 11574 4120
rect 11532 3738 11560 4111
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11532 2514 11560 3674
rect 11900 3534 11928 3878
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3194 11928 3470
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1465 11652 2246
rect 11610 1456 11666 1465
rect 11610 1391 11666 1400
rect 11992 480 12020 4519
rect 12162 4040 12218 4049
rect 12162 3975 12218 3984
rect 12176 610 12204 3975
rect 12268 3670 12296 4558
rect 12360 4078 12388 4694
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12268 2990 12296 3606
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12268 2446 12296 2926
rect 12360 2650 12388 3606
rect 12544 3466 12572 6190
rect 12636 3505 12664 7142
rect 12728 4826 12756 16390
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15434 12848 15846
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 14074 12848 14826
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13530 12848 13670
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11558 12848 11834
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11014 12848 11494
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10169 12848 10406
rect 12806 10160 12862 10169
rect 12806 10095 12862 10104
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12820 8362 12848 9590
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12806 8256 12862 8265
rect 12806 8191 12862 8200
rect 12820 7721 12848 8191
rect 12806 7712 12862 7721
rect 12806 7647 12862 7656
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12728 4078 12756 4762
rect 12820 4457 12848 7142
rect 12912 5794 12940 16934
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 14822 13032 16050
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 14550 13032 14758
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14074 13032 14486
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13004 9110 13032 13466
rect 13096 9353 13124 17070
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 13188 15450 13216 16623
rect 13280 15586 13308 17002
rect 13372 16590 13400 17138
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 15978 13400 16526
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13372 15706 13400 15914
rect 13464 15910 13492 16594
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 15978 14136 16390
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 13452 15904 13504 15910
rect 13912 15904 13964 15910
rect 13452 15846 13504 15852
rect 13542 15872 13598 15881
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13464 15609 13492 15846
rect 13912 15846 13964 15852
rect 13542 15807 13598 15816
rect 13450 15600 13506 15609
rect 13280 15558 13400 15586
rect 13188 15422 13308 15450
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 14958 13216 15302
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12306 13216 13126
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 11898 13216 12242
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13174 11792 13230 11801
rect 13174 11727 13230 11736
rect 13188 10713 13216 11727
rect 13280 11694 13308 15422
rect 13372 12442 13400 15558
rect 13450 15535 13506 15544
rect 13556 14362 13584 15807
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 15366 13676 15506
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13740 15314 13768 15370
rect 13648 15094 13676 15302
rect 13740 15286 13860 15314
rect 13832 15162 13860 15286
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13648 14482 13676 15030
rect 13924 14770 13952 15846
rect 13832 14742 13952 14770
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13556 14334 13676 14362
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11354 13308 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13464 11257 13492 13806
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 13530 13584 13738
rect 13648 13530 13676 14334
rect 13726 13560 13782 13569
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13636 13524 13688 13530
rect 13726 13495 13782 13504
rect 13636 13466 13688 13472
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13450 11248 13506 11257
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13360 11212 13412 11218
rect 13450 11183 13506 11192
rect 13360 11154 13412 11160
rect 13174 10704 13230 10713
rect 13174 10639 13230 10648
rect 13188 9654 13216 10639
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13082 9344 13138 9353
rect 13082 9279 13138 9288
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8090 13032 8910
rect 13188 8634 13216 9454
rect 13280 9042 13308 11154
rect 13372 10470 13400 11154
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13096 7936 13124 8298
rect 13280 8090 13308 8842
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13004 7908 13124 7936
rect 13004 5914 13032 7908
rect 13268 7880 13320 7886
rect 13082 7848 13138 7857
rect 13268 7822 13320 7828
rect 13082 7783 13138 7792
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12912 5766 13032 5794
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12912 5370 12940 5578
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12806 4448 12862 4457
rect 12806 4383 12862 4392
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 13004 4010 13032 5766
rect 13096 4049 13124 7783
rect 13280 7002 13308 7822
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13082 4040 13138 4049
rect 12992 4004 13044 4010
rect 13082 3975 13138 3984
rect 12992 3946 13044 3952
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12728 3534 12756 3878
rect 12716 3528 12768 3534
rect 12622 3496 12678 3505
rect 12532 3460 12584 3466
rect 12716 3470 12768 3476
rect 12622 3431 12678 3440
rect 12532 3402 12584 3408
rect 12728 2990 12756 3470
rect 12912 3398 12940 3878
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13096 3194 13124 3470
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12716 2984 12768 2990
rect 13096 2972 13124 3130
rect 12716 2926 12768 2932
rect 13004 2944 13124 2972
rect 13004 2854 13032 2944
rect 13188 2904 13216 6394
rect 13266 5264 13322 5273
rect 13266 5199 13322 5208
rect 13280 5098 13308 5199
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13372 3913 13400 10406
rect 13464 9042 13492 10610
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13464 7954 13492 8978
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7206 13492 7754
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13450 6216 13506 6225
rect 13450 6151 13506 6160
rect 13464 4457 13492 6151
rect 13450 4448 13506 4457
rect 13450 4383 13506 4392
rect 13450 4312 13506 4321
rect 13450 4247 13506 4256
rect 13358 3904 13414 3913
rect 13358 3839 13414 3848
rect 13464 3670 13492 4247
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13096 2876 13216 2904
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 13004 2582 13032 2790
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12636 2106 12664 2382
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 12164 604 12216 610
rect 12164 546 12216 552
rect 12532 604 12584 610
rect 12532 546 12584 552
rect 12544 480 12572 546
rect 13096 480 13124 2876
rect 13556 2836 13584 12922
rect 13740 12850 13768 13495
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 11218 13860 14742
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13394 13952 13670
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 11898 13952 13330
rect 14016 12782 14044 14418
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14016 12374 14044 12718
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14016 11694 14044 12310
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11286 14044 11630
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13740 10962 13768 11086
rect 13740 10934 13860 10962
rect 13634 10704 13690 10713
rect 13634 10639 13690 10648
rect 13648 8294 13676 10639
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 9217 13768 10406
rect 13832 9761 13860 10934
rect 14016 10674 14044 11086
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13818 9752 13874 9761
rect 13818 9687 13874 9696
rect 13726 9208 13782 9217
rect 13832 9178 13860 9687
rect 13726 9143 13782 9152
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13636 8016 13688 8022
rect 13634 7984 13636 7993
rect 13688 7984 13690 7993
rect 13634 7919 13690 7928
rect 13740 7834 13768 8298
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13648 7806 13768 7834
rect 13648 7342 13676 7806
rect 13832 7342 13860 8230
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13648 7177 13676 7278
rect 13634 7168 13690 7177
rect 13634 7103 13690 7112
rect 13832 6798 13860 7278
rect 13924 7274 13952 8298
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14108 6934 14136 15914
rect 14200 15094 14228 16594
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14200 12782 14228 13874
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12102 14228 12718
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 9926 14228 10406
rect 14188 9920 14240 9926
rect 14186 9888 14188 9897
rect 14240 9888 14242 9897
rect 14186 9823 14242 9832
rect 14096 6928 14148 6934
rect 14002 6896 14058 6905
rect 13912 6860 13964 6866
rect 14096 6870 14148 6876
rect 14002 6831 14058 6840
rect 13912 6802 13964 6808
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5914 13676 6122
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13648 5234 13676 5714
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 4146 13676 4422
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13740 3618 13768 6054
rect 13832 5370 13860 6054
rect 13924 5681 13952 6802
rect 14016 5914 14044 6831
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13910 5672 13966 5681
rect 13910 5607 13966 5616
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14016 4826 14044 5850
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14108 4185 14136 6734
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14200 5710 14228 6666
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5234 14228 5646
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14292 4826 14320 15846
rect 14568 15706 14596 16050
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14890 14688 15302
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14646 14784 14702 14793
rect 14646 14719 14702 14728
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 11150 14412 14214
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13462 14504 13670
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 12646 14504 13262
rect 14660 13138 14688 14719
rect 14752 14618 14780 14962
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 14249 14780 14350
rect 14738 14240 14794 14249
rect 14738 14175 14794 14184
rect 14752 14074 14780 14175
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14568 13110 14688 13138
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10577 14412 10950
rect 14370 10568 14426 10577
rect 14370 10503 14426 10512
rect 14384 10266 14412 10503
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14476 10033 14504 10134
rect 14462 10024 14518 10033
rect 14462 9959 14518 9968
rect 14464 9648 14516 9654
rect 14462 9616 14464 9625
rect 14516 9616 14518 9625
rect 14462 9551 14518 9560
rect 14568 9353 14596 13110
rect 14752 12442 14780 13398
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 11898 14780 12242
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14660 10305 14688 10775
rect 14646 10296 14702 10305
rect 14646 10231 14702 10240
rect 14554 9344 14610 9353
rect 14554 9279 14610 9288
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14384 8430 14412 8842
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14462 7576 14518 7585
rect 14462 7511 14518 7520
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6322 14412 7142
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14384 5846 14412 6258
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14384 5370 14412 5782
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14094 4176 14150 4185
rect 14094 4111 14150 4120
rect 14292 4078 14320 4762
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 3738 14044 3878
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14476 3641 14504 7511
rect 14568 6458 14596 9279
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14554 6080 14610 6089
rect 14554 6015 14610 6024
rect 14462 3632 14518 3641
rect 13740 3602 13860 3618
rect 13740 3596 13872 3602
rect 13740 3590 13820 3596
rect 14462 3567 14518 3576
rect 13820 3538 13872 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13648 2961 13676 3470
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13634 2952 13690 2961
rect 13634 2887 13690 2896
rect 13464 2808 13584 2836
rect 13740 2825 13768 3334
rect 13832 3058 13860 3538
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13924 2922 13952 3334
rect 14200 3097 14228 3334
rect 14186 3088 14242 3097
rect 14186 3023 14242 3032
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13726 2816 13782 2825
rect 13464 2666 13492 2808
rect 13726 2751 13782 2760
rect 13464 2638 13676 2666
rect 13648 480 13676 2638
rect 14476 2582 14504 2994
rect 14568 2961 14596 6015
rect 14660 5914 14688 10231
rect 14752 8888 14780 11834
rect 14844 10810 14872 15914
rect 15382 15736 15438 15745
rect 15382 15671 15438 15680
rect 15016 15496 15068 15502
rect 15014 15464 15016 15473
rect 15068 15464 15070 15473
rect 15014 15399 15070 15408
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 14657 15056 14758
rect 15014 14648 15070 14657
rect 15014 14583 15070 14592
rect 15014 14376 15070 14385
rect 15014 14311 15016 14320
rect 15068 14311 15070 14320
rect 15016 14282 15068 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13977 15332 15302
rect 15106 13968 15162 13977
rect 15106 13903 15162 13912
rect 15290 13968 15346 13977
rect 15290 13903 15346 13912
rect 15120 13870 15148 13903
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15396 13394 15424 15671
rect 15474 14920 15530 14929
rect 15474 14855 15530 14864
rect 15488 14074 15516 14855
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15580 14006 15608 18799
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16868 16998 16896 17682
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15948 15502 15976 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15660 14816 15712 14822
rect 15658 14784 15660 14793
rect 15712 14784 15714 14793
rect 15658 14719 15714 14728
rect 15764 14385 15792 15438
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15750 14376 15806 14385
rect 15750 14311 15806 14320
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15120 13274 15148 13330
rect 15476 13320 15528 13326
rect 15120 13246 15424 13274
rect 15476 13262 15528 13268
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15292 12640 15344 12646
rect 15106 12608 15162 12617
rect 15292 12582 15344 12588
rect 15106 12543 15162 12552
rect 15120 12442 15148 12543
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14924 11688 14976 11694
rect 14922 11656 14924 11665
rect 14976 11656 14978 11665
rect 15304 11626 15332 12582
rect 14922 11591 14978 11600
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15304 11354 15332 11562
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 13246
rect 15488 12889 15516 13262
rect 15474 12880 15530 12889
rect 15474 12815 15530 12824
rect 15580 12442 15608 13330
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 14844 10606 14872 10746
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 9994 15332 10474
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9738 15332 9930
rect 15384 9920 15436 9926
rect 15382 9888 15384 9897
rect 15436 9888 15438 9897
rect 15382 9823 15438 9832
rect 15304 9710 15424 9738
rect 14832 9376 14884 9382
rect 14830 9344 14832 9353
rect 14884 9344 14886 9353
rect 14830 9279 14886 9288
rect 14752 8860 14872 8888
rect 14844 7954 14872 8860
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8401 15332 8774
rect 15290 8392 15346 8401
rect 15290 8327 15346 8336
rect 14832 7948 14884 7954
rect 14752 7908 14832 7936
rect 14752 7721 14780 7908
rect 14832 7890 14884 7896
rect 14832 7744 14884 7750
rect 14738 7712 14794 7721
rect 14832 7686 14884 7692
rect 14738 7647 14794 7656
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14648 5704 14700 5710
rect 14646 5672 14648 5681
rect 14700 5672 14702 5681
rect 14646 5607 14702 5616
rect 14752 4570 14780 6870
rect 14844 6662 14872 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6390 15332 6802
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15304 5914 15332 6326
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15028 5556 15056 5850
rect 15028 5528 15332 5556
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5302 15332 5528
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15396 4842 15424 9710
rect 15488 7426 15516 11018
rect 15580 11014 15608 12038
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10674 15608 10950
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15672 10606 15700 14214
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15764 12442 15792 13942
rect 15856 12866 15884 14894
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 13734 15976 14214
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13569 15976 13670
rect 15934 13560 15990 13569
rect 15934 13495 15990 13504
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 12986 15976 13330
rect 16040 13326 16068 14418
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16132 13954 16160 14350
rect 16224 14113 16252 14758
rect 16210 14104 16266 14113
rect 16210 14039 16266 14048
rect 16132 13938 16252 13954
rect 16132 13932 16264 13938
rect 16132 13926 16212 13932
rect 16212 13874 16264 13880
rect 16028 13320 16080 13326
rect 16026 13288 16028 13297
rect 16080 13288 16082 13297
rect 16026 13223 16082 13232
rect 16224 13190 16252 13874
rect 16212 13184 16264 13190
rect 16210 13152 16212 13161
rect 16264 13152 16266 13161
rect 16210 13087 16266 13096
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16212 12912 16264 12918
rect 15856 12838 16068 12866
rect 16212 12854 16264 12860
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15934 12064 15990 12073
rect 15934 11999 15990 12008
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10266 15700 10542
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15658 9208 15714 9217
rect 15764 9178 15792 11222
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 10062 15884 10406
rect 15948 10266 15976 11999
rect 16040 11393 16068 12838
rect 16224 11898 16252 12854
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16026 11384 16082 11393
rect 16026 11319 16082 11328
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15856 9761 15884 9998
rect 16132 9926 16160 11154
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15842 9752 15898 9761
rect 15842 9687 15898 9696
rect 15658 9143 15660 9152
rect 15712 9143 15714 9152
rect 15752 9172 15804 9178
rect 15660 9114 15712 9120
rect 15752 9114 15804 9120
rect 15672 8090 15700 9114
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15764 8022 15792 9114
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8634 15884 8910
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 7449 15884 7822
rect 15842 7440 15898 7449
rect 15488 7398 15792 7426
rect 15474 7304 15530 7313
rect 15474 7239 15530 7248
rect 15488 6798 15516 7239
rect 15568 7200 15620 7206
rect 15566 7168 15568 7177
rect 15620 7168 15622 7177
rect 15566 7103 15622 7112
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15580 6254 15608 7103
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5574 15608 6190
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15396 4814 15516 4842
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 14660 4542 14780 4570
rect 14660 3777 14688 4542
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14646 3768 14702 3777
rect 14646 3703 14702 3712
rect 14752 2990 14780 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4078 15332 4422
rect 15396 4282 15424 4694
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15304 3738 15332 4014
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15396 3670 15424 4218
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 2984 14792 2990
rect 14554 2952 14610 2961
rect 14740 2926 14792 2932
rect 14830 2952 14886 2961
rect 14554 2887 14610 2896
rect 14830 2887 14886 2896
rect 15106 2952 15162 2961
rect 15106 2887 15108 2896
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14660 2689 14688 2790
rect 14646 2680 14702 2689
rect 14646 2615 14702 2624
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14004 2304 14056 2310
rect 14476 2281 14504 2518
rect 14004 2246 14056 2252
rect 14462 2272 14518 2281
rect 14016 1873 14044 2246
rect 14462 2207 14518 2216
rect 14002 1864 14058 1873
rect 14002 1799 14058 1808
rect 14278 1320 14334 1329
rect 14278 1255 14334 1264
rect 14292 480 14320 1255
rect 14844 480 14872 2887
rect 15160 2887 15162 2896
rect 15108 2858 15160 2864
rect 15304 2582 15332 3402
rect 15488 3210 15516 4814
rect 15580 4690 15608 5510
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15672 4282 15700 6122
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15764 4049 15792 7398
rect 15842 7375 15898 7384
rect 15842 5400 15898 5409
rect 15842 5335 15844 5344
rect 15896 5335 15898 5344
rect 15844 5306 15896 5312
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15844 3936 15896 3942
rect 15842 3904 15844 3913
rect 15896 3904 15898 3913
rect 15842 3839 15898 3848
rect 15842 3768 15898 3777
rect 15842 3703 15844 3712
rect 15896 3703 15898 3712
rect 15844 3674 15896 3680
rect 15488 3182 15608 3210
rect 15856 3194 15884 3674
rect 15948 3233 15976 9862
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 7206 16068 7822
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16132 6497 16160 9862
rect 16224 9518 16252 11834
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 7546 16252 8230
rect 16316 7834 16344 15846
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16408 14278 16436 15302
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 12918 16436 14214
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16394 12744 16450 12753
rect 16394 12679 16450 12688
rect 16408 12646 16436 12679
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16394 12200 16450 12209
rect 16394 12135 16450 12144
rect 16408 11665 16436 12135
rect 16500 12084 16528 13330
rect 16592 13326 16620 15302
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14550 16804 14962
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12238 16620 13262
rect 16684 12986 16712 13942
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16764 12640 16816 12646
rect 16762 12608 16764 12617
rect 16816 12608 16818 12617
rect 16762 12543 16818 12552
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16580 12232 16632 12238
rect 16578 12200 16580 12209
rect 16632 12200 16634 12209
rect 16578 12135 16634 12144
rect 16580 12096 16632 12102
rect 16500 12056 16580 12084
rect 16394 11656 16450 11665
rect 16394 11591 16450 11600
rect 16408 10130 16436 11591
rect 16500 11098 16528 12056
rect 16580 12038 16632 12044
rect 16776 11898 16804 12310
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16580 11144 16632 11150
rect 16500 11092 16580 11098
rect 16500 11086 16632 11092
rect 16500 11070 16620 11086
rect 16500 10810 16528 11070
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9450 16436 10066
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 8498 16436 8774
rect 16670 8528 16726 8537
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16580 8492 16632 8498
rect 16670 8463 16726 8472
rect 16580 8434 16632 8440
rect 16592 8022 16620 8434
rect 16684 8430 16712 8463
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16776 8090 16804 11834
rect 16868 9178 16896 16934
rect 16960 14958 16988 19207
rect 17052 16658 17080 20431
rect 17512 20369 17540 27520
rect 24030 27160 24086 27169
rect 24030 27095 24086 27104
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 23662 24440 23718 24449
rect 23662 24375 23718 24384
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 21730 22672 21786 22681
rect 21730 22607 21786 22616
rect 20810 22400 20866 22409
rect 19622 22332 19918 22352
rect 20810 22335 20866 22344
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 18234 20496 18290 20505
rect 18234 20431 18290 20440
rect 17498 20360 17554 20369
rect 17498 20295 17554 20304
rect 18248 18970 18276 20431
rect 19340 20256 19392 20262
rect 19168 20204 19340 20210
rect 19168 20198 19392 20204
rect 19168 20182 19380 20198
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18086 18000 18770
rect 19062 18728 19118 18737
rect 19062 18663 19118 18672
rect 17960 18080 18012 18086
rect 17880 18028 17960 18034
rect 17880 18022 18012 18028
rect 17880 18006 18000 18022
rect 17880 17814 17908 18006
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18432 16794 18460 17002
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17052 16250 17080 16594
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17420 15910 17448 16662
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15366 17448 15846
rect 17972 15638 18000 15914
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17960 15632 18012 15638
rect 17958 15600 17960 15609
rect 18012 15600 18014 15609
rect 17880 15558 17958 15586
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 17408 14816 17460 14822
rect 17512 14804 17540 15438
rect 17880 15162 17908 15558
rect 17958 15535 18014 15544
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17460 14776 17540 14804
rect 17408 14758 17460 14764
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13870 16988 14350
rect 17038 14240 17094 14249
rect 17038 14175 17094 14184
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12442 16988 12582
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16960 11354 16988 12378
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10606 16988 10950
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16316 7806 16436 7834
rect 16302 7712 16358 7721
rect 16302 7647 16358 7656
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16224 7410 16252 7482
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16316 7342 16344 7647
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16118 6488 16174 6497
rect 16118 6423 16174 6432
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16040 3534 16068 4694
rect 16132 4010 16160 4966
rect 16316 4690 16344 5170
rect 16408 5166 16436 7806
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 5817 16528 7142
rect 16592 6866 16620 7958
rect 16776 7478 16804 8026
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 7002 16712 7210
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16486 5808 16542 5817
rect 16486 5743 16542 5752
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5370 16712 5510
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3738 16160 3946
rect 16302 3768 16358 3777
rect 16120 3732 16172 3738
rect 16302 3703 16358 3712
rect 16120 3674 16172 3680
rect 16316 3670 16344 3703
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15934 3224 15990 3233
rect 15580 2666 15608 3182
rect 15844 3188 15896 3194
rect 15934 3159 15990 3168
rect 15844 3130 15896 3136
rect 15842 3088 15898 3097
rect 15842 3023 15898 3032
rect 15396 2638 15608 2666
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15396 480 15424 2638
rect 15474 2408 15530 2417
rect 15474 2343 15476 2352
rect 15528 2343 15530 2352
rect 15476 2314 15528 2320
rect 15856 1714 15884 3023
rect 15934 2680 15990 2689
rect 15934 2615 15936 2624
rect 15988 2615 15990 2624
rect 15936 2586 15988 2592
rect 16316 2514 16344 3606
rect 16408 2553 16436 4966
rect 16684 4758 16712 5306
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16500 4146 16528 4422
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16764 4072 16816 4078
rect 16486 4040 16542 4049
rect 16486 3975 16542 3984
rect 16762 4040 16764 4049
rect 16816 4040 16818 4049
rect 16762 3975 16818 3984
rect 16500 3777 16528 3975
rect 16486 3768 16542 3777
rect 16486 3703 16542 3712
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16578 3088 16634 3097
rect 16776 3058 16804 3334
rect 16868 3194 16896 7890
rect 16960 5409 16988 10542
rect 17052 7002 17080 14175
rect 17236 13870 17264 14418
rect 17224 13864 17276 13870
rect 17222 13832 17224 13841
rect 17276 13832 17278 13841
rect 17222 13767 17278 13776
rect 17222 13424 17278 13433
rect 17222 13359 17278 13368
rect 17130 12200 17186 12209
rect 17130 12135 17186 12144
rect 17144 11898 17172 12135
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17130 11792 17186 11801
rect 17130 11727 17186 11736
rect 17144 11529 17172 11727
rect 17130 11520 17186 11529
rect 17130 11455 17186 11464
rect 17236 11354 17264 13359
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17236 10810 17264 11290
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17052 5914 17080 6938
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16946 5400 17002 5409
rect 16946 5335 17002 5344
rect 16946 5264 17002 5273
rect 16946 5199 17002 5208
rect 16960 4010 16988 5199
rect 17038 4584 17094 4593
rect 17038 4519 17094 4528
rect 17052 4146 17080 4519
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17144 4049 17172 10406
rect 17328 10198 17356 10610
rect 17420 10538 17448 14758
rect 17592 14272 17644 14278
rect 18064 14249 18092 15846
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18248 14618 18276 15438
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 17592 14214 17644 14220
rect 18050 14240 18106 14249
rect 17604 11898 17632 14214
rect 18050 14175 18106 14184
rect 18050 13968 18106 13977
rect 18050 13903 18106 13912
rect 17958 12200 18014 12209
rect 17776 12164 17828 12170
rect 17696 12124 17776 12152
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17512 10198 17540 10678
rect 17604 10470 17632 11154
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17316 10192 17368 10198
rect 17500 10192 17552 10198
rect 17316 10134 17368 10140
rect 17406 10160 17462 10169
rect 17328 9722 17356 10134
rect 17500 10134 17552 10140
rect 17406 10095 17462 10104
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 8974 17356 9318
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 8634 17356 8910
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17420 8265 17448 10095
rect 17406 8256 17462 8265
rect 17406 8191 17462 8200
rect 17222 7576 17278 7585
rect 17222 7511 17278 7520
rect 17236 6934 17264 7511
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17236 6458 17264 6734
rect 17512 6730 17540 10134
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17222 5672 17278 5681
rect 17222 5607 17278 5616
rect 17236 4457 17264 5607
rect 17328 5030 17356 6598
rect 17512 6390 17540 6666
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17604 5681 17632 10406
rect 17696 9110 17724 12124
rect 17958 12135 18014 12144
rect 17776 12106 17828 12112
rect 17774 11928 17830 11937
rect 17774 11863 17776 11872
rect 17828 11863 17830 11872
rect 17776 11834 17828 11840
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10192 17828 10198
rect 17774 10160 17776 10169
rect 17828 10160 17830 10169
rect 17774 10095 17830 10104
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9382 17816 9862
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17774 9208 17830 9217
rect 17880 9178 17908 10406
rect 17972 9586 18000 12135
rect 18064 11354 18092 13903
rect 18144 13864 18196 13870
rect 18248 13818 18276 14350
rect 18340 14346 18368 14758
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18326 14240 18382 14249
rect 18326 14175 18382 14184
rect 18196 13812 18276 13818
rect 18144 13806 18276 13812
rect 18156 13790 18276 13806
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13190 18184 13670
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12850 18184 13126
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18248 12238 18276 13790
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18340 11778 18368 14175
rect 18432 11898 18460 16730
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18616 15910 18644 16526
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18616 14890 18644 15846
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18616 14414 18644 14826
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18510 13288 18566 13297
rect 18510 13223 18566 13232
rect 18524 12986 18552 13223
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18524 12714 18552 12922
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18156 11750 18368 11778
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18064 10606 18092 11290
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17774 9143 17830 9152
rect 17868 9172 17920 9178
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17788 8072 17816 9143
rect 17868 9114 17920 9120
rect 17880 8634 17908 9114
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17696 8044 17816 8072
rect 17590 5672 17646 5681
rect 17590 5607 17646 5616
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4486 17356 4966
rect 17498 4720 17554 4729
rect 17498 4655 17500 4664
rect 17552 4655 17554 4664
rect 17500 4626 17552 4632
rect 17316 4480 17368 4486
rect 17222 4448 17278 4457
rect 17316 4422 17368 4428
rect 17222 4383 17278 4392
rect 17130 4040 17186 4049
rect 16948 4004 17000 4010
rect 17130 3975 17186 3984
rect 16948 3946 17000 3952
rect 17500 3664 17552 3670
rect 17222 3632 17278 3641
rect 17500 3606 17552 3612
rect 17222 3567 17278 3576
rect 17040 3392 17092 3398
rect 17236 3369 17264 3567
rect 17040 3334 17092 3340
rect 17222 3360 17278 3369
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16578 3023 16634 3032
rect 16764 3052 16816 3058
rect 16592 2922 16620 3023
rect 16764 2994 16816 3000
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16592 2650 16620 2858
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16394 2544 16450 2553
rect 16304 2508 16356 2514
rect 16394 2479 16450 2488
rect 16304 2450 16356 2456
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 15856 1686 15976 1714
rect 15948 480 15976 1686
rect 16684 1442 16712 2314
rect 16776 1873 16804 2994
rect 17052 2961 17080 3334
rect 17222 3295 17278 3304
rect 17038 2952 17094 2961
rect 17038 2887 17094 2896
rect 17512 2854 17540 3606
rect 17500 2848 17552 2854
rect 17498 2816 17500 2825
rect 17552 2816 17554 2825
rect 17498 2751 17554 2760
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16868 2310 16896 2450
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16762 1864 16818 1873
rect 16762 1799 16818 1808
rect 16868 1737 16896 2246
rect 16854 1728 16910 1737
rect 16854 1663 16910 1672
rect 16500 1414 16712 1442
rect 17038 1456 17094 1465
rect 16500 480 16528 1414
rect 17038 1391 17094 1400
rect 17052 480 17080 1391
rect 17604 480 17632 5238
rect 17696 4570 17724 8044
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17788 7546 17816 7890
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17788 7274 17816 7482
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17880 5930 17908 8230
rect 17972 6254 18000 8774
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6662 18092 7278
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18064 6089 18092 6598
rect 18050 6080 18106 6089
rect 18050 6015 18106 6024
rect 17880 5902 18092 5930
rect 17866 5672 17922 5681
rect 17866 5607 17922 5616
rect 17774 5128 17830 5137
rect 17774 5063 17776 5072
rect 17828 5063 17830 5072
rect 17776 5034 17828 5040
rect 17880 4826 17908 5607
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17960 4684 18012 4690
rect 17880 4644 17960 4672
rect 17696 4542 17816 4570
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 2145 17724 4422
rect 17788 3602 17816 4542
rect 17880 4146 17908 4644
rect 17960 4626 18012 4632
rect 18064 4570 18092 5902
rect 17972 4542 18092 4570
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17788 3194 17816 3538
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17972 2650 18000 4542
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 2689 18092 3878
rect 18156 3466 18184 11750
rect 18432 11694 18460 11834
rect 18524 11762 18552 12174
rect 18616 12102 18644 12786
rect 18708 12782 18736 15846
rect 18800 15706 18828 16934
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18800 14958 18828 15642
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18892 15026 18920 15302
rect 18970 15056 19026 15065
rect 18880 15020 18932 15026
rect 18970 14991 19026 15000
rect 18880 14962 18932 14968
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18786 14512 18842 14521
rect 18892 14482 18920 14962
rect 18984 14822 19012 14991
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 19076 14657 19104 18663
rect 19062 14648 19118 14657
rect 19062 14583 19118 14592
rect 18786 14447 18842 14456
rect 18880 14476 18932 14482
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18340 11354 18368 11630
rect 18800 11354 18828 14447
rect 18880 14418 18932 14424
rect 18892 13530 18920 14418
rect 19076 13818 19104 14583
rect 18984 13790 19104 13818
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18984 13410 19012 13790
rect 18892 13382 19012 13410
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18340 9625 18368 11154
rect 18708 10674 18736 11154
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18524 10266 18552 10542
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18326 9616 18382 9625
rect 18326 9551 18382 9560
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 18340 9178 18368 9551
rect 18524 9353 18552 9551
rect 18510 9344 18566 9353
rect 18510 9279 18566 9288
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18248 8129 18276 8298
rect 18234 8120 18290 8129
rect 18234 8055 18290 8064
rect 18340 7954 18368 9114
rect 18892 8090 18920 13382
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12889 19012 13126
rect 19064 12912 19116 12918
rect 18970 12880 19026 12889
rect 19064 12854 19116 12860
rect 18970 12815 19026 12824
rect 18970 10976 19026 10985
rect 18970 10911 19026 10920
rect 18984 10198 19012 10911
rect 19076 10606 19104 12854
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 19168 9178 19196 20182
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19982 17640 20038 17649
rect 19982 17575 20038 17584
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16794 20024 17575
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16998 20760 17070
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20732 16697 20760 16934
rect 20718 16688 20774 16697
rect 19708 16652 19760 16658
rect 20718 16623 20774 16632
rect 19708 16594 19760 16600
rect 19720 15978 19748 16594
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20088 16250 20116 16526
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20364 16114 20392 16390
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 19708 15972 19760 15978
rect 19708 15914 19760 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19524 15496 19576 15502
rect 19444 15456 19524 15484
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19260 12442 19288 13466
rect 19352 13462 19380 15030
rect 19444 14822 19472 15456
rect 19524 15438 19576 15444
rect 19628 14890 19656 15506
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19432 14816 19484 14822
rect 19430 14784 19432 14793
rect 19484 14784 19486 14793
rect 19430 14719 19486 14728
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 14006 19472 14418
rect 20088 14278 20116 14826
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19430 13832 19486 13841
rect 19430 13767 19486 13776
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19352 12442 19380 13398
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19352 11937 19380 12242
rect 19444 12238 19472 13767
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20088 13326 20116 14214
rect 20166 13832 20222 13841
rect 20166 13767 20222 13776
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19904 12628 19932 13194
rect 20180 12866 20208 13767
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20272 13530 20300 13670
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 13025 20300 13126
rect 20258 13016 20314 13025
rect 20258 12951 20314 12960
rect 20076 12844 20128 12850
rect 20180 12838 20300 12866
rect 20076 12786 20128 12792
rect 19904 12600 20015 12628
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19987 12424 20015 12600
rect 20088 12442 20116 12786
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 20180 12617 20208 12650
rect 20166 12608 20222 12617
rect 20166 12543 20222 12552
rect 20076 12436 20128 12442
rect 19987 12396 20024 12424
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19524 12232 19576 12238
rect 19996 12209 20024 12396
rect 20076 12378 20128 12384
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19524 12174 19576 12180
rect 19982 12200 20038 12209
rect 19338 11928 19394 11937
rect 19444 11898 19472 12174
rect 19338 11863 19394 11872
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19352 10282 19380 11290
rect 19536 11218 19564 12174
rect 19982 12135 20038 12144
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 10810 19472 11018
rect 19720 10985 19748 11154
rect 19706 10976 19762 10985
rect 19706 10911 19762 10920
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19536 10713 19564 10746
rect 19522 10704 19578 10713
rect 19522 10639 19578 10648
rect 19430 10568 19486 10577
rect 19614 10568 19670 10577
rect 19486 10526 19614 10554
rect 19430 10503 19486 10512
rect 19996 10538 20024 11766
rect 19614 10503 19670 10512
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19260 10266 19380 10282
rect 19248 10260 19380 10266
rect 19300 10254 19380 10260
rect 19248 10202 19300 10208
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9500 19288 9862
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9512 19392 9518
rect 19260 9472 19340 9500
rect 19340 9454 19392 9460
rect 19340 9376 19392 9382
rect 19260 9324 19340 9330
rect 19260 9318 19392 9324
rect 19260 9302 19380 9318
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19076 8362 19104 8774
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7410 18276 7686
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18340 7290 18368 7890
rect 18696 7744 18748 7750
rect 18694 7712 18696 7721
rect 18748 7712 18750 7721
rect 18694 7647 18750 7656
rect 18786 7576 18842 7585
rect 18892 7546 18920 8026
rect 19076 7954 19104 8298
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18786 7511 18842 7520
rect 18880 7540 18932 7546
rect 18248 7262 18368 7290
rect 18248 6934 18276 7262
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 5545 18276 6734
rect 18234 5536 18290 5545
rect 18234 5471 18290 5480
rect 18234 5264 18290 5273
rect 18234 5199 18290 5208
rect 18248 4826 18276 5199
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3738 18276 4014
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18248 3194 18276 3470
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 3058 18276 3130
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18050 2680 18106 2689
rect 17960 2644 18012 2650
rect 18050 2615 18106 2624
rect 18144 2644 18196 2650
rect 17960 2586 18012 2592
rect 18144 2586 18196 2592
rect 18050 2544 18106 2553
rect 18156 2514 18184 2586
rect 18050 2479 18052 2488
rect 18104 2479 18106 2488
rect 18144 2508 18196 2514
rect 18052 2450 18104 2456
rect 18144 2450 18196 2456
rect 18248 2378 18276 2994
rect 18340 2553 18368 7142
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5778 18460 6190
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18432 4486 18460 5714
rect 18524 5574 18552 6122
rect 18694 5944 18750 5953
rect 18694 5879 18750 5888
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 4622 18552 5510
rect 18616 5370 18644 5714
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18616 3738 18644 4082
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18616 3194 18644 3674
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18326 2544 18382 2553
rect 18326 2479 18382 2488
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 17682 2136 17738 2145
rect 17682 2071 17684 2080
rect 17736 2071 17738 2080
rect 17684 2042 17736 2048
rect 17696 2011 17724 2042
rect 18142 2000 18198 2009
rect 18142 1935 18198 1944
rect 18156 480 18184 1935
rect 18708 480 18736 5879
rect 18800 4078 18828 7511
rect 18880 7482 18932 7488
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18892 3670 18920 7346
rect 19076 6866 19104 7890
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19168 5098 19196 8230
rect 19260 7818 19288 9302
rect 19444 9042 19472 9590
rect 19536 9382 19564 9998
rect 19996 9625 20024 9998
rect 19982 9616 20038 9625
rect 19982 9551 20038 9560
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 20088 9330 20116 12242
rect 20180 10266 20208 12378
rect 20272 11354 20300 12838
rect 20364 11540 20392 16050
rect 20456 16046 20484 16390
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15706 20484 15982
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20456 15366 20484 15438
rect 20548 15434 20576 15846
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15201 20484 15302
rect 20442 15192 20498 15201
rect 20442 15127 20498 15136
rect 20626 15192 20682 15201
rect 20626 15127 20682 15136
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 13705 20484 14758
rect 20548 14618 20576 14894
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20534 14376 20590 14385
rect 20534 14311 20590 14320
rect 20548 13734 20576 14311
rect 20536 13728 20588 13734
rect 20442 13696 20498 13705
rect 20536 13670 20588 13676
rect 20442 13631 20498 13640
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20456 12594 20484 13466
rect 20548 13190 20576 13670
rect 20640 13530 20668 15127
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 14414 20760 14554
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20640 12986 20668 13262
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20628 12640 20680 12646
rect 20456 12566 20576 12594
rect 20628 12582 20680 12588
rect 20442 12472 20498 12481
rect 20442 12407 20498 12416
rect 20456 12306 20484 12407
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20548 12186 20576 12566
rect 20456 12158 20576 12186
rect 20456 11830 20484 12158
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20548 11694 20576 12038
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20444 11552 20496 11558
rect 20364 11512 20444 11540
rect 20444 11494 20496 11500
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20456 11150 20484 11494
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 20364 10849 20392 10950
rect 20350 10840 20406 10849
rect 20350 10775 20406 10784
rect 20548 10606 20576 11630
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20180 9722 20208 10202
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20272 9450 20300 9862
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20364 9382 20392 10066
rect 20442 9888 20498 9897
rect 20442 9823 20498 9832
rect 20352 9376 20404 9382
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19338 8256 19394 8265
rect 19338 8191 19394 8200
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19352 7426 19380 8191
rect 19444 8022 19472 8978
rect 19536 8838 19564 9318
rect 20088 9302 20300 9330
rect 20352 9318 20404 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 8430 19564 8774
rect 19904 8673 19932 8910
rect 19890 8664 19946 8673
rect 19890 8599 19892 8608
rect 19944 8599 19946 8608
rect 19892 8570 19944 8576
rect 19904 8539 19932 8570
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19432 7880 19484 7886
rect 19430 7848 19432 7857
rect 19484 7848 19486 7857
rect 19430 7783 19486 7792
rect 19444 7546 19472 7783
rect 19996 7546 20024 8978
rect 20180 8634 20208 9046
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20180 8090 20208 8570
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20074 7576 20130 7585
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19984 7540 20036 7546
rect 20074 7511 20130 7520
rect 19984 7482 20036 7488
rect 19522 7440 19578 7449
rect 19352 7398 19472 7426
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 19340 6860 19392 6866
rect 19260 6730 19288 6831
rect 19340 6802 19392 6808
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19352 6458 19380 6802
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 6186 19472 7398
rect 19522 7375 19578 7384
rect 19536 7002 19564 7375
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20088 7041 20116 7511
rect 20180 7410 20208 8026
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20074 7032 20130 7041
rect 19524 6996 19576 7002
rect 20074 6967 20130 6976
rect 19524 6938 19576 6944
rect 19536 6458 19564 6938
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 20088 6118 20116 6734
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19260 5868 19472 5896
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 18880 3664 18932 3670
rect 18878 3632 18880 3641
rect 18932 3632 18934 3641
rect 18878 3567 18934 3576
rect 18892 2922 18920 3567
rect 19076 3097 19104 4422
rect 19168 4214 19196 4558
rect 19156 4208 19208 4214
rect 19154 4176 19156 4185
rect 19208 4176 19210 4185
rect 19154 4111 19210 4120
rect 19062 3088 19118 3097
rect 19062 3023 19118 3032
rect 19076 2990 19104 3023
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 19260 480 19288 5868
rect 19338 5808 19394 5817
rect 19444 5794 19472 5868
rect 19522 5808 19578 5817
rect 19444 5766 19522 5794
rect 19338 5743 19394 5752
rect 19522 5743 19578 5752
rect 19352 4690 19380 5743
rect 20088 5574 20116 6054
rect 20166 5944 20222 5953
rect 20166 5879 20222 5888
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19430 5400 19486 5409
rect 19430 5335 19486 5344
rect 19444 4758 19472 5335
rect 19720 5137 19748 5510
rect 20088 5166 20116 5510
rect 20076 5160 20128 5166
rect 19706 5128 19762 5137
rect 20076 5102 20128 5108
rect 19706 5063 19762 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20088 4826 20116 5102
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 20180 4146 20208 5879
rect 20272 4214 20300 9302
rect 20364 9081 20392 9318
rect 20350 9072 20406 9081
rect 20350 9007 20406 9016
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 8090 20392 8230
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20350 7848 20406 7857
rect 20350 7783 20352 7792
rect 20404 7783 20406 7792
rect 20352 7754 20404 7760
rect 20364 7206 20392 7754
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20456 6866 20484 9823
rect 20640 9738 20668 12582
rect 20732 12102 20760 14350
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20548 9710 20668 9738
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20548 5846 20576 9710
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20640 9178 20668 9454
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 7426 20760 8774
rect 20640 7398 20760 7426
rect 20640 7342 20668 7398
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 7002 20668 7278
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20824 6458 20852 22335
rect 21744 21146 21772 22607
rect 23202 22536 23258 22545
rect 23202 22471 23258 22480
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21560 20602 21588 20946
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 23216 18306 23244 22471
rect 23480 22432 23532 22438
rect 23478 22400 23480 22409
rect 23532 22400 23534 22409
rect 23478 22335 23534 22344
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23124 18278 23244 18306
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 21270 17776 21326 17785
rect 21270 17711 21326 17720
rect 21824 17740 21876 17746
rect 21284 17678 21312 17711
rect 21824 17682 21876 17688
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21836 16998 21864 17682
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21008 16833 21036 16934
rect 20994 16824 21050 16833
rect 20994 16759 21050 16768
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21284 15366 21312 16458
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21178 14920 21234 14929
rect 21178 14855 21234 14864
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20902 12880 20958 12889
rect 20902 12815 20958 12824
rect 20916 12306 20944 12815
rect 21008 12322 21036 13738
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21100 12986 21128 13262
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21192 12442 21220 14855
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 20904 12300 20956 12306
rect 21008 12294 21220 12322
rect 20904 12242 20956 12248
rect 20916 11354 20944 12242
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 21008 11286 21036 12174
rect 21100 12073 21128 12174
rect 21086 12064 21142 12073
rect 21086 11999 21142 12008
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21100 10810 21128 11562
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21192 10130 21220 12294
rect 21284 11558 21312 15302
rect 21376 15162 21404 16050
rect 21468 15366 21496 16662
rect 21730 16008 21786 16017
rect 21730 15943 21732 15952
rect 21784 15943 21786 15952
rect 21732 15914 21784 15920
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21376 14550 21404 15098
rect 21364 14544 21416 14550
rect 21468 14521 21496 15302
rect 21546 14920 21602 14929
rect 21546 14855 21548 14864
rect 21600 14855 21602 14864
rect 21548 14826 21600 14832
rect 21364 14486 21416 14492
rect 21454 14512 21510 14521
rect 21376 14074 21404 14486
rect 21454 14447 21510 14456
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21376 13530 21404 13738
rect 21652 13530 21680 15846
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21744 13734 21772 15302
rect 21836 14074 21864 16934
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21928 14958 21956 16730
rect 22020 16590 22048 17138
rect 22480 17066 22508 17682
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22020 16182 22048 16390
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22020 15473 22048 15982
rect 22098 15872 22154 15881
rect 22098 15807 22154 15816
rect 22112 15502 22140 15807
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22100 15496 22152 15502
rect 22006 15464 22062 15473
rect 22100 15438 22152 15444
rect 22006 15399 22062 15408
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 22112 14890 22140 15438
rect 22204 15162 22232 15574
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22296 15042 22324 17002
rect 22480 16969 22508 17002
rect 22560 16992 22612 16998
rect 22466 16960 22522 16969
rect 22560 16934 22612 16940
rect 22466 16895 22522 16904
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 15706 22508 16390
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22572 15638 22600 16934
rect 22836 16720 22888 16726
rect 22650 16688 22706 16697
rect 22836 16662 22888 16668
rect 22650 16623 22706 16632
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 15162 22416 15438
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22204 15014 22324 15042
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21560 12986 21588 13330
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21652 12442 21680 13466
rect 21744 13190 21772 13670
rect 21928 13326 21956 14214
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21744 10470 21772 11290
rect 21822 11112 21878 11121
rect 21822 11047 21824 11056
rect 21876 11047 21878 11056
rect 21824 11018 21876 11024
rect 21928 10554 21956 12718
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21836 10526 21956 10554
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 10169 21772 10406
rect 21730 10160 21786 10169
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21364 10124 21416 10130
rect 21730 10095 21786 10104
rect 21364 10066 21416 10072
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20916 9178 20944 9522
rect 21284 9382 21312 9998
rect 21376 9382 21404 10066
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20916 8362 20944 9114
rect 21284 8945 21312 9318
rect 21270 8936 21326 8945
rect 21270 8871 21326 8880
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20916 7857 20944 7890
rect 20902 7848 20958 7857
rect 20902 7783 20958 7792
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6905 20944 7142
rect 20902 6896 20958 6905
rect 20902 6831 20958 6840
rect 20996 6860 21048 6866
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20640 5370 20668 6326
rect 20916 6254 20944 6831
rect 21100 6848 21128 8366
rect 21048 6820 21128 6848
rect 20996 6802 21048 6808
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20720 4480 20772 4486
rect 20640 4440 20720 4468
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 19432 3936 19484 3942
rect 19430 3904 19432 3913
rect 19484 3904 19486 3913
rect 19430 3839 19486 3848
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19430 3768 19486 3777
rect 19622 3760 19918 3780
rect 19486 3726 19564 3754
rect 19430 3703 19486 3712
rect 19536 3618 19564 3726
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19536 3590 19748 3618
rect 19720 3505 19748 3590
rect 19892 3528 19944 3534
rect 19522 3496 19578 3505
rect 19522 3431 19578 3440
rect 19706 3496 19762 3505
rect 19892 3470 19944 3476
rect 19706 3431 19762 3440
rect 19536 2530 19564 3431
rect 19904 3194 19932 3470
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2650 20024 3674
rect 20258 3632 20314 3641
rect 20258 3567 20314 3576
rect 20272 3369 20300 3567
rect 20258 3360 20314 3369
rect 20258 3295 20314 3304
rect 20456 3126 20484 4082
rect 20640 3738 20668 4440
rect 20720 4422 20772 4428
rect 20824 4146 20852 4490
rect 21008 4146 21036 6802
rect 21376 6769 21404 9318
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 7750 21496 8910
rect 21546 8664 21602 8673
rect 21546 8599 21602 8608
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21362 6760 21418 6769
rect 21362 6695 21418 6704
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21284 6322 21312 6598
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5914 21312 6258
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21284 5681 21312 5714
rect 21364 5704 21416 5710
rect 21270 5672 21326 5681
rect 21364 5646 21416 5652
rect 21270 5607 21326 5616
rect 21376 5370 21404 5646
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20810 4040 20866 4049
rect 20810 3975 20866 3984
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19536 2502 19840 2530
rect 19812 480 19840 2502
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 1465 20208 2246
rect 20166 1456 20222 1465
rect 20166 1391 20222 1400
rect 20364 480 20392 2790
rect 20548 2650 20576 3334
rect 20732 3097 20760 3334
rect 20718 3088 20774 3097
rect 20718 3023 20774 3032
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20534 2544 20590 2553
rect 20534 2479 20536 2488
rect 20588 2479 20590 2488
rect 20536 2450 20588 2456
rect 20824 2394 20852 3975
rect 21008 3602 21036 4082
rect 21192 3738 21220 4558
rect 21284 3738 21312 4626
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20916 2582 20944 2926
rect 21008 2922 21036 3538
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20824 2366 20944 2394
rect 20916 480 20944 2366
rect 21468 2281 21496 7686
rect 21560 6866 21588 8599
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21560 6458 21588 6802
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21546 6216 21602 6225
rect 21546 6151 21602 6160
rect 21560 5681 21588 6151
rect 21652 6089 21680 9862
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 8634 21772 9046
rect 21836 8974 21864 10526
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 9489 21956 10406
rect 22020 10266 22048 12582
rect 22112 11354 22140 14486
rect 22204 13954 22232 15014
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14618 22324 14894
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22388 14346 22416 15098
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22388 14074 22416 14282
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22204 13926 22416 13954
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22204 12442 22232 12582
rect 22296 12442 22324 13194
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22204 12186 22232 12378
rect 22388 12306 22416 13926
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22204 12158 22416 12186
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22204 10266 22232 11154
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22020 9500 22048 10202
rect 22204 10033 22232 10202
rect 22190 10024 22246 10033
rect 22190 9959 22246 9968
rect 22100 9512 22152 9518
rect 21914 9480 21970 9489
rect 22020 9472 22100 9500
rect 22100 9454 22152 9460
rect 21914 9415 21970 9424
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22190 9344 22246 9353
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21730 6896 21786 6905
rect 21730 6831 21786 6840
rect 21638 6080 21694 6089
rect 21638 6015 21694 6024
rect 21546 5672 21602 5681
rect 21546 5607 21602 5616
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21560 2553 21588 3674
rect 21546 2544 21602 2553
rect 21546 2479 21602 2488
rect 21744 2394 21772 6831
rect 21836 6633 21864 7686
rect 21928 7546 21956 7822
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21822 6624 21878 6633
rect 21822 6559 21878 6568
rect 22020 6497 22048 9318
rect 22190 9279 22246 9288
rect 22098 8664 22154 8673
rect 22098 8599 22100 8608
rect 22152 8599 22154 8608
rect 22100 8570 22152 8576
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6866 22140 7142
rect 22204 6882 22232 9279
rect 22296 8090 22324 12038
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22296 7002 22324 8026
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22100 6860 22152 6866
rect 22204 6854 22324 6882
rect 22100 6802 22152 6808
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21822 6488 21878 6497
rect 21822 6423 21878 6432
rect 22006 6488 22062 6497
rect 22006 6423 22062 6432
rect 21836 6225 21864 6423
rect 21822 6216 21878 6225
rect 21822 6151 21878 6160
rect 22112 5234 22140 6598
rect 22190 6352 22246 6361
rect 22190 6287 22192 6296
rect 22244 6287 22246 6296
rect 22192 6258 22244 6264
rect 22100 5228 22152 5234
rect 22020 5188 22100 5216
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21928 5001 21956 5102
rect 21914 4992 21970 5001
rect 21914 4927 21970 4936
rect 21914 4856 21970 4865
rect 22020 4826 22048 5188
rect 22100 5170 22152 5176
rect 22112 5105 22140 5170
rect 21914 4791 21970 4800
rect 22008 4820 22060 4826
rect 21928 4758 21956 4791
rect 22008 4762 22060 4768
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 22020 4185 22048 4762
rect 22006 4176 22062 4185
rect 22006 4111 22062 4120
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22020 3194 22048 3946
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22098 3224 22154 3233
rect 22008 3188 22060 3194
rect 22204 3194 22232 3606
rect 22098 3159 22154 3168
rect 22192 3188 22244 3194
rect 22008 3130 22060 3136
rect 21560 2366 21772 2394
rect 21454 2272 21510 2281
rect 21454 2207 21510 2216
rect 21560 480 21588 2366
rect 22112 480 22140 3159
rect 22192 3130 22244 3136
rect 22296 2530 22324 6854
rect 22388 5778 22416 12158
rect 22480 11286 22508 15302
rect 22664 14550 22692 16623
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22756 16182 22784 16526
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22756 15638 22784 16118
rect 22848 16046 22876 16662
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22940 16250 22968 16594
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22744 15632 22796 15638
rect 22744 15574 22796 15580
rect 22742 14784 22798 14793
rect 22742 14719 22798 14728
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22664 12850 22692 13466
rect 22652 12844 22704 12850
rect 22572 12804 22652 12832
rect 22572 12374 22600 12804
rect 22652 12786 22704 12792
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22572 11642 22600 12174
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22664 11898 22692 12106
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22572 11614 22692 11642
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22480 10674 22508 11086
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22480 10130 22508 10610
rect 22572 10146 22600 11494
rect 22664 11218 22692 11614
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22664 10470 22692 11154
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 10266 22692 10406
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22468 10124 22520 10130
rect 22572 10118 22692 10146
rect 22468 10066 22520 10072
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22480 8362 22508 9318
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 5914 22508 7142
rect 22572 6361 22600 9318
rect 22558 6352 22614 6361
rect 22558 6287 22614 6296
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22572 5817 22600 6054
rect 22558 5808 22614 5817
rect 22376 5772 22428 5778
rect 22558 5743 22614 5752
rect 22376 5714 22428 5720
rect 22558 5400 22614 5409
rect 22558 5335 22614 5344
rect 22572 5001 22600 5335
rect 22558 4992 22614 5001
rect 22558 4927 22614 4936
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22388 3777 22416 4490
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22374 3768 22430 3777
rect 22374 3703 22430 3712
rect 22480 2650 22508 4422
rect 22664 3670 22692 10118
rect 22756 8090 22784 14719
rect 22940 14600 22968 16186
rect 22848 14572 22968 14600
rect 22848 12238 22876 14572
rect 23032 14521 23060 18022
rect 23018 14512 23074 14521
rect 23018 14447 23074 14456
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23032 13258 23060 14350
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 22926 13152 22982 13161
rect 22926 13087 22982 13096
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22848 11354 22876 12038
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22834 11112 22890 11121
rect 22834 11047 22890 11056
rect 22848 10538 22876 11047
rect 22940 10577 22968 13087
rect 23018 12608 23074 12617
rect 23018 12543 23074 12552
rect 23032 12306 23060 12543
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11558 23060 12242
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22926 10568 22982 10577
rect 22836 10532 22888 10538
rect 22926 10503 22982 10512
rect 22836 10474 22888 10480
rect 22940 10198 22968 10503
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22848 9761 22876 9862
rect 22834 9752 22890 9761
rect 22834 9687 22890 9696
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22848 8974 22876 9522
rect 22940 9178 22968 10134
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23032 9058 23060 11494
rect 22940 9030 23060 9058
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22848 8838 22876 8910
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8294 22876 8774
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22940 8106 22968 9030
rect 23124 8378 23152 18278
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 14550 23244 18022
rect 23204 14544 23256 14550
rect 23204 14486 23256 14492
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22848 8078 22968 8106
rect 23032 8350 23152 8378
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22756 5370 22784 5714
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22756 5030 22784 5306
rect 22744 5024 22796 5030
rect 22742 4992 22744 5001
rect 22796 4992 22798 5001
rect 22742 4927 22798 4936
rect 22848 4049 22876 8078
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5234 22968 5714
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23032 4826 23060 8350
rect 23216 8242 23244 13942
rect 23308 12628 23336 18702
rect 23492 18086 23520 18770
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23492 17898 23520 18022
rect 23400 17870 23520 17898
rect 23400 15026 23428 17870
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 16561 23520 17478
rect 23584 17066 23612 17682
rect 23676 17626 23704 24375
rect 23938 22128 23994 22137
rect 23938 22063 23994 22072
rect 23952 18902 23980 22063
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 24044 18714 24072 27095
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24136 23662 24164 25162
rect 24228 23866 24256 27639
rect 24490 27520 24546 28000
rect 24504 25226 24532 27520
rect 25410 26616 25466 26625
rect 25410 26551 25466 26560
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24766 24984 24822 24993
rect 24766 24919 24822 24928
rect 24780 24018 24808 24919
rect 24780 23990 24900 24018
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24766 23896 24822 23905
rect 24216 23860 24268 23866
rect 24766 23831 24822 23840
rect 24216 23802 24268 23808
rect 24124 23656 24176 23662
rect 24124 23598 24176 23604
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 24780 22794 24808 23831
rect 24872 23322 24900 23990
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 25134 23216 25190 23225
rect 25134 23151 25190 23160
rect 24780 22778 24900 22794
rect 24676 22772 24728 22778
rect 24780 22772 24912 22778
rect 24780 22766 24860 22772
rect 24676 22714 24728 22720
rect 24860 22714 24912 22720
rect 24952 22568 25004 22574
rect 24950 22536 24952 22545
rect 25004 22536 25006 22545
rect 24950 22471 25006 22480
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24766 21584 24822 21593
rect 24766 21519 24822 21528
rect 24674 21040 24730 21049
rect 24674 20975 24730 20984
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24122 19952 24178 19961
rect 24122 19887 24178 19896
rect 24216 19916 24268 19922
rect 23952 18686 24072 18714
rect 23676 17598 23796 17626
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23676 17105 23704 17478
rect 23768 17338 23796 17598
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23662 17096 23718 17105
rect 23572 17060 23624 17066
rect 23662 17031 23718 17040
rect 23572 17002 23624 17008
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23478 16552 23534 16561
rect 23478 16487 23534 16496
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23492 14906 23520 15914
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15502 23612 15846
rect 23676 15570 23704 16759
rect 23754 16008 23810 16017
rect 23754 15943 23810 15952
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23400 14878 23520 14906
rect 23400 14498 23428 14878
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 14657 23520 14758
rect 23478 14648 23534 14657
rect 23584 14618 23612 15438
rect 23676 14958 23704 15506
rect 23664 14952 23716 14958
rect 23768 14929 23796 15943
rect 23860 15586 23888 17206
rect 23952 16794 23980 18686
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23952 16114 23980 16730
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 24044 16017 24072 18566
rect 24136 18426 24164 19887
rect 24216 19858 24268 19864
rect 24228 19394 24256 19858
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24228 19366 24440 19394
rect 24412 19174 24440 19366
rect 24584 19304 24636 19310
rect 24582 19272 24584 19281
rect 24636 19272 24638 19281
rect 24582 19207 24638 19216
rect 24688 19174 24716 20975
rect 24780 20058 24808 21519
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24766 19408 24822 19417
rect 24766 19343 24822 19352
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 24228 18086 24256 18770
rect 24412 18737 24440 19110
rect 24398 18728 24454 18737
rect 24780 18714 24808 19343
rect 24398 18663 24454 18672
rect 24688 18686 24808 18714
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24582 18320 24638 18329
rect 24582 18255 24638 18264
rect 24596 18222 24624 18255
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24228 16726 24256 18022
rect 24688 17882 24716 18686
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 18193 24808 18566
rect 24766 18184 24822 18193
rect 24766 18119 24822 18128
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17270 24716 17682
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24216 16720 24268 16726
rect 24504 16697 24532 17070
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24216 16662 24268 16668
rect 24490 16688 24546 16697
rect 24490 16623 24546 16632
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24124 16108 24176 16114
rect 24176 16068 24256 16096
rect 24124 16050 24176 16056
rect 24030 16008 24086 16017
rect 24030 15943 24086 15952
rect 24124 15972 24176 15978
rect 24124 15914 24176 15920
rect 23860 15558 23980 15586
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23860 15201 23888 15438
rect 23846 15192 23902 15201
rect 23846 15127 23902 15136
rect 23860 15026 23888 15127
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23664 14894 23716 14900
rect 23754 14920 23810 14929
rect 23754 14855 23810 14864
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23478 14583 23534 14592
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23400 14470 23612 14498
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13938 23428 14214
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 13462 23428 13874
rect 23584 13818 23612 14470
rect 23676 13841 23704 14758
rect 23952 14600 23980 15558
rect 23768 14572 23980 14600
rect 23492 13790 23612 13818
rect 23662 13832 23718 13841
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23400 12986 23428 13398
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23388 12776 23440 12782
rect 23492 12764 23520 13790
rect 23662 13767 23718 13776
rect 23440 12736 23520 12764
rect 23768 12730 23796 14572
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23860 13569 23888 13670
rect 23846 13560 23902 13569
rect 23846 13495 23902 13504
rect 23388 12718 23440 12724
rect 23584 12702 23796 12730
rect 23308 12600 23520 12628
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23294 12336 23350 12345
rect 23294 12271 23350 12280
rect 23308 10452 23336 12271
rect 23400 11762 23428 12378
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23492 11354 23520 12600
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23492 10810 23520 11290
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23584 10674 23612 12702
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12481 23704 12582
rect 23662 12472 23718 12481
rect 23662 12407 23718 12416
rect 23662 12336 23718 12345
rect 23662 12271 23718 12280
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23308 10424 23520 10452
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23308 9450 23336 10202
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23400 9330 23428 9454
rect 23308 9302 23428 9330
rect 23308 8498 23336 9302
rect 23492 9217 23520 10424
rect 23478 9208 23534 9217
rect 23478 9143 23534 9152
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23124 8214 23244 8242
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23124 8022 23152 8214
rect 23112 8016 23164 8022
rect 23112 7958 23164 7964
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 6866 23244 7890
rect 23308 7750 23336 8230
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7426 23336 7686
rect 23400 7546 23428 8774
rect 23492 8430 23520 8978
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23308 7398 23428 7426
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23124 5370 23152 5646
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23032 4282 23060 4762
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23124 4146 23152 5306
rect 23308 5166 23336 7210
rect 23400 6866 23428 7398
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23400 6118 23428 6802
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23388 5568 23440 5574
rect 23492 5545 23520 8366
rect 23584 5710 23612 10474
rect 23676 8537 23704 12271
rect 23952 11234 23980 14418
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24044 13530 24072 13874
rect 24136 13802 24164 15914
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 12850 24164 13126
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 24044 11354 24072 12582
rect 24136 12306 24164 12786
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24136 11354 24164 12242
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 23952 11206 24164 11234
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 23662 8528 23718 8537
rect 23662 8463 23718 8472
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23676 6458 23704 7822
rect 23768 6769 23796 11018
rect 23952 10266 23980 11086
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 23952 9722 23980 10066
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 23846 9480 23902 9489
rect 23846 9415 23902 9424
rect 23940 9444 23992 9450
rect 23860 9178 23888 9415
rect 23940 9386 23992 9392
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23754 6760 23810 6769
rect 23754 6695 23810 6704
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23754 6352 23810 6361
rect 23754 6287 23810 6296
rect 23662 6080 23718 6089
rect 23662 6015 23718 6024
rect 23676 5846 23704 6015
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23664 5568 23716 5574
rect 23388 5510 23440 5516
rect 23478 5536 23534 5545
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22834 4040 22890 4049
rect 22834 3975 22890 3984
rect 22742 3904 22798 3913
rect 22742 3839 22798 3848
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22756 3398 22784 3839
rect 23018 3496 23074 3505
rect 23124 3466 23152 4082
rect 23216 3942 23244 4626
rect 23308 4010 23336 5102
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23018 3431 23074 3440
rect 23112 3460 23164 3466
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22756 3194 22784 3334
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 23032 2530 23060 3431
rect 23112 3402 23164 3408
rect 23124 3058 23152 3402
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23216 2689 23244 3878
rect 23400 3754 23428 5510
rect 23664 5510 23716 5516
rect 23478 5471 23534 5480
rect 23478 5400 23534 5409
rect 23478 5335 23534 5344
rect 23492 4826 23520 5335
rect 23676 5302 23704 5510
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23492 4457 23520 4626
rect 23478 4448 23534 4457
rect 23478 4383 23534 4392
rect 23492 4282 23520 4383
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23676 4078 23704 4762
rect 23768 4729 23796 6287
rect 23754 4720 23810 4729
rect 23754 4655 23810 4664
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23400 3726 23520 3754
rect 23492 3670 23520 3726
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23570 3632 23626 3641
rect 23676 3602 23704 3878
rect 23570 3567 23626 3576
rect 23664 3596 23716 3602
rect 23202 2680 23258 2689
rect 23202 2615 23258 2624
rect 22296 2502 22692 2530
rect 23032 2502 23244 2530
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 2145 22600 2246
rect 22558 2136 22614 2145
rect 22558 2071 22614 2080
rect 22664 480 22692 2502
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23032 1737 23060 2246
rect 23018 1728 23074 1737
rect 23018 1663 23074 1672
rect 23216 480 23244 2502
rect 23478 2408 23534 2417
rect 23478 2343 23480 2352
rect 23532 2343 23534 2352
rect 23480 2314 23532 2320
rect 23478 2272 23534 2281
rect 23478 2207 23534 2216
rect 23492 921 23520 2207
rect 23584 1442 23612 3567
rect 23664 3538 23716 3544
rect 23676 3194 23704 3538
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23768 2310 23796 2450
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23768 1601 23796 2246
rect 23860 2009 23888 8774
rect 23952 8634 23980 9386
rect 24044 8838 24072 9658
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23952 7886 23980 8570
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7546 23980 7822
rect 24044 7546 24072 8230
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24136 7426 24164 11206
rect 24228 10690 24256 16068
rect 24688 15638 24716 16594
rect 24676 15632 24728 15638
rect 24674 15600 24676 15609
rect 24728 15600 24730 15609
rect 24674 15535 24730 15544
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24780 15094 24808 17002
rect 24950 16960 25006 16969
rect 24950 16895 25006 16904
rect 24964 15638 24992 16895
rect 25044 15904 25096 15910
rect 25042 15872 25044 15881
rect 25096 15872 25098 15881
rect 25042 15807 25098 15816
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 25056 14278 25084 15506
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 25056 13977 25084 14214
rect 25042 13968 25098 13977
rect 25042 13903 25098 13912
rect 24766 13696 24822 13705
rect 24822 13654 24900 13682
rect 24766 13631 24822 13640
rect 24674 13152 24730 13161
rect 24289 13084 24585 13104
rect 24674 13087 24730 13096
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12782 24716 13087
rect 24872 12850 24900 13654
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24964 12374 24992 13126
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 24320 11150 24348 11562
rect 24766 11248 24822 11257
rect 24766 11183 24822 11192
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24228 10662 24348 10690
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24228 10266 24256 10474
rect 24320 10266 24348 10662
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24780 10169 24808 11183
rect 24766 10160 24822 10169
rect 24872 10130 24900 11834
rect 24964 11286 24992 12310
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 24964 10606 24992 11222
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24766 10095 24822 10104
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 24768 9920 24820 9926
rect 24820 9880 24900 9908
rect 24768 9862 24820 9868
rect 24219 9704 24247 9862
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24676 9716 24728 9722
rect 24219 9676 24256 9704
rect 24228 9602 24256 9676
rect 24676 9658 24728 9664
rect 24228 9574 24348 9602
rect 24320 8906 24348 9574
rect 24688 9194 24716 9658
rect 24872 9586 24900 9880
rect 24964 9654 24992 9998
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24688 9178 24900 9194
rect 24688 9172 24912 9178
rect 24688 9166 24860 9172
rect 24216 8900 24268 8906
rect 24216 8842 24268 8848
rect 24308 8900 24360 8906
rect 24308 8842 24360 8848
rect 24228 8362 24256 8842
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24228 7478 24256 8298
rect 24688 8090 24716 9166
rect 24860 9114 24912 9120
rect 24766 9072 24822 9081
rect 25056 9042 25084 10950
rect 25148 9178 25176 23151
rect 25320 18896 25372 18902
rect 25320 18838 25372 18844
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25240 14793 25268 14894
rect 25226 14784 25282 14793
rect 25226 14719 25282 14728
rect 25332 13512 25360 18838
rect 25424 16250 25452 26551
rect 25502 26072 25558 26081
rect 25502 26007 25558 26016
rect 25516 16794 25544 26007
rect 25870 25528 25926 25537
rect 25870 25463 25926 25472
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25792 15910 25820 16594
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25792 15065 25820 15846
rect 25778 15056 25834 15065
rect 25778 14991 25834 15000
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25332 13484 25452 13512
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25332 13297 25360 13330
rect 25318 13288 25374 13297
rect 25318 13223 25374 13232
rect 25332 12986 25360 13223
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25240 11694 25268 12038
rect 25320 11824 25372 11830
rect 25318 11792 25320 11801
rect 25372 11792 25374 11801
rect 25318 11727 25374 11736
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25424 11354 25452 13484
rect 25792 13410 25820 13670
rect 25884 13530 25912 25463
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25792 13382 25912 13410
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25700 11286 25728 11494
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25502 11112 25558 11121
rect 25502 11047 25558 11056
rect 25318 10568 25374 10577
rect 25318 10503 25374 10512
rect 25332 10470 25360 10503
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25240 9722 25268 10202
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 24766 9007 24822 9016
rect 25044 9036 25096 9042
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23952 7398 24164 7426
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 23952 5273 23980 7398
rect 24124 6724 24176 6730
rect 24124 6666 24176 6672
rect 24030 6624 24086 6633
rect 24030 6559 24086 6568
rect 24044 6254 24072 6559
rect 24136 6497 24164 6666
rect 24228 6662 24256 7414
rect 24688 7410 24716 8026
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24216 6656 24268 6662
rect 24216 6598 24268 6604
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24122 6488 24178 6497
rect 24289 6480 24585 6500
rect 24122 6423 24178 6432
rect 24136 6322 24164 6423
rect 24688 6322 24716 6598
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 24044 5930 24072 6190
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24044 5914 24164 5930
rect 24044 5908 24176 5914
rect 24044 5902 24124 5908
rect 24124 5850 24176 5856
rect 24688 5710 24716 6054
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 23938 5264 23994 5273
rect 23938 5199 23994 5208
rect 24582 5128 24638 5137
rect 24582 5063 24638 5072
rect 23938 4992 23994 5001
rect 23938 4927 23994 4936
rect 23846 2000 23902 2009
rect 23846 1935 23902 1944
rect 23952 1601 23980 4927
rect 24596 4622 24624 5063
rect 24780 5030 24808 9007
rect 25044 8978 25096 8984
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24872 7274 24900 8842
rect 25056 8498 25084 8978
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25516 8106 25544 11047
rect 25608 10470 25636 11154
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 10033 25636 10406
rect 25792 10266 25820 13194
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25594 10024 25650 10033
rect 25594 9959 25650 9968
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25608 9518 25636 9862
rect 25792 9722 25820 10202
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25596 9512 25648 9518
rect 25596 9454 25648 9460
rect 25608 9178 25636 9454
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25608 8242 25636 9114
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25700 8634 25728 9046
rect 25884 8974 25912 13382
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25700 8294 25728 8325
rect 25688 8288 25740 8294
rect 25608 8236 25688 8242
rect 25608 8230 25740 8236
rect 25608 8214 25728 8230
rect 25516 8078 25636 8106
rect 25700 8090 25728 8214
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 25148 6905 25176 7686
rect 25516 7206 25544 7890
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25134 6896 25190 6905
rect 25134 6831 25190 6840
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25042 6760 25098 6769
rect 25042 6695 25098 6704
rect 25056 6458 25084 6695
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25056 6254 25084 6394
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 25148 5914 25176 6598
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24872 4826 24900 5782
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24964 5370 24992 5646
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24674 4720 24730 4729
rect 24674 4655 24730 4664
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24032 4480 24084 4486
rect 24032 4422 24084 4428
rect 24044 2961 24072 4422
rect 24136 4321 24164 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24122 4312 24178 4321
rect 24289 4304 24585 4324
rect 24688 4321 24716 4655
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24674 4312 24730 4321
rect 24122 4247 24124 4256
rect 24176 4247 24178 4256
rect 24674 4247 24730 4256
rect 24124 4218 24176 4224
rect 24136 4187 24164 4218
rect 24872 4146 24900 4558
rect 24950 4176 25006 4185
rect 24860 4140 24912 4146
rect 24950 4111 25006 4120
rect 24860 4082 24912 4088
rect 24308 4072 24360 4078
rect 24122 4040 24178 4049
rect 24964 4026 24992 4111
rect 24308 4014 24360 4020
rect 24122 3975 24178 3984
rect 24136 3942 24164 3975
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 24136 3398 24164 3878
rect 24320 3641 24348 4014
rect 24872 3998 24992 4026
rect 24582 3768 24638 3777
rect 24582 3703 24638 3712
rect 24306 3632 24362 3641
rect 24306 3567 24362 3576
rect 24596 3534 24624 3703
rect 24584 3528 24636 3534
rect 24636 3476 24716 3482
rect 24584 3470 24716 3476
rect 24596 3454 24716 3470
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3454
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24030 2952 24086 2961
rect 24030 2887 24086 2896
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24044 2553 24072 2586
rect 24780 2553 24808 3334
rect 24030 2544 24086 2553
rect 24030 2479 24086 2488
rect 24766 2544 24822 2553
rect 24766 2479 24822 2488
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23754 1592 23810 1601
rect 23754 1527 23810 1536
rect 23938 1592 23994 1601
rect 23938 1527 23994 1536
rect 23584 1414 23796 1442
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 23768 480 23796 1414
rect 24228 598 24348 626
rect 4618 96 4674 105
rect 4618 31 4674 40
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18694 0 18750 480
rect 19246 0 19302 480
rect 19798 0 19854 480
rect 20350 0 20406 480
rect 20902 0 20958 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24228 105 24256 598
rect 24320 480 24348 598
rect 24872 480 24900 3998
rect 25148 3913 25176 5850
rect 25134 3904 25190 3913
rect 25134 3839 25190 3848
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24964 2650 24992 3130
rect 25240 2854 25268 6598
rect 25332 6089 25360 6802
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25424 6225 25452 6258
rect 25410 6216 25466 6225
rect 25410 6151 25466 6160
rect 25318 6080 25374 6089
rect 25318 6015 25374 6024
rect 25412 5636 25464 5642
rect 25412 5578 25464 5584
rect 25424 5370 25452 5578
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24964 2446 24992 2586
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 25424 480 25452 4966
rect 25516 4146 25544 7142
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25608 4078 25636 8078
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25700 6458 25728 8026
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25700 5914 25728 6394
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25700 5386 25728 5850
rect 25700 5370 25820 5386
rect 25700 5364 25832 5370
rect 25700 5358 25780 5364
rect 25700 5166 25728 5358
rect 25780 5306 25832 5312
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25700 4826 25728 5102
rect 25688 4820 25740 4826
rect 25688 4762 25740 4768
rect 25700 4146 25728 4762
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25596 4072 25648 4078
rect 25596 4014 25648 4020
rect 25700 3754 25728 4082
rect 25608 3738 25728 3754
rect 25596 3732 25728 3738
rect 25648 3726 25728 3732
rect 25596 3674 25648 3680
rect 25608 3126 25636 3674
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25700 3194 25728 3606
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25596 3120 25648 3126
rect 25884 3097 25912 8910
rect 25962 7848 26018 7857
rect 25962 7783 26018 7792
rect 25976 7546 26004 7783
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 26148 7268 26200 7274
rect 26148 7210 26200 7216
rect 25964 6112 26016 6118
rect 25962 6080 25964 6089
rect 26016 6080 26018 6089
rect 25962 6015 26018 6024
rect 26160 5778 26188 7210
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 25962 5672 26018 5681
rect 25962 5607 26018 5616
rect 25596 3062 25648 3068
rect 25870 3088 25926 3097
rect 25608 2922 25636 3062
rect 25870 3023 25926 3032
rect 25596 2916 25648 2922
rect 25596 2858 25648 2864
rect 25594 2680 25650 2689
rect 25594 2615 25596 2624
rect 25648 2615 25650 2624
rect 25596 2586 25648 2592
rect 25976 480 26004 5607
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 26068 2582 26096 3062
rect 26056 2576 26108 2582
rect 26056 2518 26108 2524
rect 24214 96 24270 105
rect 24214 31 24270 40
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26160 377 26188 5714
rect 26528 480 26556 6122
rect 27618 1728 27674 1737
rect 27618 1663 27674 1672
rect 26790 1456 26846 1465
rect 26846 1414 27108 1442
rect 26790 1391 26846 1400
rect 27080 480 27108 1414
rect 27632 480 27660 1663
rect 26146 368 26202 377
rect 26146 303 26202 312
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3422 27648 3478 27704
rect 2686 26560 2742 26616
rect 1582 24248 1638 24304
rect 1490 23160 1546 23216
rect 2594 22480 2650 22536
rect 2042 22380 2044 22400
rect 2044 22380 2096 22400
rect 2096 22380 2098 22400
rect 2042 22344 2098 22380
rect 1490 21392 1546 21448
rect 1582 20848 1638 20904
rect 1490 20304 1546 20360
rect 1398 19624 1454 19680
rect 2042 20204 2044 20224
rect 2044 20204 2096 20224
rect 2096 20204 2098 20224
rect 2042 20168 2098 20204
rect 2410 19116 2412 19136
rect 2412 19116 2464 19136
rect 2464 19116 2466 19136
rect 2410 19080 2466 19116
rect 1582 18572 1584 18592
rect 1584 18572 1636 18592
rect 1636 18572 1638 18592
rect 1582 18536 1638 18572
rect 2042 16532 2044 16552
rect 2044 16532 2096 16552
rect 2096 16532 2098 16552
rect 2042 16496 2098 16532
rect 1858 15408 1914 15464
rect 1950 13776 2006 13832
rect 1766 11600 1822 11656
rect 1582 11328 1638 11384
rect 1398 9016 1454 9072
rect 1490 7520 1546 7576
rect 1950 13232 2006 13288
rect 2410 15544 2466 15600
rect 2226 14048 2282 14104
rect 2318 12688 2374 12744
rect 2318 12416 2374 12472
rect 2226 12164 2282 12200
rect 2226 12144 2228 12164
rect 2228 12144 2280 12164
rect 2280 12144 2282 12164
rect 2226 11872 2282 11928
rect 2134 11464 2190 11520
rect 2226 11328 2282 11384
rect 2410 10920 2466 10976
rect 1674 4256 1730 4312
rect 662 3168 718 3224
rect 846 3168 902 3224
rect 294 1672 350 1728
rect 1398 2644 1454 2680
rect 1398 2624 1400 2644
rect 1400 2624 1452 2644
rect 1452 2624 1454 2644
rect 1582 3712 1638 3768
rect 1858 4120 1914 4176
rect 2134 6568 2190 6624
rect 2410 7812 2466 7848
rect 2410 7792 2412 7812
rect 2412 7792 2464 7812
rect 2464 7792 2466 7812
rect 24214 27648 24270 27704
rect 4066 27104 4122 27160
rect 3698 26036 3754 26072
rect 3698 26016 3700 26036
rect 3700 26016 3752 26036
rect 3752 26016 3754 26036
rect 4066 25336 4122 25392
rect 3514 24656 3570 24712
rect 2778 23704 2834 23760
rect 2778 23024 2834 23080
rect 2870 18944 2926 19000
rect 2778 17448 2834 17504
rect 2778 17060 2834 17096
rect 2778 17040 2780 17060
rect 2780 17040 2832 17060
rect 2832 17040 2834 17060
rect 2686 16632 2742 16688
rect 3146 16632 3202 16688
rect 2870 16516 2926 16552
rect 2870 16496 2872 16516
rect 2872 16496 2924 16516
rect 2924 16496 2926 16516
rect 2870 15680 2926 15736
rect 3054 13776 3110 13832
rect 2962 12960 3018 13016
rect 3238 14864 3294 14920
rect 3238 13912 3294 13968
rect 3146 12688 3202 12744
rect 3054 12008 3110 12064
rect 2870 9324 2872 9344
rect 2872 9324 2924 9344
rect 2924 9324 2926 9344
rect 2870 9288 2926 9324
rect 3146 10104 3202 10160
rect 3146 9424 3202 9480
rect 2226 5208 2282 5264
rect 2134 4936 2190 4992
rect 2318 4528 2374 4584
rect 3974 21936 4030 21992
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 7838 24792 7894 24848
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4710 22344 4766 22400
rect 4342 19080 4398 19136
rect 4250 17992 4306 18048
rect 3974 16496 4030 16552
rect 4066 16224 4122 16280
rect 4158 15988 4160 16008
rect 4160 15988 4212 16008
rect 4212 15988 4214 16008
rect 4158 15952 4214 15988
rect 4342 15816 4398 15872
rect 3974 14592 4030 14648
rect 3974 13912 4030 13968
rect 3882 13776 3938 13832
rect 3882 13640 3938 13696
rect 3698 13232 3754 13288
rect 3606 12688 3662 12744
rect 3514 11872 3570 11928
rect 3330 9832 3386 9888
rect 3330 9560 3386 9616
rect 3790 11736 3846 11792
rect 3974 12588 3976 12608
rect 3976 12588 4028 12608
rect 4028 12588 4030 12608
rect 3974 12552 4030 12588
rect 4158 12280 4214 12336
rect 4342 12688 4398 12744
rect 3882 11348 3938 11384
rect 3882 11328 3884 11348
rect 3884 11328 3936 11348
rect 3936 11328 3938 11348
rect 3882 11212 3938 11248
rect 3882 11192 3884 11212
rect 3884 11192 3936 11212
rect 3936 11192 3938 11212
rect 3790 10648 3846 10704
rect 4066 10376 4122 10432
rect 3790 10240 3846 10296
rect 3790 9560 3846 9616
rect 3606 9424 3662 9480
rect 3790 9424 3846 9480
rect 2962 3984 3018 4040
rect 2870 3576 2926 3632
rect 2594 3032 2650 3088
rect 2502 2796 2504 2816
rect 2504 2796 2556 2816
rect 2556 2796 2558 2816
rect 2502 2760 2558 2796
rect 2410 1944 2466 2000
rect 3238 6024 3294 6080
rect 3606 9152 3662 9208
rect 3790 8200 3846 8256
rect 3514 7948 3570 7984
rect 3514 7928 3516 7948
rect 3516 7928 3568 7948
rect 3568 7928 3570 7948
rect 3974 7540 4030 7576
rect 3974 7520 3976 7540
rect 3976 7520 4028 7540
rect 4028 7520 4030 7540
rect 3422 6024 3478 6080
rect 3330 5888 3386 5944
rect 3606 5752 3662 5808
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4618 16768 4674 16824
rect 4526 15272 4582 15328
rect 4526 11736 4582 11792
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5354 20168 5410 20224
rect 5262 17040 5318 17096
rect 4710 11872 4766 11928
rect 4618 9832 4674 9888
rect 4526 9036 4582 9072
rect 4526 9016 4528 9036
rect 4528 9016 4580 9036
rect 4580 9016 4582 9036
rect 4894 14048 4950 14104
rect 4802 10920 4858 10976
rect 3146 3576 3202 3632
rect 3422 3440 3478 3496
rect 3422 2524 3424 2544
rect 3424 2524 3476 2544
rect 3476 2524 3478 2544
rect 3422 2488 3478 2524
rect 2870 856 2926 912
rect 3974 4800 4030 4856
rect 4250 4120 4306 4176
rect 3882 3440 3938 3496
rect 4158 2896 4214 2952
rect 3790 1400 3846 1456
rect 4434 2624 4490 2680
rect 3698 312 3754 368
rect 4894 8472 4950 8528
rect 4802 8200 4858 8256
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5538 15428 5594 15464
rect 5538 15408 5540 15428
rect 5540 15408 5592 15428
rect 5592 15408 5594 15428
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 7102 16496 7158 16552
rect 7010 15544 7066 15600
rect 5446 14320 5502 14376
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6182 13368 6238 13424
rect 6734 14184 6790 14240
rect 6458 12552 6514 12608
rect 6642 12960 6698 13016
rect 6550 12416 6606 12472
rect 6090 12300 6146 12336
rect 6090 12280 6092 12300
rect 6092 12280 6144 12300
rect 6144 12280 6146 12300
rect 5998 11600 6054 11656
rect 6182 10920 6238 10976
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6366 10512 6422 10568
rect 6182 10376 6238 10432
rect 6642 10684 6644 10704
rect 6644 10684 6696 10704
rect 6696 10684 6698 10704
rect 6642 10648 6698 10684
rect 6458 10412 6460 10432
rect 6460 10412 6512 10432
rect 6512 10412 6514 10432
rect 6458 10376 6514 10412
rect 6458 10240 6514 10296
rect 6366 9832 6422 9888
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 4986 6568 5042 6624
rect 5078 6196 5080 6216
rect 5080 6196 5132 6216
rect 5132 6196 5134 6216
rect 5078 6160 5134 6196
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6366 8336 6422 8392
rect 5630 8064 5686 8120
rect 5998 7656 6054 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6090 7112 6146 7168
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5630 6316 5686 6352
rect 5630 6296 5632 6316
rect 5632 6296 5684 6316
rect 5684 6296 5686 6316
rect 5446 5616 5502 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4986 4276 5042 4312
rect 4986 4256 4988 4276
rect 4988 4256 5040 4276
rect 5040 4256 5042 4276
rect 4802 3984 4858 4040
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4894 2624 4950 2680
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6274 6704 6330 6760
rect 6274 5072 6330 5128
rect 6918 12860 6920 12880
rect 6920 12860 6972 12880
rect 6972 12860 6974 12880
rect 6918 12824 6974 12860
rect 6826 12688 6882 12744
rect 6918 12180 6920 12200
rect 6920 12180 6972 12200
rect 6972 12180 6974 12200
rect 6918 12144 6974 12180
rect 7378 11636 7380 11656
rect 7380 11636 7432 11656
rect 7432 11636 7434 11656
rect 7378 11600 7434 11636
rect 7102 11192 7158 11248
rect 7378 10004 7380 10024
rect 7380 10004 7432 10024
rect 7432 10004 7434 10024
rect 7378 9968 7434 10004
rect 7286 9560 7342 9616
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9310 23024 9366 23080
rect 8758 20304 8814 20360
rect 8482 15952 8538 16008
rect 8022 13640 8078 13696
rect 8206 13812 8208 13832
rect 8208 13812 8260 13832
rect 8260 13812 8262 13832
rect 8206 13776 8262 13812
rect 8206 11756 8262 11792
rect 8206 11736 8208 11756
rect 8208 11736 8260 11756
rect 8260 11736 8262 11756
rect 8114 11192 8170 11248
rect 8574 14320 8630 14376
rect 7470 8608 7526 8664
rect 6826 5888 6882 5944
rect 6550 4020 6552 4040
rect 6552 4020 6604 4040
rect 6604 4020 6606 4040
rect 6550 3984 6606 4020
rect 6182 1944 6238 2000
rect 7102 6740 7104 6760
rect 7104 6740 7156 6760
rect 7156 6740 7158 6760
rect 7102 6704 7158 6740
rect 7102 5888 7158 5944
rect 6918 4800 6974 4856
rect 6826 2796 6828 2816
rect 6828 2796 6880 2816
rect 6880 2796 6882 2816
rect 6826 2760 6882 2796
rect 6458 2644 6514 2680
rect 7378 6024 7434 6080
rect 7746 5344 7802 5400
rect 7654 4664 7710 4720
rect 8758 11600 8814 11656
rect 8942 11192 8998 11248
rect 8390 9560 8446 9616
rect 8298 8472 8354 8528
rect 8758 8880 8814 8936
rect 8482 8200 8538 8256
rect 8206 6160 8262 6216
rect 8298 5208 8354 5264
rect 8114 4564 8116 4584
rect 8116 4564 8168 4584
rect 8168 4564 8170 4584
rect 8114 4528 8170 4564
rect 8022 4020 8024 4040
rect 8024 4020 8076 4040
rect 8076 4020 8078 4040
rect 8022 3984 8078 4020
rect 8298 3848 8354 3904
rect 8574 6452 8630 6488
rect 8574 6432 8576 6452
rect 8576 6432 8628 6452
rect 8628 6432 8630 6452
rect 8666 6160 8722 6216
rect 8298 3596 8354 3632
rect 8298 3576 8300 3596
rect 8300 3576 8352 3596
rect 8352 3576 8354 3596
rect 6458 2624 6460 2644
rect 6460 2624 6512 2644
rect 6512 2624 6514 2644
rect 8022 3068 8024 3088
rect 8024 3068 8076 3088
rect 8076 3068 8078 3088
rect 8022 3032 8078 3068
rect 8206 2508 8262 2544
rect 8206 2488 8208 2508
rect 8208 2488 8260 2508
rect 8260 2488 8262 2508
rect 8022 1536 8078 1592
rect 8574 2760 8630 2816
rect 8850 1808 8906 1864
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 12346 24656 12402 24712
rect 10782 20440 10838 20496
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11886 17720 11942 17776
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10138 16088 10194 16144
rect 9494 15408 9550 15464
rect 9770 13640 9826 13696
rect 9586 12960 9642 13016
rect 9954 13232 10010 13288
rect 9770 13096 9826 13152
rect 9586 11328 9642 11384
rect 9310 9288 9366 9344
rect 9218 3168 9274 3224
rect 9678 10956 9680 10976
rect 9680 10956 9732 10976
rect 9732 10956 9734 10976
rect 9678 10920 9734 10956
rect 9678 10648 9734 10704
rect 9678 9036 9734 9072
rect 9678 9016 9680 9036
rect 9680 9016 9732 9036
rect 9732 9016 9734 9036
rect 9862 10920 9918 10976
rect 9402 6296 9458 6352
rect 9402 5888 9458 5944
rect 9586 6704 9642 6760
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10690 13776 10746 13832
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11702 12824 11758 12880
rect 11702 12436 11758 12472
rect 11702 12416 11704 12436
rect 11704 12416 11756 12436
rect 11756 12416 11758 12436
rect 11610 12280 11666 12336
rect 10874 11464 10930 11520
rect 10782 11328 10838 11384
rect 10322 11056 10378 11112
rect 10046 10412 10048 10432
rect 10048 10412 10100 10432
rect 10100 10412 10102 10432
rect 10046 10376 10102 10412
rect 10046 10240 10102 10296
rect 9862 8608 9918 8664
rect 9770 8336 9826 8392
rect 9862 8064 9918 8120
rect 10230 10668 10286 10704
rect 10230 10648 10232 10668
rect 10232 10648 10284 10668
rect 10284 10648 10286 10668
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9696 10194 9752
rect 11150 10376 11206 10432
rect 11426 10376 11482 10432
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11150 10240 11206 10296
rect 10966 8472 11022 8528
rect 10138 8200 10194 8256
rect 10690 8200 10746 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10138 7656 10194 7712
rect 10322 7656 10378 7712
rect 10046 7520 10102 7576
rect 10690 7248 10746 7304
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9954 5636 10010 5672
rect 9954 5616 9956 5636
rect 9956 5616 10008 5636
rect 10008 5616 10010 5636
rect 9954 5208 10010 5264
rect 9126 2624 9182 2680
rect 9034 1672 9090 1728
rect 9954 4936 10010 4992
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11242 8336 11298 8392
rect 11058 6296 11114 6352
rect 10690 5208 10746 5264
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9862 3712 9918 3768
rect 10690 3848 10746 3904
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10782 3712 10838 3768
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10322 2352 10378 2408
rect 10874 2372 10930 2408
rect 10874 2352 10876 2372
rect 10876 2352 10928 2372
rect 10928 2352 10930 2372
rect 10782 2216 10838 2272
rect 10874 1536 10930 1592
rect 11334 6296 11390 6352
rect 11426 5888 11482 5944
rect 11702 10104 11758 10160
rect 12162 9968 12218 10024
rect 12162 9696 12218 9752
rect 12162 9444 12218 9480
rect 12162 9424 12164 9444
rect 12164 9424 12216 9444
rect 12216 9424 12218 9444
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 17038 20440 17094 20496
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16946 19216 17002 19272
rect 15566 18808 15622 18864
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 12622 18264 12678 18320
rect 12438 15680 12494 15736
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 12530 13388 12586 13424
rect 12530 13368 12532 13388
rect 12532 13368 12584 13388
rect 12584 13368 12586 13388
rect 12438 11772 12440 11792
rect 12440 11772 12492 11792
rect 12492 11772 12494 11792
rect 12438 11736 12494 11772
rect 12530 11600 12586 11656
rect 12622 11056 12678 11112
rect 11610 4936 11666 4992
rect 11978 6976 12034 7032
rect 12622 9424 12678 9480
rect 12162 7792 12218 7848
rect 12162 7420 12164 7440
rect 12164 7420 12216 7440
rect 12216 7420 12218 7440
rect 12162 7384 12218 7420
rect 12438 7284 12440 7304
rect 12440 7284 12492 7304
rect 12492 7284 12494 7304
rect 12438 7248 12494 7284
rect 11242 2644 11298 2680
rect 11242 2624 11244 2644
rect 11244 2624 11296 2644
rect 11296 2624 11298 2644
rect 11058 1400 11114 1456
rect 12162 6724 12218 6760
rect 12162 6704 12164 6724
rect 12164 6704 12216 6724
rect 12216 6704 12218 6724
rect 12162 5752 12218 5808
rect 12438 4936 12494 4992
rect 11978 4528 12034 4584
rect 11794 4256 11850 4312
rect 11518 4120 11574 4176
rect 11610 1400 11666 1456
rect 12162 3984 12218 4040
rect 12806 10104 12862 10160
rect 12806 8200 12862 8256
rect 12806 7656 12862 7712
rect 13174 16632 13230 16688
rect 13542 15816 13598 15872
rect 13174 11736 13230 11792
rect 13450 15544 13506 15600
rect 13726 13504 13782 13560
rect 13450 11192 13506 11248
rect 13174 10648 13230 10704
rect 13082 9288 13138 9344
rect 13082 7792 13138 7848
rect 12806 4392 12862 4448
rect 13082 3984 13138 4040
rect 12622 3440 12678 3496
rect 13266 5208 13322 5264
rect 13450 6160 13506 6216
rect 13450 4392 13506 4448
rect 13450 4256 13506 4312
rect 13358 3848 13414 3904
rect 13634 10648 13690 10704
rect 13818 9696 13874 9752
rect 13726 9152 13782 9208
rect 13634 7964 13636 7984
rect 13636 7964 13688 7984
rect 13688 7964 13690 7984
rect 13634 7928 13690 7964
rect 13634 7112 13690 7168
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14186 9868 14188 9888
rect 14188 9868 14240 9888
rect 14240 9868 14242 9888
rect 14186 9832 14242 9868
rect 14002 6840 14058 6896
rect 13910 5616 13966 5672
rect 14646 14728 14702 14784
rect 14738 14184 14794 14240
rect 14370 10512 14426 10568
rect 14462 9968 14518 10024
rect 14462 9596 14464 9616
rect 14464 9596 14516 9616
rect 14516 9596 14518 9616
rect 14462 9560 14518 9596
rect 14646 10784 14702 10840
rect 14646 10240 14702 10296
rect 14554 9288 14610 9344
rect 14462 7520 14518 7576
rect 14094 4120 14150 4176
rect 14554 6024 14610 6080
rect 14462 3576 14518 3632
rect 13634 2896 13690 2952
rect 14186 3032 14242 3088
rect 13726 2760 13782 2816
rect 15382 15680 15438 15736
rect 15014 15444 15016 15464
rect 15016 15444 15068 15464
rect 15068 15444 15070 15464
rect 15014 15408 15070 15444
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15014 14592 15070 14648
rect 15014 14340 15070 14376
rect 15014 14320 15016 14340
rect 15016 14320 15068 14340
rect 15068 14320 15070 14340
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15106 13912 15162 13968
rect 15290 13912 15346 13968
rect 15474 14864 15530 14920
rect 15658 14764 15660 14784
rect 15660 14764 15712 14784
rect 15712 14764 15714 14784
rect 15658 14728 15714 14764
rect 15750 14320 15806 14376
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15106 12552 15162 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14922 11636 14924 11656
rect 14924 11636 14976 11656
rect 14976 11636 14978 11656
rect 14922 11600 14978 11636
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15474 12824 15530 12880
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 9868 15384 9888
rect 15384 9868 15436 9888
rect 15436 9868 15438 9888
rect 15382 9832 15438 9868
rect 14830 9324 14832 9344
rect 14832 9324 14884 9344
rect 14884 9324 14886 9344
rect 14830 9288 14886 9324
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15290 8336 15346 8392
rect 14738 7656 14794 7712
rect 14646 5652 14648 5672
rect 14648 5652 14700 5672
rect 14700 5652 14702 5672
rect 14646 5616 14702 5652
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15934 13504 15990 13560
rect 16210 14048 16266 14104
rect 16026 13268 16028 13288
rect 16028 13268 16080 13288
rect 16080 13268 16082 13288
rect 16026 13232 16082 13268
rect 16210 13132 16212 13152
rect 16212 13132 16264 13152
rect 16264 13132 16266 13152
rect 16210 13096 16266 13132
rect 15934 12008 15990 12064
rect 15658 9172 15714 9208
rect 16026 11328 16082 11384
rect 15842 9696 15898 9752
rect 15658 9152 15660 9172
rect 15660 9152 15712 9172
rect 15712 9152 15714 9172
rect 15474 7248 15530 7304
rect 15566 7148 15568 7168
rect 15568 7148 15620 7168
rect 15620 7148 15622 7168
rect 15566 7112 15622 7148
rect 14646 3712 14702 3768
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 2896 14610 2952
rect 14830 2896 14886 2952
rect 15106 2916 15162 2952
rect 15106 2896 15108 2916
rect 15108 2896 15160 2916
rect 15160 2896 15162 2916
rect 14646 2624 14702 2680
rect 14462 2216 14518 2272
rect 14002 1808 14058 1864
rect 14278 1264 14334 1320
rect 15842 7384 15898 7440
rect 15842 5364 15898 5400
rect 15842 5344 15844 5364
rect 15844 5344 15896 5364
rect 15896 5344 15898 5364
rect 15750 3984 15806 4040
rect 15842 3884 15844 3904
rect 15844 3884 15896 3904
rect 15896 3884 15898 3904
rect 15842 3848 15898 3884
rect 15842 3732 15898 3768
rect 15842 3712 15844 3732
rect 15844 3712 15896 3732
rect 15896 3712 15898 3732
rect 16394 12688 16450 12744
rect 16394 12144 16450 12200
rect 16762 12588 16764 12608
rect 16764 12588 16816 12608
rect 16816 12588 16818 12608
rect 16762 12552 16818 12588
rect 16578 12180 16580 12200
rect 16580 12180 16632 12200
rect 16632 12180 16634 12200
rect 16578 12144 16634 12180
rect 16394 11600 16450 11656
rect 16670 8472 16726 8528
rect 24030 27104 24086 27160
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 23662 24384 23718 24440
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 21730 22616 21786 22672
rect 20810 22344 20866 22400
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18234 20440 18290 20496
rect 17498 20304 17554 20360
rect 19062 18672 19118 18728
rect 17958 15580 17960 15600
rect 17960 15580 18012 15600
rect 18012 15580 18014 15600
rect 17958 15544 18014 15580
rect 17038 14184 17094 14240
rect 16302 7656 16358 7712
rect 16118 6432 16174 6488
rect 16486 5752 16542 5808
rect 16302 3712 16358 3768
rect 15934 3168 15990 3224
rect 15842 3032 15898 3088
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15474 2372 15530 2408
rect 15474 2352 15476 2372
rect 15476 2352 15528 2372
rect 15528 2352 15530 2372
rect 15934 2644 15990 2680
rect 15934 2624 15936 2644
rect 15936 2624 15988 2644
rect 15988 2624 15990 2644
rect 16486 3984 16542 4040
rect 16762 4020 16764 4040
rect 16764 4020 16816 4040
rect 16816 4020 16818 4040
rect 16762 3984 16818 4020
rect 16486 3712 16542 3768
rect 16578 3032 16634 3088
rect 17222 13812 17224 13832
rect 17224 13812 17276 13832
rect 17276 13812 17278 13832
rect 17222 13776 17278 13812
rect 17222 13368 17278 13424
rect 17130 12144 17186 12200
rect 17130 11736 17186 11792
rect 17130 11464 17186 11520
rect 16946 5344 17002 5400
rect 16946 5208 17002 5264
rect 17038 4528 17094 4584
rect 18050 14184 18106 14240
rect 18050 13912 18106 13968
rect 17406 10104 17462 10160
rect 17406 8200 17462 8256
rect 17222 7520 17278 7576
rect 17222 5616 17278 5672
rect 17958 12144 18014 12200
rect 17774 11892 17830 11928
rect 17774 11872 17776 11892
rect 17776 11872 17828 11892
rect 17828 11872 17830 11892
rect 17774 10140 17776 10160
rect 17776 10140 17828 10160
rect 17828 10140 17830 10160
rect 17774 10104 17830 10140
rect 17774 9152 17830 9208
rect 18326 14184 18382 14240
rect 18510 13232 18566 13288
rect 17590 5616 17646 5672
rect 17498 4684 17554 4720
rect 17498 4664 17500 4684
rect 17500 4664 17552 4684
rect 17552 4664 17554 4684
rect 17222 4392 17278 4448
rect 17130 3984 17186 4040
rect 17222 3576 17278 3632
rect 16394 2488 16450 2544
rect 17222 3304 17278 3360
rect 17038 2896 17094 2952
rect 17498 2796 17500 2816
rect 17500 2796 17552 2816
rect 17552 2796 17554 2816
rect 17498 2760 17554 2796
rect 16762 1808 16818 1864
rect 16854 1672 16910 1728
rect 17038 1400 17094 1456
rect 18050 6024 18106 6080
rect 17866 5616 17922 5672
rect 17774 5092 17830 5128
rect 17774 5072 17776 5092
rect 17776 5072 17828 5092
rect 17828 5072 17830 5092
rect 18970 15000 19026 15056
rect 18786 14456 18842 14512
rect 19062 14592 19118 14648
rect 18326 9560 18382 9616
rect 18510 9560 18566 9616
rect 18510 9288 18566 9344
rect 18234 8064 18290 8120
rect 18970 12824 19026 12880
rect 18970 10920 19026 10976
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19982 17584 20038 17640
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20718 16632 20774 16688
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19430 14764 19432 14784
rect 19432 14764 19484 14784
rect 19484 14764 19486 14784
rect 19430 14728 19486 14764
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13776 19486 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20166 13776 20222 13832
rect 20258 12960 20314 13016
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20166 12552 20222 12608
rect 19338 11872 19394 11928
rect 19982 12144 20038 12200
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19706 10920 19762 10976
rect 19522 10648 19578 10704
rect 19430 10512 19486 10568
rect 19614 10512 19670 10568
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18694 7692 18696 7712
rect 18696 7692 18748 7712
rect 18748 7692 18750 7712
rect 18694 7656 18750 7692
rect 18786 7520 18842 7576
rect 18234 5480 18290 5536
rect 18234 5208 18290 5264
rect 18050 2624 18106 2680
rect 18050 2508 18106 2544
rect 18050 2488 18052 2508
rect 18052 2488 18104 2508
rect 18104 2488 18106 2508
rect 18694 5888 18750 5944
rect 18326 2488 18382 2544
rect 17682 2100 17738 2136
rect 17682 2080 17684 2100
rect 17684 2080 17736 2100
rect 17736 2080 17738 2100
rect 18142 1944 18198 2000
rect 19982 9560 20038 9616
rect 20442 15136 20498 15192
rect 20626 15136 20682 15192
rect 20534 14320 20590 14376
rect 20442 13640 20498 13696
rect 20442 12416 20498 12472
rect 20350 10784 20406 10840
rect 20442 9832 20498 9888
rect 19338 8200 19394 8256
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19890 8628 19946 8664
rect 19890 8608 19892 8628
rect 19892 8608 19944 8628
rect 19944 8608 19946 8628
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19430 7828 19432 7848
rect 19432 7828 19484 7848
rect 19484 7828 19486 7848
rect 19430 7792 19486 7828
rect 20074 7520 20130 7576
rect 19246 6840 19302 6896
rect 19522 7384 19578 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20074 6976 20130 7032
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 18878 3612 18880 3632
rect 18880 3612 18932 3632
rect 18932 3612 18934 3632
rect 18878 3576 18934 3612
rect 19154 4156 19156 4176
rect 19156 4156 19208 4176
rect 19208 4156 19210 4176
rect 19154 4120 19210 4156
rect 19062 3032 19118 3088
rect 19338 5752 19394 5808
rect 19522 5752 19578 5808
rect 20166 5888 20222 5944
rect 19430 5344 19486 5400
rect 19706 5072 19762 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20350 9016 20406 9072
rect 20350 7812 20406 7848
rect 20350 7792 20352 7812
rect 20352 7792 20404 7812
rect 20404 7792 20406 7812
rect 23202 22480 23258 22536
rect 23478 22380 23480 22400
rect 23480 22380 23532 22400
rect 23532 22380 23534 22400
rect 23478 22344 23534 22380
rect 21270 17720 21326 17776
rect 20994 16768 21050 16824
rect 21178 14864 21234 14920
rect 20902 12824 20958 12880
rect 21086 12008 21142 12064
rect 21730 15972 21786 16008
rect 21730 15952 21732 15972
rect 21732 15952 21784 15972
rect 21784 15952 21786 15972
rect 21546 14884 21602 14920
rect 21546 14864 21548 14884
rect 21548 14864 21600 14884
rect 21600 14864 21602 14884
rect 21454 14456 21510 14512
rect 22098 15816 22154 15872
rect 22006 15408 22062 15464
rect 22466 16904 22522 16960
rect 22650 16632 22706 16688
rect 21822 11076 21878 11112
rect 21822 11056 21824 11076
rect 21824 11056 21876 11076
rect 21876 11056 21878 11076
rect 21730 10104 21786 10160
rect 21270 8880 21326 8936
rect 20902 7792 20958 7848
rect 20902 6840 20958 6896
rect 19430 3884 19432 3904
rect 19432 3884 19484 3904
rect 19484 3884 19486 3904
rect 19430 3848 19486 3884
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19430 3712 19486 3768
rect 19522 3440 19578 3496
rect 19706 3440 19762 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20258 3576 20314 3632
rect 20258 3304 20314 3360
rect 21546 8608 21602 8664
rect 21362 6704 21418 6760
rect 21270 5616 21326 5672
rect 20810 3984 20866 4040
rect 20166 1400 20222 1456
rect 20718 3032 20774 3088
rect 20534 2508 20590 2544
rect 20534 2488 20536 2508
rect 20536 2488 20588 2508
rect 20588 2488 20590 2508
rect 21546 6160 21602 6216
rect 22190 9968 22246 10024
rect 21914 9424 21970 9480
rect 21730 6840 21786 6896
rect 21638 6024 21694 6080
rect 21546 5616 21602 5672
rect 21546 2488 21602 2544
rect 21822 6568 21878 6624
rect 22190 9288 22246 9344
rect 22098 8628 22154 8664
rect 22098 8608 22100 8628
rect 22100 8608 22152 8628
rect 22152 8608 22154 8628
rect 21822 6432 21878 6488
rect 22006 6432 22062 6488
rect 21822 6160 21878 6216
rect 22190 6316 22246 6352
rect 22190 6296 22192 6316
rect 22192 6296 22244 6316
rect 22244 6296 22246 6316
rect 21914 4936 21970 4992
rect 21914 4800 21970 4856
rect 22006 4120 22062 4176
rect 22098 3168 22154 3224
rect 21454 2216 21510 2272
rect 22742 14728 22798 14784
rect 22558 6296 22614 6352
rect 22558 5752 22614 5808
rect 22558 5344 22614 5400
rect 22558 4936 22614 4992
rect 22374 3712 22430 3768
rect 23018 14456 23074 14512
rect 22926 13096 22982 13152
rect 22834 11056 22890 11112
rect 23018 12552 23074 12608
rect 22926 10512 22982 10568
rect 22834 9696 22890 9752
rect 22742 4972 22744 4992
rect 22744 4972 22796 4992
rect 22796 4972 22798 4992
rect 22742 4936 22798 4972
rect 23938 22072 23994 22128
rect 25410 26560 25466 26616
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24928 24822 24984
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23840 24822 23896
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25134 23160 25190 23216
rect 24950 22516 24952 22536
rect 24952 22516 25004 22536
rect 25004 22516 25006 22536
rect 24950 22480 25006 22516
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21528 24822 21584
rect 24674 20984 24730 21040
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24122 19896 24178 19952
rect 23662 17040 23718 17096
rect 23662 16768 23718 16824
rect 23478 16496 23534 16552
rect 23754 15952 23810 16008
rect 23478 14592 23534 14648
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24582 19252 24584 19272
rect 24584 19252 24636 19272
rect 24636 19252 24638 19272
rect 24582 19216 24638 19252
rect 24766 19352 24822 19408
rect 24398 18672 24454 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24582 18264 24638 18320
rect 24766 18128 24822 18184
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24490 16632 24546 16688
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24030 15952 24086 16008
rect 23846 15136 23902 15192
rect 23754 14864 23810 14920
rect 23662 13776 23718 13832
rect 23846 13504 23902 13560
rect 23294 12280 23350 12336
rect 23662 12416 23718 12472
rect 23662 12280 23718 12336
rect 23478 9152 23534 9208
rect 23662 8472 23718 8528
rect 23846 9424 23902 9480
rect 23754 6704 23810 6760
rect 23754 6296 23810 6352
rect 23662 6024 23718 6080
rect 22834 3984 22890 4040
rect 22742 3848 22798 3904
rect 23018 3440 23074 3496
rect 23478 5480 23534 5536
rect 23478 5344 23534 5400
rect 23478 4392 23534 4448
rect 23754 4664 23810 4720
rect 23570 3576 23626 3632
rect 23202 2624 23258 2680
rect 22558 2080 22614 2136
rect 23018 1672 23074 1728
rect 23478 2372 23534 2408
rect 23478 2352 23480 2372
rect 23480 2352 23532 2372
rect 23532 2352 23534 2372
rect 23478 2216 23534 2272
rect 24674 15580 24676 15600
rect 24676 15580 24728 15600
rect 24728 15580 24730 15600
rect 24674 15544 24730 15580
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24950 16904 25006 16960
rect 25042 15852 25044 15872
rect 25044 15852 25096 15872
rect 25096 15852 25098 15872
rect 25042 15816 25098 15852
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25042 13912 25098 13968
rect 24766 13640 24822 13696
rect 24674 13096 24730 13152
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11192 24822 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24766 10104 24822 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 9016 24822 9072
rect 25226 14728 25282 14784
rect 25502 26016 25558 26072
rect 25870 25472 25926 25528
rect 25778 15000 25834 15056
rect 25318 13232 25374 13288
rect 25318 11772 25320 11792
rect 25320 11772 25372 11792
rect 25372 11772 25374 11792
rect 25318 11736 25374 11772
rect 25502 11056 25558 11112
rect 25318 10512 25374 10568
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24030 6568 24086 6624
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24122 6432 24178 6488
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 23938 5208 23994 5264
rect 24582 5072 24638 5128
rect 23938 4936 23994 4992
rect 23846 1944 23902 2000
rect 25594 9968 25650 10024
rect 25134 6840 25190 6896
rect 25042 6704 25098 6760
rect 24674 4664 24730 4720
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24122 4276 24178 4312
rect 24122 4256 24124 4276
rect 24124 4256 24176 4276
rect 24176 4256 24178 4276
rect 24674 4256 24730 4312
rect 24950 4120 25006 4176
rect 24122 3984 24178 4040
rect 24582 3712 24638 3768
rect 24306 3576 24362 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24030 2896 24086 2952
rect 24030 2488 24086 2544
rect 24766 2488 24822 2544
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23754 1536 23810 1592
rect 23938 1536 23994 1592
rect 23478 856 23534 912
rect 4618 40 4674 96
rect 25134 3848 25190 3904
rect 25410 6160 25466 6216
rect 25318 6024 25374 6080
rect 25962 7792 26018 7848
rect 25962 6060 25964 6080
rect 25964 6060 26016 6080
rect 26016 6060 26018 6080
rect 25962 6024 26018 6060
rect 25962 5616 26018 5672
rect 25870 3032 25926 3088
rect 25594 2644 25650 2680
rect 25594 2624 25596 2644
rect 25596 2624 25648 2644
rect 25648 2624 25650 2644
rect 24214 40 24270 96
rect 27618 1672 27674 1728
rect 26790 1400 26846 1456
rect 26146 312 26202 368
<< metal3 >>
rect 0 27706 480 27736
rect 3417 27706 3483 27709
rect 0 27704 3483 27706
rect 0 27648 3422 27704
rect 3478 27648 3483 27704
rect 0 27646 3483 27648
rect 0 27616 480 27646
rect 3417 27643 3483 27646
rect 24209 27706 24275 27709
rect 27520 27706 28000 27736
rect 24209 27704 28000 27706
rect 24209 27648 24214 27704
rect 24270 27648 28000 27704
rect 24209 27646 28000 27648
rect 24209 27643 24275 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 4061 27162 4127 27165
rect 0 27160 4127 27162
rect 0 27104 4066 27160
rect 4122 27104 4127 27160
rect 0 27102 4127 27104
rect 0 27072 480 27102
rect 4061 27099 4127 27102
rect 24025 27162 24091 27165
rect 27520 27162 28000 27192
rect 24025 27160 28000 27162
rect 24025 27104 24030 27160
rect 24086 27104 28000 27160
rect 24025 27102 28000 27104
rect 24025 27099 24091 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 2681 26618 2747 26621
rect 0 26616 2747 26618
rect 0 26560 2686 26616
rect 2742 26560 2747 26616
rect 0 26558 2747 26560
rect 0 26528 480 26558
rect 2681 26555 2747 26558
rect 25405 26618 25471 26621
rect 27520 26618 28000 26648
rect 25405 26616 28000 26618
rect 25405 26560 25410 26616
rect 25466 26560 28000 26616
rect 25405 26558 28000 26560
rect 25405 26555 25471 26558
rect 27520 26528 28000 26558
rect 0 26074 480 26104
rect 3693 26074 3759 26077
rect 0 26072 3759 26074
rect 0 26016 3698 26072
rect 3754 26016 3759 26072
rect 0 26014 3759 26016
rect 0 25984 480 26014
rect 3693 26011 3759 26014
rect 25497 26074 25563 26077
rect 27520 26074 28000 26104
rect 25497 26072 28000 26074
rect 25497 26016 25502 26072
rect 25558 26016 28000 26072
rect 25497 26014 28000 26016
rect 25497 26011 25563 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 25865 25530 25931 25533
rect 27520 25530 28000 25560
rect 25865 25528 28000 25530
rect 25865 25472 25870 25528
rect 25926 25472 28000 25528
rect 25865 25470 28000 25472
rect 25865 25467 25931 25470
rect 27520 25440 28000 25470
rect 0 25394 480 25424
rect 4061 25394 4127 25397
rect 0 25392 4127 25394
rect 0 25336 4066 25392
rect 4122 25336 4127 25392
rect 0 25334 4127 25336
rect 0 25304 480 25334
rect 4061 25331 4127 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 24761 24986 24827 24989
rect 27520 24986 28000 25016
rect 24761 24984 28000 24986
rect 24761 24928 24766 24984
rect 24822 24928 28000 24984
rect 24761 24926 28000 24928
rect 24761 24923 24827 24926
rect 27520 24896 28000 24926
rect 0 24850 480 24880
rect 7833 24850 7899 24853
rect 0 24848 7899 24850
rect 0 24792 7838 24848
rect 7894 24792 7899 24848
rect 0 24790 7899 24792
rect 0 24760 480 24790
rect 7833 24787 7899 24790
rect 3509 24714 3575 24717
rect 12341 24714 12407 24717
rect 3509 24712 12407 24714
rect 3509 24656 3514 24712
rect 3570 24656 12346 24712
rect 12402 24656 12407 24712
rect 3509 24654 12407 24656
rect 3509 24651 3575 24654
rect 12341 24651 12407 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 23657 24442 23723 24445
rect 27520 24442 28000 24472
rect 23657 24440 28000 24442
rect 23657 24384 23662 24440
rect 23718 24384 28000 24440
rect 23657 24382 28000 24384
rect 23657 24379 23723 24382
rect 27520 24352 28000 24382
rect 0 24306 480 24336
rect 1577 24306 1643 24309
rect 0 24304 1643 24306
rect 0 24248 1582 24304
rect 1638 24248 1643 24304
rect 0 24246 1643 24248
rect 0 24216 480 24246
rect 1577 24243 1643 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24761 23898 24827 23901
rect 27520 23898 28000 23928
rect 24761 23896 28000 23898
rect 24761 23840 24766 23896
rect 24822 23840 28000 23896
rect 24761 23838 28000 23840
rect 24761 23835 24827 23838
rect 27520 23808 28000 23838
rect 0 23762 480 23792
rect 2773 23762 2839 23765
rect 0 23760 2839 23762
rect 0 23704 2778 23760
rect 2834 23704 2839 23760
rect 0 23702 2839 23704
rect 0 23672 480 23702
rect 2773 23699 2839 23702
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 480 23158
rect 1485 23155 1551 23158
rect 25129 23218 25195 23221
rect 27520 23218 28000 23248
rect 25129 23216 28000 23218
rect 25129 23160 25134 23216
rect 25190 23160 28000 23216
rect 25129 23158 28000 23160
rect 25129 23155 25195 23158
rect 27520 23128 28000 23158
rect 2773 23082 2839 23085
rect 9305 23082 9371 23085
rect 2773 23080 9371 23082
rect 2773 23024 2778 23080
rect 2834 23024 9310 23080
rect 9366 23024 9371 23080
rect 2773 23022 9371 23024
rect 2773 23019 2839 23022
rect 9305 23019 9371 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 21725 22674 21791 22677
rect 27520 22674 28000 22704
rect 21725 22672 28000 22674
rect 21725 22616 21730 22672
rect 21786 22616 28000 22672
rect 21725 22614 28000 22616
rect 21725 22611 21791 22614
rect 27520 22584 28000 22614
rect 0 22538 480 22568
rect 2589 22538 2655 22541
rect 0 22536 2655 22538
rect 0 22480 2594 22536
rect 2650 22480 2655 22536
rect 0 22478 2655 22480
rect 0 22448 480 22478
rect 2589 22475 2655 22478
rect 23197 22538 23263 22541
rect 24945 22538 25011 22541
rect 23197 22536 25011 22538
rect 23197 22480 23202 22536
rect 23258 22480 24950 22536
rect 25006 22480 25011 22536
rect 23197 22478 25011 22480
rect 23197 22475 23263 22478
rect 24945 22475 25011 22478
rect 2037 22402 2103 22405
rect 4705 22402 4771 22405
rect 2037 22400 4771 22402
rect 2037 22344 2042 22400
rect 2098 22344 4710 22400
rect 4766 22344 4771 22400
rect 2037 22342 4771 22344
rect 2037 22339 2103 22342
rect 4705 22339 4771 22342
rect 20805 22402 20871 22405
rect 23473 22402 23539 22405
rect 20805 22400 23539 22402
rect 20805 22344 20810 22400
rect 20866 22344 23478 22400
rect 23534 22344 23539 22400
rect 20805 22342 23539 22344
rect 20805 22339 20871 22342
rect 23473 22339 23539 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 23933 22130 23999 22133
rect 27520 22130 28000 22160
rect 23933 22128 28000 22130
rect 23933 22072 23938 22128
rect 23994 22072 28000 22128
rect 23933 22070 28000 22072
rect 23933 22067 23999 22070
rect 27520 22040 28000 22070
rect 0 21994 480 22024
rect 3969 21994 4035 21997
rect 0 21992 4035 21994
rect 0 21936 3974 21992
rect 4030 21936 4035 21992
rect 0 21934 4035 21936
rect 0 21904 480 21934
rect 3969 21931 4035 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24761 21586 24827 21589
rect 27520 21586 28000 21616
rect 24761 21584 28000 21586
rect 24761 21528 24766 21584
rect 24822 21528 28000 21584
rect 24761 21526 28000 21528
rect 24761 21523 24827 21526
rect 27520 21496 28000 21526
rect 0 21450 480 21480
rect 1485 21450 1551 21453
rect 0 21448 1551 21450
rect 0 21392 1490 21448
rect 1546 21392 1551 21448
rect 0 21390 1551 21392
rect 0 21360 480 21390
rect 1485 21387 1551 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 24669 21042 24735 21045
rect 27520 21042 28000 21072
rect 24669 21040 28000 21042
rect 24669 20984 24674 21040
rect 24730 20984 28000 21040
rect 24669 20982 28000 20984
rect 24669 20979 24735 20982
rect 27520 20952 28000 20982
rect 0 20906 480 20936
rect 1577 20906 1643 20909
rect 0 20904 1643 20906
rect 0 20848 1582 20904
rect 1638 20848 1643 20904
rect 0 20846 1643 20848
rect 0 20816 480 20846
rect 1577 20843 1643 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10777 20498 10843 20501
rect 17033 20498 17099 20501
rect 10777 20496 17099 20498
rect 10777 20440 10782 20496
rect 10838 20440 17038 20496
rect 17094 20440 17099 20496
rect 10777 20438 17099 20440
rect 10777 20435 10843 20438
rect 17033 20435 17099 20438
rect 18229 20498 18295 20501
rect 27520 20498 28000 20528
rect 18229 20496 28000 20498
rect 18229 20440 18234 20496
rect 18290 20440 28000 20496
rect 18229 20438 28000 20440
rect 18229 20435 18295 20438
rect 27520 20408 28000 20438
rect 0 20362 480 20392
rect 1485 20362 1551 20365
rect 0 20360 1551 20362
rect 0 20304 1490 20360
rect 1546 20304 1551 20360
rect 0 20302 1551 20304
rect 0 20272 480 20302
rect 1485 20299 1551 20302
rect 8753 20362 8819 20365
rect 17493 20362 17559 20365
rect 8753 20360 17559 20362
rect 8753 20304 8758 20360
rect 8814 20304 17498 20360
rect 17554 20304 17559 20360
rect 8753 20302 17559 20304
rect 8753 20299 8819 20302
rect 17493 20299 17559 20302
rect 2037 20226 2103 20229
rect 5349 20226 5415 20229
rect 2037 20224 5415 20226
rect 2037 20168 2042 20224
rect 2098 20168 5354 20224
rect 5410 20168 5415 20224
rect 2037 20166 5415 20168
rect 2037 20163 2103 20166
rect 5349 20163 5415 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 24117 19954 24183 19957
rect 27520 19954 28000 19984
rect 24117 19952 28000 19954
rect 24117 19896 24122 19952
rect 24178 19896 28000 19952
rect 24117 19894 28000 19896
rect 24117 19891 24183 19894
rect 27520 19864 28000 19894
rect 0 19682 480 19712
rect 1393 19682 1459 19685
rect 0 19680 1459 19682
rect 0 19624 1398 19680
rect 1454 19624 1459 19680
rect 0 19622 1459 19624
rect 0 19592 480 19622
rect 1393 19619 1459 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 24761 19410 24827 19413
rect 27520 19410 28000 19440
rect 24761 19408 28000 19410
rect 24761 19352 24766 19408
rect 24822 19352 28000 19408
rect 24761 19350 28000 19352
rect 24761 19347 24827 19350
rect 27520 19320 28000 19350
rect 16941 19274 17007 19277
rect 24577 19274 24643 19277
rect 16941 19272 24643 19274
rect 16941 19216 16946 19272
rect 17002 19216 24582 19272
rect 24638 19216 24643 19272
rect 16941 19214 24643 19216
rect 16941 19211 17007 19214
rect 24577 19211 24643 19214
rect 0 19138 480 19168
rect 2405 19138 2471 19141
rect 4337 19138 4403 19141
rect 0 19078 1594 19138
rect 0 19048 480 19078
rect 1534 19002 1594 19078
rect 2405 19136 4403 19138
rect 2405 19080 2410 19136
rect 2466 19080 4342 19136
rect 4398 19080 4403 19136
rect 2405 19078 4403 19080
rect 2405 19075 2471 19078
rect 4337 19075 4403 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2865 19002 2931 19005
rect 1534 19000 2931 19002
rect 1534 18944 2870 19000
rect 2926 18944 2931 19000
rect 1534 18942 2931 18944
rect 2865 18939 2931 18942
rect 20118 18942 24962 19002
rect 15561 18866 15627 18869
rect 20118 18866 20178 18942
rect 15561 18864 20178 18866
rect 15561 18808 15566 18864
rect 15622 18808 20178 18864
rect 15561 18806 20178 18808
rect 15561 18803 15627 18806
rect 19057 18730 19123 18733
rect 24393 18730 24459 18733
rect 19057 18728 24459 18730
rect 19057 18672 19062 18728
rect 19118 18672 24398 18728
rect 24454 18672 24459 18728
rect 19057 18670 24459 18672
rect 24902 18730 24962 18942
rect 27520 18730 28000 18760
rect 24902 18670 28000 18730
rect 19057 18667 19123 18670
rect 24393 18667 24459 18670
rect 27520 18640 28000 18670
rect 0 18594 480 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 480 18534
rect 1577 18531 1643 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 12617 18322 12683 18325
rect 24577 18322 24643 18325
rect 12617 18320 24643 18322
rect 12617 18264 12622 18320
rect 12678 18264 24582 18320
rect 24638 18264 24643 18320
rect 12617 18262 24643 18264
rect 12617 18259 12683 18262
rect 24577 18259 24643 18262
rect 24761 18186 24827 18189
rect 27520 18186 28000 18216
rect 24761 18184 28000 18186
rect 24761 18128 24766 18184
rect 24822 18128 28000 18184
rect 24761 18126 28000 18128
rect 24761 18123 24827 18126
rect 27520 18096 28000 18126
rect 0 18050 480 18080
rect 4245 18050 4311 18053
rect 0 18048 4311 18050
rect 0 17992 4250 18048
rect 4306 17992 4311 18048
rect 0 17990 4311 17992
rect 0 17960 480 17990
rect 4245 17987 4311 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 11881 17778 11947 17781
rect 21265 17778 21331 17781
rect 11881 17776 21331 17778
rect 11881 17720 11886 17776
rect 11942 17720 21270 17776
rect 21326 17720 21331 17776
rect 11881 17718 21331 17720
rect 11881 17715 11947 17718
rect 21265 17715 21331 17718
rect 19977 17642 20043 17645
rect 27520 17642 28000 17672
rect 19977 17640 28000 17642
rect 19977 17584 19982 17640
rect 20038 17584 28000 17640
rect 19977 17582 28000 17584
rect 19977 17579 20043 17582
rect 27520 17552 28000 17582
rect 0 17506 480 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 480 17446
rect 2773 17443 2839 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 2773 17098 2839 17101
rect 5257 17098 5323 17101
rect 2773 17096 5323 17098
rect 2773 17040 2778 17096
rect 2834 17040 5262 17096
rect 5318 17040 5323 17096
rect 2773 17038 5323 17040
rect 2773 17035 2839 17038
rect 5257 17035 5323 17038
rect 23657 17098 23723 17101
rect 27520 17098 28000 17128
rect 23657 17096 28000 17098
rect 23657 17040 23662 17096
rect 23718 17040 28000 17096
rect 23657 17038 28000 17040
rect 23657 17035 23723 17038
rect 27520 17008 28000 17038
rect 22461 16962 22527 16965
rect 24945 16962 25011 16965
rect 22461 16960 25011 16962
rect 22461 16904 22466 16960
rect 22522 16904 24950 16960
rect 25006 16904 25011 16960
rect 22461 16902 25011 16904
rect 22461 16899 22527 16902
rect 24945 16899 25011 16902
rect 10277 16896 10597 16897
rect 0 16826 480 16856
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4613 16826 4679 16829
rect 0 16824 4679 16826
rect 0 16768 4618 16824
rect 4674 16768 4679 16824
rect 0 16766 4679 16768
rect 0 16736 480 16766
rect 4613 16763 4679 16766
rect 20989 16826 21055 16829
rect 23657 16826 23723 16829
rect 20989 16824 23723 16826
rect 20989 16768 20994 16824
rect 21050 16768 23662 16824
rect 23718 16768 23723 16824
rect 20989 16766 23723 16768
rect 20989 16763 21055 16766
rect 23657 16763 23723 16766
rect 2681 16690 2747 16693
rect 3141 16690 3207 16693
rect 2681 16688 3207 16690
rect 2681 16632 2686 16688
rect 2742 16632 3146 16688
rect 3202 16632 3207 16688
rect 2681 16630 3207 16632
rect 2681 16627 2747 16630
rect 3141 16627 3207 16630
rect 13169 16690 13235 16693
rect 20713 16690 20779 16693
rect 13169 16688 20779 16690
rect 13169 16632 13174 16688
rect 13230 16632 20718 16688
rect 20774 16632 20779 16688
rect 13169 16630 20779 16632
rect 13169 16627 13235 16630
rect 20713 16627 20779 16630
rect 22645 16690 22711 16693
rect 24485 16690 24551 16693
rect 22645 16688 24551 16690
rect 22645 16632 22650 16688
rect 22706 16632 24490 16688
rect 24546 16632 24551 16688
rect 22645 16630 24551 16632
rect 22645 16627 22711 16630
rect 24485 16627 24551 16630
rect 2037 16556 2103 16557
rect 2037 16554 2084 16556
rect 1992 16552 2084 16554
rect 2148 16554 2154 16556
rect 2865 16554 2931 16557
rect 2148 16552 2931 16554
rect 1992 16496 2042 16552
rect 2148 16496 2870 16552
rect 2926 16496 2931 16552
rect 1992 16494 2084 16496
rect 2037 16492 2084 16494
rect 2148 16494 2931 16496
rect 2148 16492 2154 16494
rect 2037 16491 2103 16492
rect 2865 16491 2931 16494
rect 3969 16554 4035 16557
rect 7097 16554 7163 16557
rect 3969 16552 7163 16554
rect 3969 16496 3974 16552
rect 4030 16496 7102 16552
rect 7158 16496 7163 16552
rect 3969 16494 7163 16496
rect 3969 16491 4035 16494
rect 7097 16491 7163 16494
rect 23473 16554 23539 16557
rect 27520 16554 28000 16584
rect 23473 16552 28000 16554
rect 23473 16496 23478 16552
rect 23534 16496 28000 16552
rect 23473 16494 28000 16496
rect 23473 16491 23539 16494
rect 27520 16464 28000 16494
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 480 16222
rect 4061 16219 4127 16222
rect 10133 16146 10199 16149
rect 2454 16144 10199 16146
rect 2454 16088 10138 16144
rect 10194 16088 10199 16144
rect 2454 16086 10199 16088
rect 0 15738 480 15768
rect 2454 15738 2514 16086
rect 10133 16083 10199 16086
rect 4153 16010 4219 16013
rect 6494 16010 6500 16012
rect 4153 16008 6500 16010
rect 4153 15952 4158 16008
rect 4214 15952 6500 16008
rect 4153 15950 6500 15952
rect 4153 15947 4219 15950
rect 6494 15948 6500 15950
rect 6564 15948 6570 16012
rect 8477 16010 8543 16013
rect 21725 16010 21791 16013
rect 23749 16010 23815 16013
rect 6686 16008 23815 16010
rect 6686 15952 8482 16008
rect 8538 15952 21730 16008
rect 21786 15952 23754 16008
rect 23810 15952 23815 16008
rect 6686 15950 23815 15952
rect 4337 15874 4403 15877
rect 6686 15874 6746 15950
rect 8477 15947 8543 15950
rect 21725 15947 21791 15950
rect 23749 15947 23815 15950
rect 24025 16010 24091 16013
rect 27520 16010 28000 16040
rect 24025 16008 28000 16010
rect 24025 15952 24030 16008
rect 24086 15952 28000 16008
rect 24025 15950 28000 15952
rect 24025 15947 24091 15950
rect 27520 15920 28000 15950
rect 4337 15872 6746 15874
rect 4337 15816 4342 15872
rect 4398 15816 6746 15872
rect 4337 15814 6746 15816
rect 13537 15874 13603 15877
rect 22093 15874 22159 15877
rect 25037 15874 25103 15877
rect 13537 15872 18154 15874
rect 13537 15816 13542 15872
rect 13598 15816 18154 15872
rect 13537 15814 18154 15816
rect 4337 15811 4403 15814
rect 13537 15811 13603 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 0 15678 2514 15738
rect 2865 15738 2931 15741
rect 12433 15738 12499 15741
rect 15377 15738 15443 15741
rect 2865 15736 7850 15738
rect 2865 15680 2870 15736
rect 2926 15680 7850 15736
rect 2865 15678 7850 15680
rect 0 15648 480 15678
rect 2865 15675 2931 15678
rect 2405 15602 2471 15605
rect 7005 15602 7071 15605
rect 2405 15600 7071 15602
rect 2405 15544 2410 15600
rect 2466 15544 7010 15600
rect 7066 15544 7071 15600
rect 2405 15542 7071 15544
rect 7790 15602 7850 15678
rect 12433 15736 15443 15738
rect 12433 15680 12438 15736
rect 12494 15680 15382 15736
rect 15438 15680 15443 15736
rect 12433 15678 15443 15680
rect 12433 15675 12499 15678
rect 15377 15675 15443 15678
rect 13445 15602 13511 15605
rect 17953 15602 18019 15605
rect 7790 15600 18019 15602
rect 7790 15544 13450 15600
rect 13506 15544 17958 15600
rect 18014 15544 18019 15600
rect 7790 15542 18019 15544
rect 18094 15602 18154 15814
rect 22093 15872 25103 15874
rect 22093 15816 22098 15872
rect 22154 15816 25042 15872
rect 25098 15816 25103 15872
rect 22093 15814 25103 15816
rect 22093 15811 22159 15814
rect 25037 15811 25103 15814
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 24669 15602 24735 15605
rect 18094 15600 24735 15602
rect 18094 15544 24674 15600
rect 24730 15544 24735 15600
rect 18094 15542 24735 15544
rect 2405 15539 2471 15542
rect 7005 15539 7071 15542
rect 13445 15539 13511 15542
rect 17953 15539 18019 15542
rect 24669 15539 24735 15542
rect 1853 15466 1919 15469
rect 5533 15466 5599 15469
rect 1853 15464 5599 15466
rect 1853 15408 1858 15464
rect 1914 15408 5538 15464
rect 5594 15408 5599 15464
rect 1853 15406 5599 15408
rect 1853 15403 1919 15406
rect 5533 15403 5599 15406
rect 9489 15466 9555 15469
rect 15009 15466 15075 15469
rect 9489 15464 15075 15466
rect 9489 15408 9494 15464
rect 9550 15408 15014 15464
rect 15070 15408 15075 15464
rect 9489 15406 15075 15408
rect 9489 15403 9555 15406
rect 15009 15403 15075 15406
rect 22001 15466 22067 15469
rect 27520 15466 28000 15496
rect 22001 15464 28000 15466
rect 22001 15408 22006 15464
rect 22062 15408 28000 15464
rect 22001 15406 28000 15408
rect 22001 15403 22067 15406
rect 27520 15376 28000 15406
rect 4286 15268 4292 15332
rect 4356 15330 4362 15332
rect 4521 15330 4587 15333
rect 4356 15328 4587 15330
rect 4356 15272 4526 15328
rect 4582 15272 4587 15328
rect 4356 15270 4587 15272
rect 4356 15268 4362 15270
rect 4521 15267 4587 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 20437 15194 20503 15197
rect 20621 15194 20687 15197
rect 23841 15194 23907 15197
rect 0 15134 2698 15194
rect 0 15104 480 15134
rect 2638 15058 2698 15134
rect 20437 15192 23907 15194
rect 20437 15136 20442 15192
rect 20498 15136 20626 15192
rect 20682 15136 23846 15192
rect 23902 15136 23907 15192
rect 20437 15134 23907 15136
rect 20437 15131 20503 15134
rect 20621 15131 20687 15134
rect 23841 15131 23907 15134
rect 18965 15058 19031 15061
rect 25773 15058 25839 15061
rect 2638 15024 2744 15058
rect 2822 15024 18890 15058
rect 2638 14998 18890 15024
rect 2684 14964 2882 14998
rect 3233 14922 3299 14925
rect 15469 14922 15535 14925
rect 3233 14920 15535 14922
rect 3233 14864 3238 14920
rect 3294 14864 15474 14920
rect 15530 14864 15535 14920
rect 3233 14862 15535 14864
rect 18830 14922 18890 14998
rect 18965 15056 25839 15058
rect 18965 15000 18970 15056
rect 19026 15000 25778 15056
rect 25834 15000 25839 15056
rect 18965 14998 25839 15000
rect 18965 14995 19031 14998
rect 25773 14995 25839 14998
rect 21173 14922 21239 14925
rect 21541 14922 21607 14925
rect 18830 14920 21607 14922
rect 18830 14864 21178 14920
rect 21234 14864 21546 14920
rect 21602 14864 21607 14920
rect 18830 14862 21607 14864
rect 3233 14859 3299 14862
rect 15469 14859 15535 14862
rect 21173 14859 21239 14862
rect 21541 14859 21607 14862
rect 23749 14922 23815 14925
rect 27520 14922 28000 14952
rect 23749 14920 28000 14922
rect 23749 14864 23754 14920
rect 23810 14864 28000 14920
rect 23749 14862 28000 14864
rect 23749 14859 23815 14862
rect 27520 14832 28000 14862
rect 14641 14786 14707 14789
rect 15653 14786 15719 14789
rect 19425 14788 19491 14789
rect 14641 14784 15719 14786
rect 14641 14728 14646 14784
rect 14702 14728 15658 14784
rect 15714 14728 15719 14784
rect 14641 14726 15719 14728
rect 14641 14723 14707 14726
rect 15653 14723 15719 14726
rect 19374 14724 19380 14788
rect 19444 14786 19491 14788
rect 22737 14786 22803 14789
rect 25221 14786 25287 14789
rect 19444 14784 19536 14786
rect 19486 14728 19536 14784
rect 19444 14726 19536 14728
rect 22737 14784 25287 14786
rect 22737 14728 22742 14784
rect 22798 14728 25226 14784
rect 25282 14728 25287 14784
rect 22737 14726 25287 14728
rect 19444 14724 19491 14726
rect 19425 14723 19491 14724
rect 22737 14723 22803 14726
rect 25221 14723 25287 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3969 14650 4035 14653
rect 0 14648 4035 14650
rect 0 14592 3974 14648
rect 4030 14592 4035 14648
rect 0 14590 4035 14592
rect 0 14560 480 14590
rect 3969 14587 4035 14590
rect 14406 14588 14412 14652
rect 14476 14650 14482 14652
rect 15009 14650 15075 14653
rect 19057 14650 19123 14653
rect 23473 14652 23539 14653
rect 14476 14648 19123 14650
rect 14476 14592 15014 14648
rect 15070 14592 19062 14648
rect 19118 14592 19123 14648
rect 14476 14590 19123 14592
rect 14476 14588 14482 14590
rect 15009 14587 15075 14590
rect 19057 14587 19123 14590
rect 23422 14588 23428 14652
rect 23492 14650 23539 14652
rect 23492 14648 23584 14650
rect 23534 14592 23584 14648
rect 23492 14590 23584 14592
rect 23492 14588 23539 14590
rect 23473 14587 23539 14588
rect 18781 14514 18847 14517
rect 21449 14514 21515 14517
rect 23013 14516 23079 14517
rect 23013 14514 23060 14516
rect 18781 14512 21515 14514
rect 18781 14456 18786 14512
rect 18842 14456 21454 14512
rect 21510 14456 21515 14512
rect 18781 14454 21515 14456
rect 22968 14512 23060 14514
rect 22968 14456 23018 14512
rect 22968 14454 23060 14456
rect 18781 14451 18847 14454
rect 21449 14451 21515 14454
rect 23013 14452 23060 14454
rect 23124 14452 23130 14516
rect 23013 14451 23079 14452
rect 5441 14378 5507 14381
rect 8569 14378 8635 14381
rect 15009 14378 15075 14381
rect 15745 14378 15811 14381
rect 5441 14376 6148 14378
rect 5441 14320 5446 14376
rect 5502 14320 6148 14376
rect 5441 14318 6148 14320
rect 5441 14315 5507 14318
rect 6088 14242 6148 14318
rect 8569 14376 15811 14378
rect 8569 14320 8574 14376
rect 8630 14320 15014 14376
rect 15070 14320 15750 14376
rect 15806 14320 15811 14376
rect 8569 14318 15811 14320
rect 8569 14315 8635 14318
rect 15009 14315 15075 14318
rect 15745 14315 15811 14318
rect 20529 14378 20595 14381
rect 27520 14378 28000 14408
rect 20529 14376 28000 14378
rect 20529 14320 20534 14376
rect 20590 14320 28000 14376
rect 20529 14318 28000 14320
rect 20529 14315 20595 14318
rect 27520 14288 28000 14318
rect 6729 14242 6795 14245
rect 14733 14242 14799 14245
rect 6088 14240 14799 14242
rect 6088 14184 6734 14240
rect 6790 14184 14738 14240
rect 14794 14184 14799 14240
rect 6088 14182 14799 14184
rect 6729 14179 6795 14182
rect 14733 14179 14799 14182
rect 17033 14242 17099 14245
rect 18045 14242 18111 14245
rect 17033 14240 18111 14242
rect 17033 14184 17038 14240
rect 17094 14184 18050 14240
rect 18106 14184 18111 14240
rect 17033 14182 18111 14184
rect 17033 14179 17099 14182
rect 18045 14179 18111 14182
rect 18321 14242 18387 14245
rect 18321 14240 24042 14242
rect 18321 14184 18326 14240
rect 18382 14184 24042 14240
rect 18321 14182 24042 14184
rect 18321 14179 18387 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 2221 14106 2287 14109
rect 4889 14106 4955 14109
rect 2221 14104 4955 14106
rect 2221 14048 2226 14104
rect 2282 14048 4894 14104
rect 4950 14048 4955 14104
rect 2221 14046 4955 14048
rect 2221 14043 2287 14046
rect 4889 14043 4955 14046
rect 16205 14106 16271 14109
rect 16205 14104 19442 14106
rect 16205 14048 16210 14104
rect 16266 14048 19442 14104
rect 16205 14046 19442 14048
rect 16205 14043 16271 14046
rect 0 13970 480 14000
rect 3233 13970 3299 13973
rect 0 13968 3299 13970
rect 0 13912 3238 13968
rect 3294 13912 3299 13968
rect 0 13910 3299 13912
rect 0 13880 480 13910
rect 3233 13907 3299 13910
rect 3969 13970 4035 13973
rect 15101 13970 15167 13973
rect 3969 13968 15167 13970
rect 3969 13912 3974 13968
rect 4030 13912 15106 13968
rect 15162 13912 15167 13968
rect 3969 13910 15167 13912
rect 3969 13907 4035 13910
rect 15101 13907 15167 13910
rect 15285 13970 15351 13973
rect 18045 13970 18111 13973
rect 15285 13968 18111 13970
rect 15285 13912 15290 13968
rect 15346 13912 18050 13968
rect 18106 13912 18111 13968
rect 15285 13910 18111 13912
rect 15285 13907 15351 13910
rect 18045 13907 18111 13910
rect 19382 13837 19442 14046
rect 23982 13970 24042 14182
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 25037 13970 25103 13973
rect 23982 13968 25103 13970
rect 23982 13912 25042 13968
rect 25098 13912 25103 13968
rect 23982 13910 25103 13912
rect 25037 13907 25103 13910
rect 1945 13834 2011 13837
rect 3049 13834 3115 13837
rect 3877 13834 3943 13837
rect 1945 13832 3943 13834
rect 1945 13776 1950 13832
rect 2006 13776 3054 13832
rect 3110 13776 3882 13832
rect 3938 13776 3943 13832
rect 1945 13774 3943 13776
rect 1945 13771 2011 13774
rect 3049 13771 3115 13774
rect 3877 13771 3943 13774
rect 7966 13772 7972 13836
rect 8036 13834 8042 13836
rect 8201 13834 8267 13837
rect 8036 13832 8267 13834
rect 8036 13776 8206 13832
rect 8262 13776 8267 13832
rect 8036 13774 8267 13776
rect 8036 13772 8042 13774
rect 8201 13771 8267 13774
rect 10685 13834 10751 13837
rect 17217 13834 17283 13837
rect 10685 13832 17283 13834
rect 10685 13776 10690 13832
rect 10746 13776 17222 13832
rect 17278 13776 17283 13832
rect 10685 13774 17283 13776
rect 19382 13832 19491 13837
rect 19382 13776 19430 13832
rect 19486 13776 19491 13832
rect 19382 13774 19491 13776
rect 10685 13771 10751 13774
rect 17217 13771 17283 13774
rect 19425 13771 19491 13774
rect 20161 13834 20227 13837
rect 23657 13834 23723 13837
rect 20161 13832 23723 13834
rect 20161 13776 20166 13832
rect 20222 13776 23662 13832
rect 23718 13776 23723 13832
rect 20161 13774 23723 13776
rect 20161 13771 20227 13774
rect 23657 13771 23723 13774
rect 3877 13698 3943 13701
rect 8017 13698 8083 13701
rect 9765 13698 9831 13701
rect 3877 13696 9831 13698
rect 3877 13640 3882 13696
rect 3938 13640 8022 13696
rect 8078 13640 9770 13696
rect 9826 13640 9831 13696
rect 3877 13638 9831 13640
rect 3877 13635 3943 13638
rect 8017 13635 8083 13638
rect 9765 13635 9831 13638
rect 20437 13698 20503 13701
rect 24761 13698 24827 13701
rect 27520 13698 28000 13728
rect 20437 13696 24827 13698
rect 20437 13640 20442 13696
rect 20498 13640 24766 13696
rect 24822 13640 24827 13696
rect 20437 13638 24827 13640
rect 20437 13635 20503 13638
rect 24761 13635 24827 13638
rect 24902 13638 28000 13698
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 13721 13562 13787 13565
rect 15929 13562 15995 13565
rect 13721 13560 15995 13562
rect 13721 13504 13726 13560
rect 13782 13504 15934 13560
rect 15990 13504 15995 13560
rect 13721 13502 15995 13504
rect 13721 13499 13787 13502
rect 15929 13499 15995 13502
rect 23606 13500 23612 13564
rect 23676 13562 23682 13564
rect 23841 13562 23907 13565
rect 23676 13560 23907 13562
rect 23676 13504 23846 13560
rect 23902 13504 23907 13560
rect 23676 13502 23907 13504
rect 23676 13500 23682 13502
rect 23841 13499 23907 13502
rect 0 13426 480 13456
rect 6177 13426 6243 13429
rect 12525 13426 12591 13429
rect 17217 13426 17283 13429
rect 24902 13426 24962 13638
rect 27520 13608 28000 13638
rect 0 13366 6010 13426
rect 0 13336 480 13366
rect 1945 13290 2011 13293
rect 3693 13290 3759 13293
rect 1945 13288 3759 13290
rect 1945 13232 1950 13288
rect 2006 13232 3698 13288
rect 3754 13232 3759 13288
rect 1945 13230 3759 13232
rect 5950 13290 6010 13366
rect 6177 13424 12591 13426
rect 6177 13368 6182 13424
rect 6238 13368 12530 13424
rect 12586 13368 12591 13424
rect 6177 13366 12591 13368
rect 6177 13363 6243 13366
rect 12525 13363 12591 13366
rect 14644 13424 24962 13426
rect 14644 13368 17222 13424
rect 17278 13368 24962 13424
rect 14644 13366 24962 13368
rect 9949 13290 10015 13293
rect 5950 13288 10015 13290
rect 5950 13232 9954 13288
rect 10010 13232 10015 13288
rect 5950 13230 10015 13232
rect 1945 13227 2011 13230
rect 3693 13227 3759 13230
rect 9949 13227 10015 13230
rect 9765 13154 9831 13157
rect 14644 13154 14704 13366
rect 17217 13363 17283 13366
rect 16021 13290 16087 13293
rect 9765 13152 14704 13154
rect 9765 13096 9770 13152
rect 9826 13096 14704 13152
rect 9765 13094 14704 13096
rect 14782 13288 16087 13290
rect 14782 13232 16026 13288
rect 16082 13232 16087 13288
rect 14782 13230 16087 13232
rect 9765 13091 9831 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 2957 13020 3023 13021
rect 2957 13018 3004 13020
rect 2912 13016 3004 13018
rect 2912 12960 2962 13016
rect 2912 12958 3004 12960
rect 2957 12956 3004 12958
rect 3068 12956 3074 13020
rect 6637 13018 6703 13021
rect 9581 13018 9647 13021
rect 14782 13018 14842 13230
rect 16021 13227 16087 13230
rect 18505 13290 18571 13293
rect 25313 13290 25379 13293
rect 18505 13288 25379 13290
rect 18505 13232 18510 13288
rect 18566 13232 25318 13288
rect 25374 13232 25379 13288
rect 18505 13230 25379 13232
rect 18505 13227 18571 13230
rect 25313 13227 25379 13230
rect 16205 13154 16271 13157
rect 22921 13154 22987 13157
rect 16205 13152 22987 13154
rect 16205 13096 16210 13152
rect 16266 13096 22926 13152
rect 22982 13096 22987 13152
rect 16205 13094 22987 13096
rect 16205 13091 16271 13094
rect 22921 13091 22987 13094
rect 24669 13154 24735 13157
rect 27520 13154 28000 13184
rect 24669 13152 28000 13154
rect 24669 13096 24674 13152
rect 24730 13096 28000 13152
rect 24669 13094 28000 13096
rect 24669 13091 24735 13094
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 20253 13018 20319 13021
rect 6637 13016 14842 13018
rect 6637 12960 6642 13016
rect 6698 12960 9586 13016
rect 9642 12960 14842 13016
rect 6637 12958 14842 12960
rect 16254 13016 20319 13018
rect 16254 12960 20258 13016
rect 20314 12960 20319 13016
rect 16254 12958 20319 12960
rect 2957 12955 3023 12956
rect 6637 12955 6703 12958
rect 9581 12955 9647 12958
rect 0 12882 480 12912
rect 6913 12882 6979 12885
rect 11697 12882 11763 12885
rect 0 12822 6746 12882
rect 0 12792 480 12822
rect 2313 12746 2379 12749
rect 3141 12746 3207 12749
rect 2313 12744 3207 12746
rect 2313 12688 2318 12744
rect 2374 12688 3146 12744
rect 3202 12688 3207 12744
rect 2313 12686 3207 12688
rect 2313 12683 2379 12686
rect 3141 12683 3207 12686
rect 3601 12746 3667 12749
rect 4337 12746 4403 12749
rect 3601 12744 4403 12746
rect 3601 12688 3606 12744
rect 3662 12688 4342 12744
rect 4398 12688 4403 12744
rect 3601 12686 4403 12688
rect 3601 12683 3667 12686
rect 4337 12683 4403 12686
rect 3969 12610 4035 12613
rect 6453 12610 6519 12613
rect 3969 12608 6519 12610
rect 3969 12552 3974 12608
rect 4030 12552 6458 12608
rect 6514 12552 6519 12608
rect 3969 12550 6519 12552
rect 3969 12547 4035 12550
rect 6453 12547 6519 12550
rect 2313 12474 2379 12477
rect 6545 12474 6611 12477
rect 2313 12472 6611 12474
rect 2313 12416 2318 12472
rect 2374 12416 6550 12472
rect 6606 12416 6611 12472
rect 2313 12414 6611 12416
rect 6686 12474 6746 12822
rect 6913 12880 11763 12882
rect 6913 12824 6918 12880
rect 6974 12824 11702 12880
rect 11758 12824 11763 12880
rect 6913 12822 11763 12824
rect 6913 12819 6979 12822
rect 11697 12819 11763 12822
rect 13854 12820 13860 12884
rect 13924 12882 13930 12884
rect 15469 12882 15535 12885
rect 13924 12880 15535 12882
rect 13924 12824 15474 12880
rect 15530 12824 15535 12880
rect 13924 12822 15535 12824
rect 13924 12820 13930 12822
rect 15469 12819 15535 12822
rect 6821 12746 6887 12749
rect 16254 12746 16314 12958
rect 20253 12955 20319 12958
rect 18965 12882 19031 12885
rect 20897 12882 20963 12885
rect 18965 12880 20963 12882
rect 18965 12824 18970 12880
rect 19026 12824 20902 12880
rect 20958 12824 20963 12880
rect 18965 12822 20963 12824
rect 18965 12819 19031 12822
rect 20897 12819 20963 12822
rect 6821 12744 16314 12746
rect 6821 12688 6826 12744
rect 6882 12688 16314 12744
rect 6821 12686 16314 12688
rect 16389 12746 16455 12749
rect 20478 12746 20484 12748
rect 16389 12744 20484 12746
rect 16389 12688 16394 12744
rect 16450 12688 20484 12744
rect 16389 12686 20484 12688
rect 6821 12683 6887 12686
rect 16389 12683 16455 12686
rect 20478 12684 20484 12686
rect 20548 12684 20554 12748
rect 15101 12610 15167 12613
rect 16757 12610 16823 12613
rect 15101 12608 16823 12610
rect 15101 12552 15106 12608
rect 15162 12552 16762 12608
rect 16818 12552 16823 12608
rect 15101 12550 16823 12552
rect 15101 12547 15167 12550
rect 16757 12547 16823 12550
rect 20161 12610 20227 12613
rect 23013 12610 23079 12613
rect 20161 12608 23079 12610
rect 20161 12552 20166 12608
rect 20222 12552 23018 12608
rect 23074 12552 23079 12608
rect 20161 12550 23079 12552
rect 20161 12547 20227 12550
rect 23013 12547 23079 12550
rect 23790 12548 23796 12612
rect 23860 12610 23866 12612
rect 27520 12610 28000 12640
rect 23860 12550 28000 12610
rect 23860 12548 23866 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 11697 12474 11763 12477
rect 20437 12474 20503 12477
rect 23657 12474 23723 12477
rect 6686 12414 10196 12474
rect 2313 12411 2379 12414
rect 6545 12411 6611 12414
rect 0 12338 480 12368
rect 3918 12338 3924 12340
rect 0 12278 3924 12338
rect 0 12248 480 12278
rect 3918 12276 3924 12278
rect 3988 12276 3994 12340
rect 4153 12338 4219 12341
rect 6085 12338 6151 12341
rect 4153 12336 6151 12338
rect 4153 12280 4158 12336
rect 4214 12280 6090 12336
rect 6146 12280 6151 12336
rect 4153 12278 6151 12280
rect 10136 12338 10196 12414
rect 11697 12472 12818 12474
rect 11697 12416 11702 12472
rect 11758 12416 12818 12472
rect 11697 12414 12818 12416
rect 11697 12411 11763 12414
rect 11605 12338 11671 12341
rect 10136 12336 11671 12338
rect 10136 12280 11610 12336
rect 11666 12280 11671 12336
rect 10136 12278 11671 12280
rect 12758 12338 12818 12414
rect 20437 12472 23723 12474
rect 20437 12416 20442 12472
rect 20498 12416 23662 12472
rect 23718 12416 23723 12472
rect 20437 12414 23723 12416
rect 20437 12411 20503 12414
rect 23657 12411 23723 12414
rect 23289 12338 23355 12341
rect 12758 12336 23355 12338
rect 12758 12280 23294 12336
rect 23350 12280 23355 12336
rect 12758 12278 23355 12280
rect 4153 12275 4219 12278
rect 6085 12275 6151 12278
rect 11605 12275 11671 12278
rect 23289 12275 23355 12278
rect 23657 12338 23723 12341
rect 23790 12338 23796 12340
rect 23657 12336 23796 12338
rect 23657 12280 23662 12336
rect 23718 12280 23796 12336
rect 23657 12278 23796 12280
rect 23657 12275 23723 12278
rect 23790 12276 23796 12278
rect 23860 12276 23866 12340
rect 2221 12202 2287 12205
rect 6913 12202 6979 12205
rect 2221 12200 6979 12202
rect 2221 12144 2226 12200
rect 2282 12144 6918 12200
rect 6974 12144 6979 12200
rect 2221 12142 6979 12144
rect 2221 12139 2287 12142
rect 6913 12139 6979 12142
rect 16389 12202 16455 12205
rect 16573 12202 16639 12205
rect 17125 12202 17191 12205
rect 17953 12202 18019 12205
rect 19977 12202 20043 12205
rect 16389 12200 20043 12202
rect 16389 12144 16394 12200
rect 16450 12144 16578 12200
rect 16634 12144 17130 12200
rect 17186 12144 17958 12200
rect 18014 12144 19982 12200
rect 20038 12144 20043 12200
rect 16389 12142 20043 12144
rect 16389 12139 16455 12142
rect 16573 12139 16639 12142
rect 17125 12139 17191 12142
rect 17953 12139 18019 12142
rect 19977 12139 20043 12142
rect 23974 12140 23980 12204
rect 24044 12202 24050 12204
rect 24044 12142 24778 12202
rect 24044 12140 24050 12142
rect 3049 12068 3115 12069
rect 2998 12004 3004 12068
rect 3068 12066 3115 12068
rect 15929 12066 15995 12069
rect 21081 12066 21147 12069
rect 3068 12064 3160 12066
rect 3110 12008 3160 12064
rect 3068 12006 3160 12008
rect 15929 12064 21147 12066
rect 15929 12008 15934 12064
rect 15990 12008 21086 12064
rect 21142 12008 21147 12064
rect 15929 12006 21147 12008
rect 24718 12066 24778 12142
rect 27520 12066 28000 12096
rect 24718 12006 28000 12066
rect 3068 12004 3115 12006
rect 3049 12003 3115 12004
rect 15929 12003 15995 12006
rect 21081 12003 21147 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 27520 11976 28000 12006
rect 24277 11935 24597 11936
rect 2221 11930 2287 11933
rect 3509 11930 3575 11933
rect 2221 11928 3575 11930
rect 2221 11872 2226 11928
rect 2282 11872 3514 11928
rect 3570 11872 3575 11928
rect 2221 11870 3575 11872
rect 2221 11867 2287 11870
rect 3509 11867 3575 11870
rect 4705 11928 4771 11933
rect 4705 11872 4710 11928
rect 4766 11872 4771 11928
rect 4705 11867 4771 11872
rect 17769 11930 17835 11933
rect 19333 11930 19399 11933
rect 17769 11928 19399 11930
rect 17769 11872 17774 11928
rect 17830 11872 19338 11928
rect 19394 11872 19399 11928
rect 17769 11870 19399 11872
rect 17769 11867 17835 11870
rect 19333 11867 19399 11870
rect 0 11794 480 11824
rect 3785 11794 3851 11797
rect 0 11792 3851 11794
rect 0 11736 3790 11792
rect 3846 11736 3851 11792
rect 0 11734 3851 11736
rect 0 11704 480 11734
rect 3785 11731 3851 11734
rect 4521 11794 4587 11797
rect 4708 11794 4768 11867
rect 4521 11792 4768 11794
rect 4521 11736 4526 11792
rect 4582 11736 4768 11792
rect 4521 11734 4768 11736
rect 8201 11794 8267 11797
rect 12433 11794 12499 11797
rect 8201 11792 12499 11794
rect 8201 11736 8206 11792
rect 8262 11736 12438 11792
rect 12494 11736 12499 11792
rect 8201 11734 12499 11736
rect 4521 11731 4587 11734
rect 8201 11731 8267 11734
rect 12433 11731 12499 11734
rect 13169 11794 13235 11797
rect 17125 11794 17191 11797
rect 25313 11794 25379 11797
rect 13169 11792 16636 11794
rect 13169 11736 13174 11792
rect 13230 11736 16636 11792
rect 13169 11734 16636 11736
rect 13169 11731 13235 11734
rect 1761 11658 1827 11661
rect 5993 11658 6059 11661
rect 1761 11656 6059 11658
rect 1761 11600 1766 11656
rect 1822 11600 5998 11656
rect 6054 11600 6059 11656
rect 1761 11598 6059 11600
rect 1761 11595 1827 11598
rect 5993 11595 6059 11598
rect 7373 11658 7439 11661
rect 8753 11658 8819 11661
rect 12525 11658 12591 11661
rect 7373 11656 12591 11658
rect 7373 11600 7378 11656
rect 7434 11600 8758 11656
rect 8814 11600 12530 11656
rect 12586 11600 12591 11656
rect 7373 11598 12591 11600
rect 7373 11595 7439 11598
rect 8753 11595 8819 11598
rect 12525 11595 12591 11598
rect 14917 11658 14983 11661
rect 16389 11658 16455 11661
rect 14917 11656 16455 11658
rect 14917 11600 14922 11656
rect 14978 11600 16394 11656
rect 16450 11600 16455 11656
rect 14917 11598 16455 11600
rect 16576 11658 16636 11734
rect 17125 11792 25379 11794
rect 17125 11736 17130 11792
rect 17186 11736 25318 11792
rect 25374 11736 25379 11792
rect 17125 11734 25379 11736
rect 17125 11731 17191 11734
rect 25313 11731 25379 11734
rect 16576 11598 24962 11658
rect 14917 11595 14983 11598
rect 16389 11595 16455 11598
rect 2129 11524 2195 11525
rect 2078 11522 2084 11524
rect 2038 11462 2084 11522
rect 2148 11520 2195 11524
rect 2190 11464 2195 11520
rect 2078 11460 2084 11462
rect 2148 11460 2195 11464
rect 2129 11459 2195 11460
rect 10869 11522 10935 11525
rect 17125 11522 17191 11525
rect 10869 11520 17191 11522
rect 10869 11464 10874 11520
rect 10930 11464 17130 11520
rect 17186 11464 17191 11520
rect 10869 11462 17191 11464
rect 24902 11522 24962 11598
rect 27520 11522 28000 11552
rect 24902 11462 28000 11522
rect 10869 11459 10935 11462
rect 17125 11459 17191 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 27520 11432 28000 11462
rect 19610 11391 19930 11392
rect 1577 11386 1643 11389
rect 2221 11386 2287 11389
rect 1577 11384 2287 11386
rect 1577 11328 1582 11384
rect 1638 11328 2226 11384
rect 2282 11328 2287 11384
rect 1577 11326 2287 11328
rect 1577 11323 1643 11326
rect 2221 11323 2287 11326
rect 3877 11386 3943 11389
rect 9581 11386 9647 11389
rect 3877 11384 9647 11386
rect 3877 11328 3882 11384
rect 3938 11328 9586 11384
rect 9642 11328 9647 11384
rect 3877 11326 9647 11328
rect 3877 11323 3943 11326
rect 9581 11323 9647 11326
rect 10777 11386 10843 11389
rect 16021 11386 16087 11389
rect 10777 11384 16087 11386
rect 10777 11328 10782 11384
rect 10838 11328 16026 11384
rect 16082 11328 16087 11384
rect 10777 11326 16087 11328
rect 10777 11323 10843 11326
rect 16021 11323 16087 11326
rect 3877 11250 3943 11253
rect 7097 11250 7163 11253
rect 3877 11248 7163 11250
rect 3877 11192 3882 11248
rect 3938 11192 7102 11248
rect 7158 11192 7163 11248
rect 3877 11190 7163 11192
rect 3877 11187 3943 11190
rect 7097 11187 7163 11190
rect 8109 11250 8175 11253
rect 8937 11250 9003 11253
rect 13445 11250 13511 11253
rect 24761 11250 24827 11253
rect 8109 11248 24827 11250
rect 8109 11192 8114 11248
rect 8170 11192 8942 11248
rect 8998 11192 13450 11248
rect 13506 11192 24766 11248
rect 24822 11192 24827 11248
rect 8109 11190 24827 11192
rect 8109 11187 8175 11190
rect 8937 11187 9003 11190
rect 13445 11187 13511 11190
rect 24761 11187 24827 11190
rect 0 11114 480 11144
rect 10317 11114 10383 11117
rect 12617 11114 12683 11117
rect 0 11112 10383 11114
rect 0 11056 10322 11112
rect 10378 11056 10383 11112
rect 0 11054 10383 11056
rect 0 11024 480 11054
rect 10317 11051 10383 11054
rect 10550 11112 12683 11114
rect 10550 11056 12622 11112
rect 12678 11056 12683 11112
rect 10550 11054 12683 11056
rect 2405 10978 2471 10981
rect 4797 10978 4863 10981
rect 2405 10976 4863 10978
rect 2405 10920 2410 10976
rect 2466 10920 4802 10976
rect 4858 10920 4863 10976
rect 2405 10918 4863 10920
rect 2405 10915 2471 10918
rect 4797 10915 4863 10918
rect 6177 10978 6243 10981
rect 9673 10978 9739 10981
rect 6177 10976 9739 10978
rect 6177 10920 6182 10976
rect 6238 10920 9678 10976
rect 9734 10920 9739 10976
rect 6177 10918 9739 10920
rect 6177 10915 6243 10918
rect 9673 10915 9739 10918
rect 9857 10978 9923 10981
rect 10550 10978 10610 11054
rect 12617 11051 12683 11054
rect 21817 11114 21883 11117
rect 22829 11114 22895 11117
rect 25497 11114 25563 11117
rect 21817 11112 22895 11114
rect 21817 11056 21822 11112
rect 21878 11056 22834 11112
rect 22890 11056 22895 11112
rect 21817 11054 22895 11056
rect 21817 11051 21883 11054
rect 22829 11051 22895 11054
rect 24028 11112 25563 11114
rect 24028 11056 25502 11112
rect 25558 11056 25563 11112
rect 24028 11054 25563 11056
rect 9857 10976 10610 10978
rect 9857 10920 9862 10976
rect 9918 10920 10610 10976
rect 9857 10918 10610 10920
rect 18965 10978 19031 10981
rect 19701 10978 19767 10981
rect 18965 10976 19767 10978
rect 18965 10920 18970 10976
rect 19026 10920 19706 10976
rect 19762 10920 19767 10976
rect 18965 10918 19767 10920
rect 9857 10915 9923 10918
rect 18965 10915 19031 10918
rect 19701 10915 19767 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 14641 10842 14707 10845
rect 6134 10840 14707 10842
rect 6134 10784 14646 10840
rect 14702 10784 14707 10840
rect 6134 10782 14707 10784
rect 3785 10706 3851 10709
rect 6134 10706 6194 10782
rect 14641 10779 14707 10782
rect 19374 10780 19380 10844
rect 19444 10842 19450 10844
rect 20345 10842 20411 10845
rect 19444 10840 20411 10842
rect 19444 10784 20350 10840
rect 20406 10784 20411 10840
rect 19444 10782 20411 10784
rect 19444 10780 19450 10782
rect 20345 10779 20411 10782
rect 20478 10780 20484 10844
rect 20548 10842 20554 10844
rect 24028 10842 24088 11054
rect 25497 11051 25563 11054
rect 27520 10978 28000 11008
rect 24718 10918 28000 10978
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 20548 10782 24088 10842
rect 20548 10780 20554 10782
rect 3785 10704 6194 10706
rect 3785 10648 3790 10704
rect 3846 10648 6194 10704
rect 3785 10646 6194 10648
rect 6637 10706 6703 10709
rect 9673 10706 9739 10709
rect 6637 10704 9739 10706
rect 6637 10648 6642 10704
rect 6698 10648 9678 10704
rect 9734 10648 9739 10704
rect 6637 10646 9739 10648
rect 3785 10643 3851 10646
rect 6637 10643 6703 10646
rect 9673 10643 9739 10646
rect 10225 10706 10291 10709
rect 13169 10706 13235 10709
rect 10225 10704 13235 10706
rect 10225 10648 10230 10704
rect 10286 10648 13174 10704
rect 13230 10648 13235 10704
rect 10225 10646 13235 10648
rect 10225 10643 10291 10646
rect 13169 10643 13235 10646
rect 13629 10706 13695 10709
rect 19517 10706 19583 10709
rect 13629 10704 19583 10706
rect 13629 10648 13634 10704
rect 13690 10648 19522 10704
rect 19578 10648 19583 10704
rect 13629 10646 19583 10648
rect 13629 10643 13695 10646
rect 19517 10643 19583 10646
rect 23974 10644 23980 10708
rect 24044 10706 24050 10708
rect 24718 10706 24778 10918
rect 27520 10888 28000 10918
rect 24044 10646 24778 10706
rect 24044 10644 24050 10646
rect 0 10570 480 10600
rect 6361 10570 6427 10573
rect 0 10568 6427 10570
rect 0 10512 6366 10568
rect 6422 10512 6427 10568
rect 0 10510 6427 10512
rect 0 10480 480 10510
rect 6361 10507 6427 10510
rect 14365 10570 14431 10573
rect 19425 10570 19491 10573
rect 14365 10568 19491 10570
rect 14365 10512 14370 10568
rect 14426 10512 19430 10568
rect 19486 10512 19491 10568
rect 14365 10510 19491 10512
rect 14365 10507 14431 10510
rect 19425 10507 19491 10510
rect 19609 10570 19675 10573
rect 22921 10570 22987 10573
rect 25313 10570 25379 10573
rect 19609 10568 22800 10570
rect 19609 10512 19614 10568
rect 19670 10512 22800 10568
rect 19609 10510 22800 10512
rect 19609 10507 19675 10510
rect 4061 10434 4127 10437
rect 6177 10434 6243 10437
rect 4061 10432 6243 10434
rect 4061 10376 4066 10432
rect 4122 10376 6182 10432
rect 6238 10376 6243 10432
rect 4061 10374 6243 10376
rect 4061 10371 4127 10374
rect 6177 10371 6243 10374
rect 6453 10434 6519 10437
rect 10041 10434 10107 10437
rect 11145 10436 11211 10437
rect 11094 10434 11100 10436
rect 6453 10432 10107 10434
rect 6453 10376 6458 10432
rect 6514 10376 10046 10432
rect 10102 10376 10107 10432
rect 6453 10374 10107 10376
rect 11018 10374 11100 10434
rect 11164 10434 11211 10436
rect 11421 10434 11487 10437
rect 11164 10432 11487 10434
rect 11206 10376 11426 10432
rect 11482 10376 11487 10432
rect 6453 10371 6519 10374
rect 10041 10371 10107 10374
rect 11094 10372 11100 10374
rect 11164 10374 11487 10376
rect 22740 10434 22800 10510
rect 22921 10568 25379 10570
rect 22921 10512 22926 10568
rect 22982 10512 25318 10568
rect 25374 10512 25379 10568
rect 22921 10510 25379 10512
rect 22921 10507 22987 10510
rect 25313 10507 25379 10510
rect 27520 10434 28000 10464
rect 22740 10374 28000 10434
rect 11164 10372 11211 10374
rect 11145 10371 11211 10372
rect 11421 10371 11487 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 27520 10344 28000 10374
rect 19610 10303 19930 10304
rect 3785 10298 3851 10301
rect 4286 10298 4292 10300
rect 3785 10296 4292 10298
rect 3785 10240 3790 10296
rect 3846 10240 4292 10296
rect 3785 10238 4292 10240
rect 3785 10235 3851 10238
rect 4286 10236 4292 10238
rect 4356 10236 4362 10300
rect 6453 10298 6519 10301
rect 10041 10298 10107 10301
rect 6453 10296 10107 10298
rect 6453 10240 6458 10296
rect 6514 10240 10046 10296
rect 10102 10240 10107 10296
rect 6453 10238 10107 10240
rect 6453 10235 6519 10238
rect 10041 10235 10107 10238
rect 11145 10298 11211 10301
rect 13854 10298 13860 10300
rect 11145 10296 13860 10298
rect 11145 10240 11150 10296
rect 11206 10240 13860 10296
rect 11145 10238 13860 10240
rect 11145 10235 11211 10238
rect 13854 10236 13860 10238
rect 13924 10236 13930 10300
rect 14641 10298 14707 10301
rect 19328 10298 19334 10300
rect 14641 10296 19334 10298
rect 14641 10240 14646 10296
rect 14702 10240 19334 10296
rect 14641 10238 19334 10240
rect 14641 10235 14707 10238
rect 19328 10236 19334 10238
rect 19398 10236 19404 10300
rect 3141 10162 3207 10165
rect 11697 10162 11763 10165
rect 3141 10160 11763 10162
rect 3141 10104 3146 10160
rect 3202 10104 11702 10160
rect 11758 10104 11763 10160
rect 3141 10102 11763 10104
rect 3141 10099 3207 10102
rect 11697 10099 11763 10102
rect 12801 10162 12867 10165
rect 17401 10162 17467 10165
rect 12801 10160 17467 10162
rect 12801 10104 12806 10160
rect 12862 10104 17406 10160
rect 17462 10104 17467 10160
rect 12801 10102 17467 10104
rect 12801 10099 12867 10102
rect 17401 10099 17467 10102
rect 17769 10162 17835 10165
rect 21725 10162 21791 10165
rect 17769 10160 21791 10162
rect 17769 10104 17774 10160
rect 17830 10104 21730 10160
rect 21786 10104 21791 10160
rect 17769 10102 21791 10104
rect 17769 10099 17835 10102
rect 21725 10099 21791 10102
rect 24761 10162 24827 10165
rect 24761 10160 25882 10162
rect 24761 10104 24766 10160
rect 24822 10104 25882 10160
rect 24761 10102 25882 10104
rect 24761 10099 24827 10102
rect 0 10026 480 10056
rect 6126 10026 6132 10028
rect 0 9966 6132 10026
rect 0 9936 480 9966
rect 6126 9964 6132 9966
rect 6196 9964 6202 10028
rect 7373 10026 7439 10029
rect 12157 10026 12223 10029
rect 7373 10024 12223 10026
rect 7373 9968 7378 10024
rect 7434 9968 12162 10024
rect 12218 9968 12223 10024
rect 7373 9966 12223 9968
rect 7373 9963 7439 9966
rect 12157 9963 12223 9966
rect 14457 10026 14523 10029
rect 22185 10026 22251 10029
rect 25589 10026 25655 10029
rect 14457 10024 22251 10026
rect 14457 9968 14462 10024
rect 14518 9968 22190 10024
rect 22246 9968 22251 10024
rect 14457 9966 22251 9968
rect 14457 9963 14523 9966
rect 22185 9963 22251 9966
rect 24028 10024 25655 10026
rect 24028 9968 25594 10024
rect 25650 9968 25655 10024
rect 24028 9966 25655 9968
rect 3325 9890 3391 9893
rect 4613 9890 4679 9893
rect 3325 9888 4679 9890
rect 3325 9832 3330 9888
rect 3386 9832 4618 9888
rect 4674 9832 4679 9888
rect 3325 9830 4679 9832
rect 3325 9827 3391 9830
rect 4613 9827 4679 9830
rect 6361 9890 6427 9893
rect 14181 9890 14247 9893
rect 6361 9888 14247 9890
rect 6361 9832 6366 9888
rect 6422 9832 14186 9888
rect 14242 9832 14247 9888
rect 6361 9830 14247 9832
rect 6361 9827 6427 9830
rect 14181 9827 14247 9830
rect 15377 9890 15443 9893
rect 20437 9890 20503 9893
rect 24028 9890 24088 9966
rect 25589 9963 25655 9966
rect 15377 9888 24088 9890
rect 15377 9832 15382 9888
rect 15438 9832 20442 9888
rect 20498 9832 24088 9888
rect 15377 9830 24088 9832
rect 25822 9890 25882 10102
rect 27520 9890 28000 9920
rect 25822 9830 28000 9890
rect 15377 9827 15443 9830
rect 20437 9827 20503 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9830
rect 24277 9759 24597 9760
rect 10133 9754 10199 9757
rect 3052 9694 5504 9754
rect 3052 9618 3112 9694
rect 5444 9652 5504 9694
rect 5996 9752 10199 9754
rect 5996 9696 10138 9752
rect 10194 9696 10199 9752
rect 5996 9694 10199 9696
rect 3006 9558 3112 9618
rect 3325 9618 3391 9621
rect 3785 9618 3851 9621
rect 3325 9616 3851 9618
rect 3325 9560 3330 9616
rect 3386 9560 3790 9616
rect 3846 9560 3851 9616
rect 5444 9618 5596 9652
rect 5996 9618 6056 9694
rect 10133 9691 10199 9694
rect 12157 9754 12223 9757
rect 13813 9754 13879 9757
rect 12157 9752 13879 9754
rect 12157 9696 12162 9752
rect 12218 9696 13818 9752
rect 13874 9696 13879 9752
rect 12157 9694 13879 9696
rect 12157 9691 12223 9694
rect 13813 9691 13879 9694
rect 15837 9754 15903 9757
rect 22829 9754 22895 9757
rect 15837 9752 22895 9754
rect 15837 9696 15842 9752
rect 15898 9696 22834 9752
rect 22890 9696 22895 9752
rect 15837 9694 22895 9696
rect 15837 9691 15903 9694
rect 22829 9691 22895 9694
rect 5444 9592 6056 9618
rect 3325 9558 3851 9560
rect 5536 9558 6056 9592
rect 7281 9618 7347 9621
rect 8385 9618 8451 9621
rect 14457 9618 14523 9621
rect 18321 9618 18387 9621
rect 7281 9616 18387 9618
rect 7281 9560 7286 9616
rect 7342 9560 8390 9616
rect 8446 9560 14462 9616
rect 14518 9560 18326 9616
rect 18382 9560 18387 9616
rect 7281 9558 18387 9560
rect 0 9482 480 9512
rect 3006 9482 3066 9558
rect 3325 9555 3391 9558
rect 3785 9555 3851 9558
rect 7281 9555 7347 9558
rect 8385 9555 8451 9558
rect 14457 9555 14523 9558
rect 18321 9555 18387 9558
rect 18505 9618 18571 9621
rect 19977 9618 20043 9621
rect 18505 9616 20043 9618
rect 18505 9560 18510 9616
rect 18566 9560 19982 9616
rect 20038 9560 20043 9616
rect 18505 9558 20043 9560
rect 18505 9555 18571 9558
rect 19977 9555 20043 9558
rect 0 9422 3066 9482
rect 3141 9482 3207 9485
rect 3601 9482 3667 9485
rect 3141 9480 3667 9482
rect 3141 9424 3146 9480
rect 3202 9424 3606 9480
rect 3662 9424 3667 9480
rect 3141 9422 3667 9424
rect 0 9392 480 9422
rect 3141 9419 3207 9422
rect 3601 9419 3667 9422
rect 3785 9482 3851 9485
rect 12157 9482 12223 9485
rect 3785 9480 12223 9482
rect 3785 9424 3790 9480
rect 3846 9424 12162 9480
rect 12218 9424 12223 9480
rect 3785 9422 12223 9424
rect 3785 9419 3851 9422
rect 12157 9419 12223 9422
rect 12617 9482 12683 9485
rect 21909 9482 21975 9485
rect 23841 9482 23907 9485
rect 12617 9480 20178 9482
rect 12617 9424 12622 9480
rect 12678 9424 20178 9480
rect 12617 9422 20178 9424
rect 12617 9419 12683 9422
rect 2865 9346 2931 9349
rect 9305 9346 9371 9349
rect 2865 9344 9371 9346
rect 2865 9288 2870 9344
rect 2926 9288 9310 9344
rect 9366 9288 9371 9344
rect 2865 9286 9371 9288
rect 2865 9283 2931 9286
rect 9305 9283 9371 9286
rect 13077 9346 13143 9349
rect 13302 9346 13308 9348
rect 13077 9344 13308 9346
rect 13077 9288 13082 9344
rect 13138 9288 13308 9344
rect 13077 9286 13308 9288
rect 13077 9283 13143 9286
rect 13302 9284 13308 9286
rect 13372 9284 13378 9348
rect 14222 9284 14228 9348
rect 14292 9346 14298 9348
rect 14549 9346 14615 9349
rect 14292 9344 14615 9346
rect 14292 9288 14554 9344
rect 14610 9288 14615 9344
rect 14292 9286 14615 9288
rect 14292 9284 14298 9286
rect 14549 9283 14615 9286
rect 14825 9346 14891 9349
rect 18505 9346 18571 9349
rect 14825 9344 18571 9346
rect 14825 9288 14830 9344
rect 14886 9288 18510 9344
rect 18566 9288 18571 9344
rect 14825 9286 18571 9288
rect 20118 9346 20178 9422
rect 21909 9480 23907 9482
rect 21909 9424 21914 9480
rect 21970 9424 23846 9480
rect 23902 9424 23907 9480
rect 21909 9422 23907 9424
rect 21909 9419 21975 9422
rect 23841 9419 23907 9422
rect 22185 9346 22251 9349
rect 20118 9344 22251 9346
rect 20118 9288 22190 9344
rect 22246 9288 22251 9344
rect 20118 9286 22251 9288
rect 14825 9283 14891 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 17726 9213 17786 9286
rect 18505 9283 18571 9286
rect 22185 9283 22251 9286
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3601 9210 3667 9213
rect 3734 9210 3740 9212
rect 3601 9208 3740 9210
rect 3601 9152 3606 9208
rect 3662 9152 3740 9208
rect 3601 9150 3740 9152
rect 3601 9147 3667 9150
rect 3734 9148 3740 9150
rect 3804 9148 3810 9212
rect 13721 9210 13787 9213
rect 15653 9210 15719 9213
rect 13721 9208 15719 9210
rect 13721 9152 13726 9208
rect 13782 9152 15658 9208
rect 15714 9152 15719 9208
rect 13721 9150 15719 9152
rect 17726 9208 17835 9213
rect 17726 9152 17774 9208
rect 17830 9152 17835 9208
rect 17726 9150 17835 9152
rect 13721 9147 13787 9150
rect 15653 9147 15719 9150
rect 17769 9147 17835 9150
rect 23473 9210 23539 9213
rect 27520 9210 28000 9240
rect 23473 9208 28000 9210
rect 23473 9152 23478 9208
rect 23534 9152 28000 9208
rect 23473 9150 28000 9152
rect 23473 9147 23539 9150
rect 27520 9120 28000 9150
rect 1393 9074 1459 9077
rect 4521 9074 4587 9077
rect 1393 9072 4587 9074
rect 1393 9016 1398 9072
rect 1454 9016 4526 9072
rect 4582 9016 4587 9072
rect 1393 9014 4587 9016
rect 1393 9011 1459 9014
rect 4521 9011 4587 9014
rect 9673 9074 9739 9077
rect 20345 9074 20411 9077
rect 9673 9072 20411 9074
rect 9673 9016 9678 9072
rect 9734 9016 20350 9072
rect 20406 9016 20411 9072
rect 9673 9014 20411 9016
rect 9673 9011 9739 9014
rect 20345 9011 20411 9014
rect 23054 9012 23060 9076
rect 23124 9074 23130 9076
rect 24761 9074 24827 9077
rect 23124 9072 24827 9074
rect 23124 9016 24766 9072
rect 24822 9016 24827 9072
rect 23124 9014 24827 9016
rect 23124 9012 23130 9014
rect 24761 9011 24827 9014
rect 0 8938 480 8968
rect 8753 8938 8819 8941
rect 0 8936 8819 8938
rect 0 8880 8758 8936
rect 8814 8880 8819 8936
rect 0 8878 8819 8880
rect 0 8848 480 8878
rect 8753 8875 8819 8878
rect 9806 8876 9812 8940
rect 9876 8938 9882 8940
rect 21265 8938 21331 8941
rect 9876 8936 21331 8938
rect 9876 8880 21270 8936
rect 21326 8880 21331 8936
rect 9876 8878 21331 8880
rect 9876 8876 9882 8878
rect 21265 8875 21331 8878
rect 23974 8876 23980 8940
rect 24044 8938 24050 8940
rect 24044 8878 24778 8938
rect 24044 8876 24050 8878
rect 7966 8802 7972 8804
rect 6134 8742 7972 8802
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 4889 8530 4955 8533
rect 6134 8530 6194 8742
rect 7966 8740 7972 8742
rect 8036 8802 8042 8804
rect 8036 8742 10794 8802
rect 8036 8740 8042 8742
rect 7465 8666 7531 8669
rect 9857 8666 9923 8669
rect 7465 8664 9923 8666
rect 7465 8608 7470 8664
rect 7526 8608 9862 8664
rect 9918 8608 9923 8664
rect 7465 8606 9923 8608
rect 10734 8666 10794 8742
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 19885 8666 19951 8669
rect 21541 8666 21607 8669
rect 22093 8666 22159 8669
rect 10734 8606 12634 8666
rect 7465 8603 7531 8606
rect 9857 8603 9923 8606
rect 4889 8528 6194 8530
rect 4889 8472 4894 8528
rect 4950 8472 6194 8528
rect 4889 8470 6194 8472
rect 8293 8530 8359 8533
rect 10961 8530 11027 8533
rect 8293 8528 11027 8530
rect 8293 8472 8298 8528
rect 8354 8472 10966 8528
rect 11022 8472 11027 8528
rect 8293 8470 11027 8472
rect 12574 8530 12634 8606
rect 19885 8664 22159 8666
rect 19885 8608 19890 8664
rect 19946 8608 21546 8664
rect 21602 8608 22098 8664
rect 22154 8608 22159 8664
rect 19885 8606 22159 8608
rect 24718 8666 24778 8878
rect 27520 8666 28000 8696
rect 24718 8606 28000 8666
rect 19885 8603 19951 8606
rect 21541 8603 21607 8606
rect 22093 8603 22159 8606
rect 27520 8576 28000 8606
rect 16665 8530 16731 8533
rect 23657 8530 23723 8533
rect 12574 8528 23723 8530
rect 12574 8472 16670 8528
rect 16726 8472 23662 8528
rect 23718 8472 23723 8528
rect 12574 8470 23723 8472
rect 4889 8467 4955 8470
rect 8293 8467 8359 8470
rect 10961 8467 11027 8470
rect 16665 8467 16731 8470
rect 23657 8467 23723 8470
rect 6361 8394 6427 8397
rect 9765 8394 9831 8397
rect 6361 8392 9831 8394
rect 6361 8336 6366 8392
rect 6422 8336 9770 8392
rect 9826 8336 9831 8392
rect 6361 8334 9831 8336
rect 6361 8331 6427 8334
rect 9765 8331 9831 8334
rect 11237 8394 11303 8397
rect 15285 8394 15351 8397
rect 11237 8392 15351 8394
rect 11237 8336 11242 8392
rect 11298 8336 15290 8392
rect 15346 8336 15351 8392
rect 11237 8334 15351 8336
rect 11237 8331 11303 8334
rect 15285 8331 15351 8334
rect 0 8258 480 8288
rect 3785 8258 3851 8261
rect 4797 8260 4863 8261
rect 4797 8258 4844 8260
rect 0 8256 3851 8258
rect 0 8200 3790 8256
rect 3846 8200 3851 8256
rect 0 8198 3851 8200
rect 4752 8256 4844 8258
rect 4752 8200 4802 8256
rect 4752 8198 4844 8200
rect 0 8168 480 8198
rect 3785 8195 3851 8198
rect 4797 8196 4844 8198
rect 4908 8196 4914 8260
rect 8477 8258 8543 8261
rect 10133 8258 10199 8261
rect 8477 8256 10199 8258
rect 8477 8200 8482 8256
rect 8538 8200 10138 8256
rect 10194 8200 10199 8256
rect 8477 8198 10199 8200
rect 4797 8195 4863 8196
rect 8477 8195 8543 8198
rect 10133 8195 10199 8198
rect 10685 8258 10751 8261
rect 12801 8258 12867 8261
rect 10685 8256 12867 8258
rect 10685 8200 10690 8256
rect 10746 8200 12806 8256
rect 12862 8200 12867 8256
rect 10685 8198 12867 8200
rect 10685 8195 10751 8198
rect 12801 8195 12867 8198
rect 17401 8258 17467 8261
rect 19333 8258 19399 8261
rect 17401 8256 19399 8258
rect 17401 8200 17406 8256
rect 17462 8200 19338 8256
rect 19394 8200 19399 8256
rect 17401 8198 19399 8200
rect 17401 8195 17467 8198
rect 19333 8195 19399 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 5625 8122 5691 8125
rect 9857 8122 9923 8125
rect 18229 8122 18295 8125
rect 27520 8122 28000 8152
rect 5625 8120 9923 8122
rect 5625 8064 5630 8120
rect 5686 8064 9862 8120
rect 9918 8064 9923 8120
rect 5625 8062 9923 8064
rect 5625 8059 5691 8062
rect 9857 8059 9923 8062
rect 13494 8120 18295 8122
rect 13494 8064 18234 8120
rect 18290 8064 18295 8120
rect 13494 8062 18295 8064
rect 3509 7986 3575 7989
rect 13494 7986 13554 8062
rect 18229 8059 18295 8062
rect 24902 8062 28000 8122
rect 3509 7984 13554 7986
rect 3509 7928 3514 7984
rect 3570 7928 13554 7984
rect 3509 7926 13554 7928
rect 13629 7986 13695 7989
rect 24902 7986 24962 8062
rect 27520 8032 28000 8062
rect 13629 7984 24962 7986
rect 13629 7928 13634 7984
rect 13690 7928 24962 7984
rect 13629 7926 24962 7928
rect 3509 7923 3575 7926
rect 13629 7923 13695 7926
rect 2405 7850 2471 7853
rect 2630 7850 2636 7852
rect 2405 7848 2636 7850
rect 2405 7792 2410 7848
rect 2466 7792 2636 7848
rect 2405 7790 2636 7792
rect 2405 7787 2471 7790
rect 2630 7788 2636 7790
rect 2700 7788 2706 7852
rect 12157 7850 12223 7853
rect 5398 7848 12223 7850
rect 5398 7792 12162 7848
rect 12218 7792 12223 7848
rect 5398 7790 12223 7792
rect 0 7714 480 7744
rect 5398 7714 5458 7790
rect 12157 7787 12223 7790
rect 13077 7850 13143 7853
rect 19425 7850 19491 7853
rect 20345 7852 20411 7853
rect 13077 7848 19491 7850
rect 13077 7792 13082 7848
rect 13138 7792 19430 7848
rect 19486 7792 19491 7848
rect 13077 7790 19491 7792
rect 13077 7787 13143 7790
rect 19425 7787 19491 7790
rect 20294 7788 20300 7852
rect 20364 7850 20411 7852
rect 20897 7850 20963 7853
rect 25957 7850 26023 7853
rect 20364 7848 20456 7850
rect 20406 7792 20456 7848
rect 20364 7790 20456 7792
rect 20532 7848 26023 7850
rect 20532 7792 20902 7848
rect 20958 7792 25962 7848
rect 26018 7792 26023 7848
rect 20532 7790 26023 7792
rect 20364 7788 20411 7790
rect 20345 7787 20411 7788
rect 0 7654 5458 7714
rect 5993 7714 6059 7717
rect 10133 7714 10199 7717
rect 5993 7712 10199 7714
rect 5993 7656 5998 7712
rect 6054 7656 10138 7712
rect 10194 7656 10199 7712
rect 5993 7654 10199 7656
rect 0 7624 480 7654
rect 5993 7651 6059 7654
rect 10133 7651 10199 7654
rect 10317 7714 10383 7717
rect 10910 7714 10916 7716
rect 10317 7712 10916 7714
rect 10317 7656 10322 7712
rect 10378 7656 10916 7712
rect 10317 7654 10916 7656
rect 10317 7651 10383 7654
rect 10910 7652 10916 7654
rect 10980 7652 10986 7716
rect 12801 7714 12867 7717
rect 14733 7714 14799 7717
rect 12801 7712 14799 7714
rect 12801 7656 12806 7712
rect 12862 7656 14738 7712
rect 14794 7656 14799 7712
rect 12801 7654 14799 7656
rect 12801 7651 12867 7654
rect 14733 7651 14799 7654
rect 16297 7714 16363 7717
rect 18689 7714 18755 7717
rect 20532 7714 20592 7790
rect 20897 7787 20963 7790
rect 25957 7787 26023 7790
rect 16297 7712 20592 7714
rect 16297 7656 16302 7712
rect 16358 7656 18694 7712
rect 18750 7656 20592 7712
rect 16297 7654 20592 7656
rect 16297 7651 16363 7654
rect 18689 7651 18755 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 1485 7578 1551 7581
rect 3969 7578 4035 7581
rect 1485 7576 4035 7578
rect 1485 7520 1490 7576
rect 1546 7520 3974 7576
rect 4030 7520 4035 7576
rect 1485 7518 4035 7520
rect 1485 7515 1551 7518
rect 3969 7515 4035 7518
rect 10041 7578 10107 7581
rect 14457 7578 14523 7581
rect 16062 7578 16068 7580
rect 10041 7576 14523 7578
rect 10041 7520 10046 7576
rect 10102 7520 14462 7576
rect 14518 7520 14523 7576
rect 10041 7518 14523 7520
rect 10041 7515 10107 7518
rect 14457 7515 14523 7518
rect 15702 7518 16068 7578
rect 3972 7442 4032 7515
rect 12157 7442 12223 7445
rect 15702 7442 15762 7518
rect 16062 7516 16068 7518
rect 16132 7516 16138 7580
rect 17217 7578 17283 7581
rect 18781 7578 18847 7581
rect 20069 7578 20135 7581
rect 27520 7578 28000 7608
rect 17217 7576 20135 7578
rect 17217 7520 17222 7576
rect 17278 7520 18786 7576
rect 18842 7520 20074 7576
rect 20130 7520 20135 7576
rect 17217 7518 20135 7520
rect 17217 7515 17283 7518
rect 18781 7515 18847 7518
rect 20069 7515 20135 7518
rect 24902 7518 28000 7578
rect 3972 7382 10932 7442
rect 10685 7306 10751 7309
rect 1396 7304 10751 7306
rect 1396 7248 10690 7304
rect 10746 7248 10751 7304
rect 1396 7246 10751 7248
rect 0 7170 480 7200
rect 1396 7170 1456 7246
rect 10685 7243 10751 7246
rect 0 7110 1456 7170
rect 6085 7170 6151 7173
rect 6678 7170 6684 7172
rect 6085 7168 6684 7170
rect 6085 7112 6090 7168
rect 6146 7112 6684 7168
rect 6085 7110 6684 7112
rect 0 7080 480 7110
rect 6085 7107 6151 7110
rect 6678 7108 6684 7110
rect 6748 7108 6754 7172
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 10872 7034 10932 7382
rect 12157 7440 15762 7442
rect 12157 7384 12162 7440
rect 12218 7384 15762 7440
rect 12157 7382 15762 7384
rect 15837 7442 15903 7445
rect 19517 7442 19583 7445
rect 15837 7440 19583 7442
rect 15837 7384 15842 7440
rect 15898 7384 19522 7440
rect 19578 7384 19583 7440
rect 15837 7382 19583 7384
rect 12157 7379 12223 7382
rect 15837 7379 15903 7382
rect 19517 7379 19583 7382
rect 12433 7306 12499 7309
rect 15469 7306 15535 7309
rect 24902 7306 24962 7518
rect 27520 7488 28000 7518
rect 12433 7304 15535 7306
rect 12433 7248 12438 7304
rect 12494 7248 15474 7304
rect 15530 7248 15535 7304
rect 12433 7246 15535 7248
rect 12433 7243 12499 7246
rect 15469 7243 15535 7246
rect 17174 7246 24962 7306
rect 13629 7170 13695 7173
rect 15561 7170 15627 7173
rect 13629 7168 15627 7170
rect 13629 7112 13634 7168
rect 13690 7112 15566 7168
rect 15622 7112 15627 7168
rect 13629 7110 15627 7112
rect 13629 7107 13695 7110
rect 15561 7107 15627 7110
rect 11973 7034 12039 7037
rect 17174 7034 17234 7246
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 10872 7032 17234 7034
rect 10872 6976 11978 7032
rect 12034 6976 17234 7032
rect 10872 6974 17234 6976
rect 20069 7034 20135 7037
rect 27520 7034 28000 7064
rect 20069 7032 28000 7034
rect 20069 6976 20074 7032
rect 20130 6976 28000 7032
rect 20069 6974 28000 6976
rect 11973 6971 12039 6974
rect 20069 6971 20135 6974
rect 27520 6944 28000 6974
rect 4061 6898 4127 6901
rect 13997 6898 14063 6901
rect 4061 6896 14063 6898
rect 4061 6840 4066 6896
rect 4122 6840 14002 6896
rect 14058 6840 14063 6896
rect 4061 6838 14063 6840
rect 4061 6835 4127 6838
rect 13997 6835 14063 6838
rect 19241 6898 19307 6901
rect 20897 6898 20963 6901
rect 19241 6896 20963 6898
rect 19241 6840 19246 6896
rect 19302 6840 20902 6896
rect 20958 6840 20963 6896
rect 19241 6838 20963 6840
rect 19241 6835 19307 6838
rect 20897 6835 20963 6838
rect 21725 6898 21791 6901
rect 25129 6898 25195 6901
rect 21725 6896 25195 6898
rect 21725 6840 21730 6896
rect 21786 6840 25134 6896
rect 25190 6840 25195 6896
rect 21725 6838 25195 6840
rect 21725 6835 21791 6838
rect 25129 6835 25195 6838
rect 6269 6764 6335 6765
rect 6269 6762 6316 6764
rect 6188 6760 6316 6762
rect 6380 6762 6386 6764
rect 7097 6762 7163 6765
rect 9581 6762 9647 6765
rect 12157 6762 12223 6765
rect 21357 6762 21423 6765
rect 6380 6760 8034 6762
rect 6188 6704 6274 6760
rect 6380 6704 7102 6760
rect 7158 6704 8034 6760
rect 6188 6702 6316 6704
rect 6269 6700 6316 6702
rect 6380 6702 8034 6704
rect 6380 6700 6386 6702
rect 6269 6699 6335 6700
rect 7097 6699 7163 6702
rect 0 6626 480 6656
rect 2129 6626 2195 6629
rect 4981 6626 5047 6629
rect 0 6566 1456 6626
rect 0 6536 480 6566
rect 1396 6490 1456 6566
rect 2129 6624 5047 6626
rect 2129 6568 2134 6624
rect 2190 6568 4986 6624
rect 5042 6568 5047 6624
rect 2129 6566 5047 6568
rect 7974 6626 8034 6702
rect 9581 6760 12223 6762
rect 9581 6704 9586 6760
rect 9642 6704 12162 6760
rect 12218 6704 12223 6760
rect 9581 6702 12223 6704
rect 9581 6699 9647 6702
rect 12157 6699 12223 6702
rect 14414 6760 21423 6762
rect 14414 6704 21362 6760
rect 21418 6704 21423 6760
rect 14414 6702 21423 6704
rect 13302 6626 13308 6628
rect 7974 6566 13308 6626
rect 2129 6563 2195 6566
rect 4981 6563 5047 6566
rect 13302 6564 13308 6566
rect 13372 6626 13378 6628
rect 13670 6626 13676 6628
rect 13372 6566 13676 6626
rect 13372 6564 13378 6566
rect 13670 6564 13676 6566
rect 13740 6564 13746 6628
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 3734 6490 3740 6492
rect 1396 6430 3740 6490
rect 3734 6428 3740 6430
rect 3804 6428 3810 6492
rect 8569 6490 8635 6493
rect 14414 6492 14474 6702
rect 21357 6699 21423 6702
rect 23749 6762 23815 6765
rect 25037 6762 25103 6765
rect 23749 6760 25103 6762
rect 23749 6704 23754 6760
rect 23810 6704 25042 6760
rect 25098 6704 25103 6760
rect 23749 6702 25103 6704
rect 23749 6699 23815 6702
rect 25037 6699 25103 6702
rect 21817 6626 21883 6629
rect 24025 6626 24091 6629
rect 21817 6624 24091 6626
rect 21817 6568 21822 6624
rect 21878 6568 24030 6624
rect 24086 6568 24091 6624
rect 21817 6566 24091 6568
rect 21817 6563 21883 6566
rect 24025 6563 24091 6566
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 8702 6490 8708 6492
rect 8569 6488 8708 6490
rect 8569 6432 8574 6488
rect 8630 6432 8708 6488
rect 8569 6430 8708 6432
rect 8569 6427 8635 6430
rect 8702 6428 8708 6430
rect 8772 6428 8778 6492
rect 14406 6490 14412 6492
rect 8894 6430 14412 6490
rect 5625 6354 5691 6357
rect 8894 6354 8954 6430
rect 14406 6428 14412 6430
rect 14476 6428 14482 6492
rect 16113 6490 16179 6493
rect 21817 6490 21883 6493
rect 16113 6488 21883 6490
rect 16113 6432 16118 6488
rect 16174 6432 21822 6488
rect 21878 6432 21883 6488
rect 16113 6430 21883 6432
rect 16113 6427 16179 6430
rect 21817 6427 21883 6430
rect 22001 6490 22067 6493
rect 24117 6490 24183 6493
rect 27520 6490 28000 6520
rect 22001 6488 24183 6490
rect 22001 6432 22006 6488
rect 22062 6432 24122 6488
rect 24178 6432 24183 6488
rect 22001 6430 24183 6432
rect 22001 6427 22067 6430
rect 24117 6427 24183 6430
rect 24718 6430 28000 6490
rect 5625 6352 8954 6354
rect 5625 6296 5630 6352
rect 5686 6296 8954 6352
rect 5625 6294 8954 6296
rect 9397 6354 9463 6357
rect 11053 6354 11119 6357
rect 9397 6352 11119 6354
rect 9397 6296 9402 6352
rect 9458 6296 11058 6352
rect 11114 6296 11119 6352
rect 9397 6294 11119 6296
rect 5625 6291 5691 6294
rect 9397 6291 9463 6294
rect 11053 6291 11119 6294
rect 11329 6354 11395 6357
rect 22185 6354 22251 6357
rect 11329 6352 22251 6354
rect 11329 6296 11334 6352
rect 11390 6296 22190 6352
rect 22246 6296 22251 6352
rect 11329 6294 22251 6296
rect 11329 6291 11395 6294
rect 22185 6291 22251 6294
rect 22553 6354 22619 6357
rect 23749 6354 23815 6357
rect 22553 6352 23815 6354
rect 22553 6296 22558 6352
rect 22614 6296 23754 6352
rect 23810 6296 23815 6352
rect 22553 6294 23815 6296
rect 22553 6291 22619 6294
rect 23749 6291 23815 6294
rect 23974 6292 23980 6356
rect 24044 6354 24050 6356
rect 24718 6354 24778 6430
rect 27520 6400 28000 6430
rect 24044 6294 24778 6354
rect 24044 6292 24050 6294
rect 5073 6218 5139 6221
rect 8201 6218 8267 6221
rect 5073 6216 8267 6218
rect 5073 6160 5078 6216
rect 5134 6160 8206 6216
rect 8262 6160 8267 6216
rect 5073 6158 8267 6160
rect 5073 6155 5139 6158
rect 8201 6155 8267 6158
rect 8661 6218 8727 6221
rect 13445 6218 13511 6221
rect 8661 6216 13511 6218
rect 8661 6160 8666 6216
rect 8722 6160 13450 6216
rect 13506 6160 13511 6216
rect 8661 6158 13511 6160
rect 8661 6155 8727 6158
rect 13445 6155 13511 6158
rect 14590 6156 14596 6220
rect 14660 6218 14666 6220
rect 21541 6218 21607 6221
rect 14660 6216 21607 6218
rect 14660 6160 21546 6216
rect 21602 6160 21607 6216
rect 14660 6158 21607 6160
rect 14660 6156 14666 6158
rect 21541 6155 21607 6158
rect 21817 6218 21883 6221
rect 25405 6218 25471 6221
rect 21817 6216 25471 6218
rect 21817 6160 21822 6216
rect 21878 6160 25410 6216
rect 25466 6160 25471 6216
rect 21817 6158 25471 6160
rect 21817 6155 21883 6158
rect 25405 6155 25471 6158
rect 0 6082 480 6112
rect 3233 6082 3299 6085
rect 0 6080 3299 6082
rect 0 6024 3238 6080
rect 3294 6024 3299 6080
rect 0 6022 3299 6024
rect 0 5992 480 6022
rect 3233 6019 3299 6022
rect 3417 6082 3483 6085
rect 7373 6082 7439 6085
rect 3417 6080 7439 6082
rect 3417 6024 3422 6080
rect 3478 6024 7378 6080
rect 7434 6024 7439 6080
rect 3417 6022 7439 6024
rect 3417 6019 3483 6022
rect 7373 6019 7439 6022
rect 14549 6082 14615 6085
rect 18045 6082 18111 6085
rect 14549 6080 18111 6082
rect 14549 6024 14554 6080
rect 14610 6024 18050 6080
rect 18106 6024 18111 6080
rect 14549 6022 18111 6024
rect 14549 6019 14615 6022
rect 18045 6019 18111 6022
rect 21633 6082 21699 6085
rect 23657 6082 23723 6085
rect 25313 6082 25379 6085
rect 25957 6082 26023 6085
rect 21633 6080 23723 6082
rect 21633 6024 21638 6080
rect 21694 6024 23662 6080
rect 23718 6024 23723 6080
rect 21633 6022 23723 6024
rect 21633 6019 21699 6022
rect 23657 6019 23723 6022
rect 23798 6080 26023 6082
rect 23798 6024 25318 6080
rect 25374 6024 25962 6080
rect 26018 6024 26023 6080
rect 23798 6022 26023 6024
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 3325 5946 3391 5949
rect 6821 5946 6887 5949
rect 3325 5944 6887 5946
rect 3325 5888 3330 5944
rect 3386 5888 6826 5944
rect 6882 5888 6887 5944
rect 3325 5886 6887 5888
rect 3325 5883 3391 5886
rect 6821 5883 6887 5886
rect 7097 5946 7163 5949
rect 9397 5946 9463 5949
rect 7097 5944 9463 5946
rect 7097 5888 7102 5944
rect 7158 5888 9402 5944
rect 9458 5888 9463 5944
rect 7097 5886 9463 5888
rect 7097 5883 7163 5886
rect 9397 5883 9463 5886
rect 11421 5946 11487 5949
rect 18689 5946 18755 5949
rect 11421 5944 18755 5946
rect 11421 5888 11426 5944
rect 11482 5888 18694 5944
rect 18750 5888 18755 5944
rect 11421 5886 18755 5888
rect 11421 5883 11487 5886
rect 18689 5883 18755 5886
rect 20161 5946 20227 5949
rect 23798 5946 23858 6022
rect 25313 6019 25379 6022
rect 25957 6019 26023 6022
rect 20161 5944 23858 5946
rect 20161 5888 20166 5944
rect 20222 5888 23858 5944
rect 20161 5886 23858 5888
rect 20161 5883 20227 5886
rect 23974 5884 23980 5948
rect 24044 5946 24050 5948
rect 27520 5946 28000 5976
rect 24044 5886 28000 5946
rect 24044 5884 24050 5886
rect 27520 5856 28000 5886
rect 3601 5810 3667 5813
rect 12157 5810 12223 5813
rect 16481 5810 16547 5813
rect 19333 5810 19399 5813
rect 3601 5808 16314 5810
rect 3601 5752 3606 5808
rect 3662 5752 12162 5808
rect 12218 5752 16314 5808
rect 3601 5750 16314 5752
rect 3601 5747 3667 5750
rect 12157 5747 12223 5750
rect 5441 5674 5507 5677
rect 9806 5674 9812 5676
rect 5441 5672 9812 5674
rect 5441 5616 5446 5672
rect 5502 5616 9812 5672
rect 5441 5614 9812 5616
rect 5441 5611 5507 5614
rect 9806 5612 9812 5614
rect 9876 5612 9882 5676
rect 9949 5674 10015 5677
rect 13905 5674 13971 5677
rect 14641 5674 14707 5677
rect 9949 5672 14707 5674
rect 9949 5616 9954 5672
rect 10010 5616 13910 5672
rect 13966 5616 14646 5672
rect 14702 5616 14707 5672
rect 9949 5614 14707 5616
rect 16254 5674 16314 5750
rect 16481 5808 19399 5810
rect 16481 5752 16486 5808
rect 16542 5752 19338 5808
rect 19394 5752 19399 5808
rect 16481 5750 19399 5752
rect 16481 5747 16547 5750
rect 19333 5747 19399 5750
rect 19517 5810 19583 5813
rect 22553 5810 22619 5813
rect 19517 5808 22619 5810
rect 19517 5752 19522 5808
rect 19578 5752 22558 5808
rect 22614 5752 22619 5808
rect 19517 5750 22619 5752
rect 19517 5747 19583 5750
rect 22553 5747 22619 5750
rect 17217 5674 17283 5677
rect 17585 5674 17651 5677
rect 16254 5672 17651 5674
rect 16254 5616 17222 5672
rect 17278 5616 17590 5672
rect 17646 5616 17651 5672
rect 16254 5614 17651 5616
rect 9949 5611 10015 5614
rect 13905 5611 13971 5614
rect 14641 5611 14707 5614
rect 17217 5611 17283 5614
rect 17585 5611 17651 5614
rect 17861 5674 17927 5677
rect 21265 5674 21331 5677
rect 17861 5672 21331 5674
rect 17861 5616 17866 5672
rect 17922 5616 21270 5672
rect 21326 5616 21331 5672
rect 17861 5614 21331 5616
rect 17861 5611 17927 5614
rect 21265 5611 21331 5614
rect 21541 5674 21607 5677
rect 25957 5674 26023 5677
rect 21541 5672 26023 5674
rect 21541 5616 21546 5672
rect 21602 5616 25962 5672
rect 26018 5616 26023 5672
rect 21541 5614 26023 5616
rect 21541 5611 21607 5614
rect 25957 5611 26023 5614
rect 18229 5538 18295 5541
rect 23473 5538 23539 5541
rect 18229 5536 23539 5538
rect 18229 5480 18234 5536
rect 18290 5480 23478 5536
rect 23534 5480 23539 5536
rect 18229 5478 23539 5480
rect 18229 5475 18295 5478
rect 23473 5475 23539 5478
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 3366 5402 3372 5404
rect 0 5342 3372 5402
rect 0 5312 480 5342
rect 3366 5340 3372 5342
rect 3436 5340 3442 5404
rect 7741 5402 7807 5405
rect 7741 5400 14842 5402
rect 7741 5344 7746 5400
rect 7802 5344 14842 5400
rect 7741 5342 14842 5344
rect 7741 5339 7807 5342
rect 2221 5266 2287 5269
rect 8293 5266 8359 5269
rect 2221 5264 8359 5266
rect 2221 5208 2226 5264
rect 2282 5208 8298 5264
rect 8354 5208 8359 5264
rect 2221 5206 8359 5208
rect 2221 5203 2287 5206
rect 8293 5203 8359 5206
rect 9949 5266 10015 5269
rect 10685 5266 10751 5269
rect 13261 5266 13327 5269
rect 9949 5264 13327 5266
rect 9949 5208 9954 5264
rect 10010 5208 10690 5264
rect 10746 5208 13266 5264
rect 13322 5208 13327 5264
rect 9949 5206 13327 5208
rect 14782 5266 14842 5342
rect 15510 5340 15516 5404
rect 15580 5402 15586 5404
rect 15837 5402 15903 5405
rect 15580 5400 15903 5402
rect 15580 5344 15842 5400
rect 15898 5344 15903 5400
rect 15580 5342 15903 5344
rect 15580 5340 15586 5342
rect 15837 5339 15903 5342
rect 16941 5402 17007 5405
rect 19425 5402 19491 5405
rect 16941 5400 19491 5402
rect 16941 5344 16946 5400
rect 17002 5344 19430 5400
rect 19486 5344 19491 5400
rect 16941 5342 19491 5344
rect 16941 5339 17007 5342
rect 19425 5339 19491 5342
rect 22553 5402 22619 5405
rect 23473 5402 23539 5405
rect 23606 5402 23612 5404
rect 22553 5400 23612 5402
rect 22553 5344 22558 5400
rect 22614 5344 23478 5400
rect 23534 5344 23612 5400
rect 22553 5342 23612 5344
rect 22553 5339 22619 5342
rect 23473 5339 23539 5342
rect 23606 5340 23612 5342
rect 23676 5340 23682 5404
rect 27520 5402 28000 5432
rect 24718 5342 28000 5402
rect 16941 5266 17007 5269
rect 18229 5266 18295 5269
rect 14782 5264 18295 5266
rect 14782 5208 16946 5264
rect 17002 5208 18234 5264
rect 18290 5208 18295 5264
rect 14782 5206 18295 5208
rect 9949 5203 10015 5206
rect 10685 5203 10751 5206
rect 13261 5203 13327 5206
rect 16941 5203 17007 5206
rect 18229 5203 18295 5206
rect 23933 5266 23999 5269
rect 24718 5266 24778 5342
rect 27520 5312 28000 5342
rect 23933 5264 24778 5266
rect 23933 5208 23938 5264
rect 23994 5208 24778 5264
rect 23933 5206 24778 5208
rect 23933 5203 23999 5206
rect 6269 5130 6335 5133
rect 17769 5130 17835 5133
rect 19701 5130 19767 5133
rect 24577 5130 24643 5133
rect 6269 5128 17835 5130
rect 6269 5072 6274 5128
rect 6330 5072 17774 5128
rect 17830 5072 17835 5128
rect 6269 5070 17835 5072
rect 6269 5067 6335 5070
rect 17769 5067 17835 5070
rect 17910 5128 24643 5130
rect 17910 5072 19706 5128
rect 19762 5072 24582 5128
rect 24638 5072 24643 5128
rect 17910 5070 24643 5072
rect 2129 4994 2195 4997
rect 9949 4994 10015 4997
rect 2129 4992 10015 4994
rect 2129 4936 2134 4992
rect 2190 4936 9954 4992
rect 10010 4936 10015 4992
rect 2129 4934 10015 4936
rect 2129 4931 2195 4934
rect 9949 4931 10015 4934
rect 11605 4994 11671 4997
rect 12433 4994 12499 4997
rect 17910 4994 17970 5070
rect 19701 5067 19767 5070
rect 24577 5067 24643 5070
rect 11605 4992 17970 4994
rect 11605 4936 11610 4992
rect 11666 4936 12438 4992
rect 12494 4936 17970 4992
rect 11605 4934 17970 4936
rect 21909 4994 21975 4997
rect 22553 4994 22619 4997
rect 21909 4992 22619 4994
rect 21909 4936 21914 4992
rect 21970 4936 22558 4992
rect 22614 4936 22619 4992
rect 21909 4934 22619 4936
rect 11605 4931 11671 4934
rect 12433 4931 12499 4934
rect 21909 4931 21975 4934
rect 22553 4931 22619 4934
rect 22737 4994 22803 4997
rect 23933 4994 23999 4997
rect 22737 4992 23999 4994
rect 22737 4936 22742 4992
rect 22798 4936 23938 4992
rect 23994 4936 23999 4992
rect 22737 4934 23999 4936
rect 22737 4931 22803 4934
rect 23933 4931 23999 4934
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 480 4798
rect 3969 4795 4035 4798
rect 6913 4858 6979 4861
rect 21909 4858 21975 4861
rect 6913 4856 10058 4858
rect 6913 4800 6918 4856
rect 6974 4800 10058 4856
rect 6913 4798 10058 4800
rect 6913 4795 6979 4798
rect 7649 4722 7715 4725
rect 9998 4722 10058 4798
rect 20164 4856 21975 4858
rect 20164 4800 21914 4856
rect 21970 4800 21975 4856
rect 20164 4798 21975 4800
rect 17493 4722 17559 4725
rect 20164 4722 20224 4798
rect 21909 4795 21975 4798
rect 7649 4720 9874 4722
rect 7649 4664 7654 4720
rect 7710 4664 9874 4720
rect 7649 4662 9874 4664
rect 9998 4662 17234 4722
rect 7649 4659 7715 4662
rect 2313 4586 2379 4589
rect 8109 4586 8175 4589
rect 2313 4584 8175 4586
rect 2313 4528 2318 4584
rect 2374 4528 8114 4584
rect 8170 4528 8175 4584
rect 2313 4526 8175 4528
rect 9814 4586 9874 4662
rect 11973 4586 12039 4589
rect 17033 4586 17099 4589
rect 9814 4584 17099 4586
rect 9814 4528 11978 4584
rect 12034 4528 17038 4584
rect 17094 4528 17099 4584
rect 9814 4526 17099 4528
rect 17174 4586 17234 4662
rect 17493 4720 20224 4722
rect 17493 4664 17498 4720
rect 17554 4664 20224 4720
rect 17493 4662 20224 4664
rect 23749 4722 23815 4725
rect 24669 4722 24735 4725
rect 27520 4722 28000 4752
rect 23749 4720 24735 4722
rect 23749 4664 23754 4720
rect 23810 4664 24674 4720
rect 24730 4664 24735 4720
rect 23749 4662 24735 4664
rect 17493 4659 17559 4662
rect 23749 4659 23815 4662
rect 24669 4659 24735 4662
rect 24902 4662 28000 4722
rect 24902 4586 24962 4662
rect 27520 4632 28000 4662
rect 17174 4526 24962 4586
rect 2313 4523 2379 4526
rect 8109 4523 8175 4526
rect 11973 4523 12039 4526
rect 17033 4523 17099 4526
rect 12801 4452 12867 4453
rect 12750 4388 12756 4452
rect 12820 4450 12867 4452
rect 13445 4450 13511 4453
rect 17217 4450 17283 4453
rect 23473 4452 23539 4453
rect 12820 4448 12912 4450
rect 12862 4392 12912 4448
rect 12820 4390 12912 4392
rect 13445 4448 14290 4450
rect 13445 4392 13450 4448
rect 13506 4392 14290 4448
rect 13445 4390 14290 4392
rect 12820 4388 12867 4390
rect 12801 4387 12867 4388
rect 13445 4387 13511 4390
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 480 4254
rect 1669 4251 1735 4254
rect 4981 4314 5047 4317
rect 5206 4314 5212 4316
rect 4981 4312 5212 4314
rect 4981 4256 4986 4312
rect 5042 4256 5212 4312
rect 4981 4254 5212 4256
rect 4981 4251 5047 4254
rect 5206 4252 5212 4254
rect 5276 4252 5282 4316
rect 11789 4314 11855 4317
rect 13445 4314 13511 4317
rect 11789 4312 13511 4314
rect 11789 4256 11794 4312
rect 11850 4256 13450 4312
rect 13506 4256 13511 4312
rect 11789 4254 13511 4256
rect 11789 4251 11855 4254
rect 13445 4251 13511 4254
rect 1853 4178 1919 4181
rect 4245 4178 4311 4181
rect 1853 4176 4311 4178
rect 1853 4120 1858 4176
rect 1914 4120 4250 4176
rect 4306 4120 4311 4176
rect 1853 4118 4311 4120
rect 1853 4115 1919 4118
rect 4245 4115 4311 4118
rect 11513 4178 11579 4181
rect 14089 4178 14155 4181
rect 11513 4176 14155 4178
rect 11513 4120 11518 4176
rect 11574 4120 14094 4176
rect 14150 4120 14155 4176
rect 11513 4118 14155 4120
rect 14230 4178 14290 4390
rect 17217 4448 23306 4450
rect 17217 4392 17222 4448
rect 17278 4392 23306 4448
rect 17217 4390 23306 4392
rect 17217 4387 17283 4390
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 23246 4314 23306 4390
rect 23422 4388 23428 4452
rect 23492 4450 23539 4452
rect 23492 4448 23584 4450
rect 23534 4392 23584 4448
rect 23492 4390 23584 4392
rect 23492 4388 23539 4390
rect 23473 4387 23539 4388
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 24117 4314 24183 4317
rect 15334 4254 23122 4314
rect 23246 4312 24183 4314
rect 23246 4256 24122 4312
rect 24178 4256 24183 4312
rect 23246 4254 24183 4256
rect 15334 4178 15394 4254
rect 14230 4118 15394 4178
rect 19149 4178 19215 4181
rect 22001 4178 22067 4181
rect 19149 4176 22067 4178
rect 19149 4120 19154 4176
rect 19210 4120 22006 4176
rect 22062 4120 22067 4176
rect 19149 4118 22067 4120
rect 23062 4178 23122 4254
rect 24117 4251 24183 4254
rect 24669 4314 24735 4317
rect 24669 4312 25146 4314
rect 24669 4256 24674 4312
rect 24730 4256 25146 4312
rect 24669 4254 25146 4256
rect 24669 4251 24735 4254
rect 24945 4178 25011 4181
rect 23062 4176 25011 4178
rect 23062 4120 24950 4176
rect 25006 4120 25011 4176
rect 23062 4118 25011 4120
rect 25086 4178 25146 4254
rect 27520 4178 28000 4208
rect 25086 4118 28000 4178
rect 11513 4115 11579 4118
rect 14089 4115 14155 4118
rect 19149 4115 19215 4118
rect 22001 4115 22067 4118
rect 24945 4115 25011 4118
rect 27520 4088 28000 4118
rect 2957 4042 3023 4045
rect 4797 4042 4863 4045
rect 6545 4042 6611 4045
rect 2957 4040 6611 4042
rect 2957 3984 2962 4040
rect 3018 3984 4802 4040
rect 4858 3984 6550 4040
rect 6606 3984 6611 4040
rect 2957 3982 6611 3984
rect 2957 3979 3023 3982
rect 4797 3979 4863 3982
rect 6545 3979 6611 3982
rect 8017 4042 8083 4045
rect 12157 4042 12223 4045
rect 13077 4042 13143 4045
rect 8017 4040 13143 4042
rect 8017 3984 8022 4040
rect 8078 3984 12162 4040
rect 12218 3984 13082 4040
rect 13138 3984 13143 4040
rect 8017 3982 13143 3984
rect 8017 3979 8083 3982
rect 12157 3979 12223 3982
rect 13077 3979 13143 3982
rect 15745 4042 15811 4045
rect 16481 4042 16547 4045
rect 15745 4040 16547 4042
rect 15745 3984 15750 4040
rect 15806 3984 16486 4040
rect 16542 3984 16547 4040
rect 15745 3982 16547 3984
rect 15745 3979 15811 3982
rect 16481 3979 16547 3982
rect 16614 3980 16620 4044
rect 16684 4042 16690 4044
rect 16757 4042 16823 4045
rect 16684 4040 16823 4042
rect 16684 3984 16762 4040
rect 16818 3984 16823 4040
rect 16684 3982 16823 3984
rect 16684 3980 16690 3982
rect 16757 3979 16823 3982
rect 17125 4042 17191 4045
rect 20805 4042 20871 4045
rect 17125 4040 20871 4042
rect 17125 3984 17130 4040
rect 17186 3984 20810 4040
rect 20866 3984 20871 4040
rect 17125 3982 20871 3984
rect 17125 3979 17191 3982
rect 20805 3979 20871 3982
rect 22829 4042 22895 4045
rect 24117 4042 24183 4045
rect 22829 4040 24183 4042
rect 22829 3984 22834 4040
rect 22890 3984 24122 4040
rect 24178 3984 24183 4040
rect 22829 3982 24183 3984
rect 22829 3979 22895 3982
rect 24117 3979 24183 3982
rect 8293 3908 8359 3909
rect 8293 3906 8340 3908
rect 8248 3904 8340 3906
rect 8248 3848 8298 3904
rect 8248 3846 8340 3848
rect 8293 3844 8340 3846
rect 8404 3844 8410 3908
rect 10685 3906 10751 3909
rect 13353 3906 13419 3909
rect 10685 3904 13419 3906
rect 10685 3848 10690 3904
rect 10746 3848 13358 3904
rect 13414 3848 13419 3904
rect 10685 3846 13419 3848
rect 8293 3843 8359 3844
rect 10685 3843 10751 3846
rect 13353 3843 13419 3846
rect 15837 3906 15903 3909
rect 19425 3906 19491 3909
rect 15837 3904 19491 3906
rect 15837 3848 15842 3904
rect 15898 3848 19430 3904
rect 19486 3848 19491 3904
rect 15837 3846 19491 3848
rect 15837 3843 15903 3846
rect 19425 3843 19491 3846
rect 22737 3906 22803 3909
rect 25129 3906 25195 3909
rect 22737 3904 25195 3906
rect 22737 3848 22742 3904
rect 22798 3848 25134 3904
rect 25190 3848 25195 3904
rect 22737 3846 25195 3848
rect 22737 3843 22803 3846
rect 25129 3843 25195 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1577 3770 1643 3773
rect 9857 3770 9923 3773
rect 0 3710 1456 3770
rect 0 3680 480 3710
rect 1396 3498 1456 3710
rect 1577 3768 9923 3770
rect 1577 3712 1582 3768
rect 1638 3712 9862 3768
rect 9918 3712 9923 3768
rect 1577 3710 9923 3712
rect 1577 3707 1643 3710
rect 9857 3707 9923 3710
rect 10777 3770 10843 3773
rect 14641 3770 14707 3773
rect 15837 3770 15903 3773
rect 10777 3768 15903 3770
rect 10777 3712 10782 3768
rect 10838 3712 14646 3768
rect 14702 3712 15842 3768
rect 15898 3712 15903 3768
rect 10777 3710 15903 3712
rect 10777 3707 10843 3710
rect 14641 3707 14707 3710
rect 15837 3707 15903 3710
rect 16062 3708 16068 3772
rect 16132 3770 16138 3772
rect 16297 3770 16363 3773
rect 16132 3768 16363 3770
rect 16132 3712 16302 3768
rect 16358 3712 16363 3768
rect 16132 3710 16363 3712
rect 16132 3708 16138 3710
rect 16297 3707 16363 3710
rect 16481 3770 16547 3773
rect 19425 3770 19491 3773
rect 22369 3770 22435 3773
rect 24577 3770 24643 3773
rect 16481 3768 19491 3770
rect 16481 3712 16486 3768
rect 16542 3712 19430 3768
rect 19486 3712 19491 3768
rect 16481 3710 19491 3712
rect 16481 3707 16547 3710
rect 19425 3707 19491 3710
rect 20118 3768 24643 3770
rect 20118 3712 22374 3768
rect 22430 3712 24582 3768
rect 24638 3712 24643 3768
rect 20118 3710 24643 3712
rect 2865 3634 2931 3637
rect 3141 3634 3207 3637
rect 8293 3634 8359 3637
rect 2865 3632 8359 3634
rect 2865 3576 2870 3632
rect 2926 3576 3146 3632
rect 3202 3576 8298 3632
rect 8354 3576 8359 3632
rect 2865 3574 8359 3576
rect 2865 3571 2931 3574
rect 3141 3571 3207 3574
rect 8293 3571 8359 3574
rect 14457 3634 14523 3637
rect 17217 3634 17283 3637
rect 14457 3632 17283 3634
rect 14457 3576 14462 3632
rect 14518 3576 17222 3632
rect 17278 3576 17283 3632
rect 14457 3574 17283 3576
rect 14457 3571 14523 3574
rect 17217 3571 17283 3574
rect 18873 3634 18939 3637
rect 20118 3634 20178 3710
rect 22369 3707 22435 3710
rect 24577 3707 24643 3710
rect 18873 3632 20178 3634
rect 18873 3576 18878 3632
rect 18934 3576 20178 3632
rect 18873 3574 20178 3576
rect 20253 3634 20319 3637
rect 23565 3634 23631 3637
rect 20253 3632 23631 3634
rect 20253 3576 20258 3632
rect 20314 3576 23570 3632
rect 23626 3576 23631 3632
rect 20253 3574 23631 3576
rect 18873 3571 18939 3574
rect 20253 3571 20319 3574
rect 23565 3571 23631 3574
rect 24301 3634 24367 3637
rect 27520 3634 28000 3664
rect 24301 3632 28000 3634
rect 24301 3576 24306 3632
rect 24362 3576 28000 3632
rect 24301 3574 28000 3576
rect 24301 3571 24367 3574
rect 27520 3544 28000 3574
rect 3417 3498 3483 3501
rect 3877 3498 3943 3501
rect 1396 3496 3943 3498
rect 1396 3440 3422 3496
rect 3478 3440 3882 3496
rect 3938 3440 3943 3496
rect 1396 3438 3943 3440
rect 3417 3435 3483 3438
rect 3877 3435 3943 3438
rect 12617 3498 12683 3501
rect 19517 3498 19583 3501
rect 12617 3496 19583 3498
rect 12617 3440 12622 3496
rect 12678 3440 19522 3496
rect 19578 3440 19583 3496
rect 12617 3438 19583 3440
rect 12617 3435 12683 3438
rect 19517 3435 19583 3438
rect 19701 3498 19767 3501
rect 23013 3498 23079 3501
rect 19701 3496 23079 3498
rect 19701 3440 19706 3496
rect 19762 3440 23018 3496
rect 23074 3440 23079 3496
rect 19701 3438 23079 3440
rect 19701 3435 19767 3438
rect 23013 3435 23079 3438
rect 17217 3362 17283 3365
rect 20253 3362 20319 3365
rect 17217 3360 20319 3362
rect 17217 3304 17222 3360
rect 17278 3304 20258 3360
rect 20314 3304 20319 3360
rect 17217 3302 20319 3304
rect 17217 3299 17283 3302
rect 20253 3299 20319 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 657 3226 723 3229
rect 0 3224 723 3226
rect 0 3168 662 3224
rect 718 3168 723 3224
rect 0 3166 723 3168
rect 0 3136 480 3166
rect 657 3163 723 3166
rect 841 3226 907 3229
rect 1158 3226 1164 3228
rect 841 3224 1164 3226
rect 841 3168 846 3224
rect 902 3168 1164 3224
rect 841 3166 1164 3168
rect 841 3163 907 3166
rect 1158 3164 1164 3166
rect 1228 3164 1234 3228
rect 9213 3226 9279 3229
rect 7790 3224 9279 3226
rect 7790 3168 9218 3224
rect 9274 3168 9279 3224
rect 7790 3166 9279 3168
rect 2589 3090 2655 3093
rect 7790 3090 7850 3166
rect 9213 3163 9279 3166
rect 15929 3226 15995 3229
rect 22093 3226 22159 3229
rect 15929 3224 22159 3226
rect 15929 3168 15934 3224
rect 15990 3168 22098 3224
rect 22154 3168 22159 3224
rect 15929 3166 22159 3168
rect 15929 3163 15995 3166
rect 22093 3163 22159 3166
rect 2589 3088 7850 3090
rect 2589 3032 2594 3088
rect 2650 3032 7850 3088
rect 2589 3030 7850 3032
rect 8017 3090 8083 3093
rect 14181 3090 14247 3093
rect 15837 3090 15903 3093
rect 16573 3092 16639 3093
rect 16573 3090 16620 3092
rect 8017 3088 14106 3090
rect 8017 3032 8022 3088
rect 8078 3032 14106 3088
rect 8017 3030 14106 3032
rect 2589 3027 2655 3030
rect 8017 3027 8083 3030
rect 4153 2954 4219 2957
rect 13629 2954 13695 2957
rect 4153 2952 13695 2954
rect 4153 2896 4158 2952
rect 4214 2896 13634 2952
rect 13690 2896 13695 2952
rect 4153 2894 13695 2896
rect 14046 2954 14106 3030
rect 14181 3088 15903 3090
rect 14181 3032 14186 3088
rect 14242 3032 15842 3088
rect 15898 3032 15903 3088
rect 14181 3030 15903 3032
rect 16528 3088 16620 3090
rect 16528 3032 16578 3088
rect 16528 3030 16620 3032
rect 14181 3027 14247 3030
rect 15837 3027 15903 3030
rect 16573 3028 16620 3030
rect 16684 3028 16690 3092
rect 19057 3090 19123 3093
rect 20713 3090 20779 3093
rect 19057 3088 20779 3090
rect 19057 3032 19062 3088
rect 19118 3032 20718 3088
rect 20774 3032 20779 3088
rect 19057 3030 20779 3032
rect 16573 3027 16639 3028
rect 19057 3027 19123 3030
rect 20713 3027 20779 3030
rect 25865 3090 25931 3093
rect 27520 3090 28000 3120
rect 25865 3088 28000 3090
rect 25865 3032 25870 3088
rect 25926 3032 28000 3088
rect 25865 3030 28000 3032
rect 25865 3027 25931 3030
rect 27520 3000 28000 3030
rect 14549 2954 14615 2957
rect 14825 2954 14891 2957
rect 14046 2952 14891 2954
rect 14046 2896 14554 2952
rect 14610 2896 14830 2952
rect 14886 2896 14891 2952
rect 14046 2894 14891 2896
rect 4153 2891 4219 2894
rect 13629 2891 13695 2894
rect 14549 2891 14615 2894
rect 14825 2891 14891 2894
rect 15101 2954 15167 2957
rect 17033 2954 17099 2957
rect 24025 2954 24091 2957
rect 15101 2952 17099 2954
rect 15101 2896 15106 2952
rect 15162 2896 17038 2952
rect 17094 2896 17099 2952
rect 15101 2894 17099 2896
rect 15101 2891 15167 2894
rect 17033 2891 17099 2894
rect 17174 2952 24091 2954
rect 17174 2896 24030 2952
rect 24086 2896 24091 2952
rect 17174 2894 24091 2896
rect 2497 2818 2563 2821
rect 6821 2818 6887 2821
rect 8569 2818 8635 2821
rect 2497 2816 8635 2818
rect 2497 2760 2502 2816
rect 2558 2760 6826 2816
rect 6882 2760 8574 2816
rect 8630 2760 8635 2816
rect 2497 2758 8635 2760
rect 2497 2755 2563 2758
rect 6821 2755 6887 2758
rect 8569 2755 8635 2758
rect 13721 2818 13787 2821
rect 17174 2818 17234 2894
rect 24025 2891 24091 2894
rect 13721 2816 17234 2818
rect 13721 2760 13726 2816
rect 13782 2760 17234 2816
rect 13721 2758 17234 2760
rect 13721 2755 13787 2758
rect 17350 2756 17356 2820
rect 17420 2818 17426 2820
rect 17493 2818 17559 2821
rect 17420 2816 17559 2818
rect 17420 2760 17498 2816
rect 17554 2760 17559 2816
rect 17420 2758 17559 2760
rect 17420 2756 17426 2758
rect 17493 2755 17559 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1393 2682 1459 2685
rect 4429 2682 4495 2685
rect 4889 2684 4955 2685
rect 4838 2682 4844 2684
rect 1393 2680 4495 2682
rect 1393 2624 1398 2680
rect 1454 2624 4434 2680
rect 4490 2624 4495 2680
rect 1393 2622 4495 2624
rect 4798 2622 4844 2682
rect 4908 2680 4955 2684
rect 4950 2624 4955 2680
rect 1393 2619 1459 2622
rect 4429 2619 4495 2622
rect 4838 2620 4844 2622
rect 4908 2620 4955 2624
rect 4889 2619 4955 2620
rect 6453 2682 6519 2685
rect 9121 2682 9187 2685
rect 6453 2680 9187 2682
rect 6453 2624 6458 2680
rect 6514 2624 9126 2680
rect 9182 2624 9187 2680
rect 6453 2622 9187 2624
rect 6453 2619 6519 2622
rect 9121 2619 9187 2622
rect 11237 2682 11303 2685
rect 14641 2682 14707 2685
rect 11237 2680 14707 2682
rect 11237 2624 11242 2680
rect 11298 2624 14646 2680
rect 14702 2624 14707 2680
rect 11237 2622 14707 2624
rect 11237 2619 11303 2622
rect 14641 2619 14707 2622
rect 15929 2682 15995 2685
rect 18045 2682 18111 2685
rect 15929 2680 18111 2682
rect 15929 2624 15934 2680
rect 15990 2624 18050 2680
rect 18106 2624 18111 2680
rect 15929 2622 18111 2624
rect 15929 2619 15995 2622
rect 18045 2619 18111 2622
rect 23197 2682 23263 2685
rect 25589 2682 25655 2685
rect 23197 2680 25655 2682
rect 23197 2624 23202 2680
rect 23258 2624 25594 2680
rect 25650 2624 25655 2680
rect 23197 2622 25655 2624
rect 23197 2619 23263 2622
rect 25589 2619 25655 2622
rect 0 2546 480 2576
rect 3417 2546 3483 2549
rect 0 2544 3483 2546
rect 0 2488 3422 2544
rect 3478 2488 3483 2544
rect 0 2486 3483 2488
rect 0 2456 480 2486
rect 3417 2483 3483 2486
rect 8201 2546 8267 2549
rect 16389 2546 16455 2549
rect 18045 2546 18111 2549
rect 8201 2544 15762 2546
rect 8201 2488 8206 2544
rect 8262 2488 15762 2544
rect 8201 2486 15762 2488
rect 8201 2483 8267 2486
rect 9806 2348 9812 2412
rect 9876 2410 9882 2412
rect 10317 2410 10383 2413
rect 9876 2408 10383 2410
rect 9876 2352 10322 2408
rect 10378 2352 10383 2408
rect 9876 2350 10383 2352
rect 9876 2348 9882 2350
rect 10317 2347 10383 2350
rect 10869 2410 10935 2413
rect 15469 2410 15535 2413
rect 10869 2408 15535 2410
rect 10869 2352 10874 2408
rect 10930 2352 15474 2408
rect 15530 2352 15535 2408
rect 10869 2350 15535 2352
rect 15702 2410 15762 2486
rect 16389 2544 18111 2546
rect 16389 2488 16394 2544
rect 16450 2488 18050 2544
rect 18106 2488 18111 2544
rect 16389 2486 18111 2488
rect 16389 2483 16455 2486
rect 18045 2483 18111 2486
rect 18321 2546 18387 2549
rect 20529 2546 20595 2549
rect 18321 2544 20595 2546
rect 18321 2488 18326 2544
rect 18382 2488 20534 2544
rect 20590 2488 20595 2544
rect 18321 2486 20595 2488
rect 18321 2483 18387 2486
rect 20529 2483 20595 2486
rect 21541 2546 21607 2549
rect 24025 2546 24091 2549
rect 21541 2544 24091 2546
rect 21541 2488 21546 2544
rect 21602 2488 24030 2544
rect 24086 2488 24091 2544
rect 21541 2486 24091 2488
rect 21541 2483 21607 2486
rect 24025 2483 24091 2486
rect 24761 2546 24827 2549
rect 27520 2546 28000 2576
rect 24761 2544 28000 2546
rect 24761 2488 24766 2544
rect 24822 2488 28000 2544
rect 24761 2486 28000 2488
rect 24761 2483 24827 2486
rect 27520 2456 28000 2486
rect 23473 2410 23539 2413
rect 15702 2408 23539 2410
rect 15702 2352 23478 2408
rect 23534 2352 23539 2408
rect 15702 2350 23539 2352
rect 10869 2347 10935 2350
rect 15469 2347 15535 2350
rect 23473 2347 23539 2350
rect 10777 2274 10843 2277
rect 14457 2274 14523 2277
rect 10777 2272 14523 2274
rect 10777 2216 10782 2272
rect 10838 2216 14462 2272
rect 14518 2216 14523 2272
rect 10777 2214 14523 2216
rect 10777 2211 10843 2214
rect 14457 2211 14523 2214
rect 21449 2274 21515 2277
rect 23473 2274 23539 2277
rect 21449 2272 23539 2274
rect 21449 2216 21454 2272
rect 21510 2216 23478 2272
rect 23534 2216 23539 2272
rect 21449 2214 23539 2216
rect 21449 2211 21515 2214
rect 23473 2211 23539 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 17677 2138 17743 2141
rect 22553 2138 22619 2141
rect 17677 2136 22619 2138
rect 17677 2080 17682 2136
rect 17738 2080 22558 2136
rect 22614 2080 22619 2136
rect 17677 2078 22619 2080
rect 17677 2075 17743 2078
rect 22553 2075 22619 2078
rect 0 2002 480 2032
rect 2405 2002 2471 2005
rect 0 2000 2471 2002
rect 0 1944 2410 2000
rect 2466 1944 2471 2000
rect 0 1942 2471 1944
rect 0 1912 480 1942
rect 2405 1939 2471 1942
rect 6177 2002 6243 2005
rect 18137 2002 18203 2005
rect 6177 2000 18203 2002
rect 6177 1944 6182 2000
rect 6238 1944 18142 2000
rect 18198 1944 18203 2000
rect 6177 1942 18203 1944
rect 6177 1939 6243 1942
rect 18137 1939 18203 1942
rect 23841 2002 23907 2005
rect 27520 2002 28000 2032
rect 23841 2000 28000 2002
rect 23841 1944 23846 2000
rect 23902 1944 28000 2000
rect 23841 1942 28000 1944
rect 23841 1939 23907 1942
rect 27520 1912 28000 1942
rect 8845 1866 8911 1869
rect 13997 1866 14063 1869
rect 16757 1866 16823 1869
rect 8845 1864 16823 1866
rect 8845 1808 8850 1864
rect 8906 1808 14002 1864
rect 14058 1808 16762 1864
rect 16818 1808 16823 1864
rect 8845 1806 16823 1808
rect 8845 1803 8911 1806
rect 13997 1803 14063 1806
rect 16757 1803 16823 1806
rect 289 1730 355 1733
rect 9029 1730 9095 1733
rect 16849 1730 16915 1733
rect 289 1728 6930 1730
rect 289 1672 294 1728
rect 350 1672 6930 1728
rect 289 1670 6930 1672
rect 289 1667 355 1670
rect 0 1458 480 1488
rect 3785 1458 3851 1461
rect 0 1456 3851 1458
rect 0 1400 3790 1456
rect 3846 1400 3851 1456
rect 0 1398 3851 1400
rect 6870 1458 6930 1670
rect 9029 1728 16915 1730
rect 9029 1672 9034 1728
rect 9090 1672 16854 1728
rect 16910 1672 16915 1728
rect 9029 1670 16915 1672
rect 9029 1667 9095 1670
rect 16849 1667 16915 1670
rect 23013 1730 23079 1733
rect 27613 1730 27679 1733
rect 23013 1728 27679 1730
rect 23013 1672 23018 1728
rect 23074 1672 27618 1728
rect 27674 1672 27679 1728
rect 23013 1670 27679 1672
rect 23013 1667 23079 1670
rect 27613 1667 27679 1670
rect 8017 1594 8083 1597
rect 10869 1594 10935 1597
rect 23749 1594 23815 1597
rect 8017 1592 23815 1594
rect 8017 1536 8022 1592
rect 8078 1536 10874 1592
rect 10930 1536 23754 1592
rect 23810 1536 23815 1592
rect 8017 1534 23815 1536
rect 8017 1531 8083 1534
rect 10869 1531 10935 1534
rect 23749 1531 23815 1534
rect 23933 1594 23999 1597
rect 23933 1592 26986 1594
rect 23933 1536 23938 1592
rect 23994 1536 26986 1592
rect 23933 1534 26986 1536
rect 23933 1531 23999 1534
rect 11053 1458 11119 1461
rect 6870 1456 11119 1458
rect 6870 1400 11058 1456
rect 11114 1400 11119 1456
rect 6870 1398 11119 1400
rect 0 1368 480 1398
rect 3785 1395 3851 1398
rect 11053 1395 11119 1398
rect 11605 1458 11671 1461
rect 17033 1458 17099 1461
rect 11605 1456 17099 1458
rect 11605 1400 11610 1456
rect 11666 1400 17038 1456
rect 17094 1400 17099 1456
rect 11605 1398 17099 1400
rect 11605 1395 11671 1398
rect 17033 1395 17099 1398
rect 20161 1458 20227 1461
rect 26785 1458 26851 1461
rect 20161 1456 26851 1458
rect 20161 1400 20166 1456
rect 20222 1400 26790 1456
rect 26846 1400 26851 1456
rect 20161 1398 26851 1400
rect 26926 1458 26986 1534
rect 27520 1458 28000 1488
rect 26926 1398 28000 1458
rect 20161 1395 20227 1398
rect 26785 1395 26851 1398
rect 27520 1368 28000 1398
rect 14273 1322 14339 1325
rect 14406 1322 14412 1324
rect 14273 1320 14412 1322
rect 14273 1264 14278 1320
rect 14334 1264 14412 1320
rect 14273 1262 14412 1264
rect 14273 1259 14339 1262
rect 14406 1260 14412 1262
rect 14476 1260 14482 1324
rect 0 914 480 944
rect 2865 914 2931 917
rect 0 912 2931 914
rect 0 856 2870 912
rect 2926 856 2931 912
rect 0 854 2931 856
rect 0 824 480 854
rect 2865 851 2931 854
rect 23473 914 23539 917
rect 27520 914 28000 944
rect 23473 912 28000 914
rect 23473 856 23478 912
rect 23534 856 28000 912
rect 23473 854 28000 856
rect 23473 851 23539 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 3693 370 3759 373
rect 0 368 3759 370
rect 0 312 3698 368
rect 3754 312 3759 368
rect 0 310 3759 312
rect 0 280 480 310
rect 3693 307 3759 310
rect 26141 370 26207 373
rect 27520 370 28000 400
rect 26141 368 28000 370
rect 26141 312 26146 368
rect 26202 312 28000 368
rect 26141 310 28000 312
rect 26141 307 26207 310
rect 27520 280 28000 310
rect 4613 98 4679 101
rect 24209 98 24275 101
rect 4613 96 24275 98
rect 4613 40 4618 96
rect 4674 40 24214 96
rect 24270 40 24275 96
rect 4613 38 24275 40
rect 4613 35 4679 38
rect 24209 35 24275 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 2084 16552 2148 16556
rect 2084 16496 2098 16552
rect 2098 16496 2148 16552
rect 2084 16492 2148 16496
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 6500 15948 6564 16012
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 4292 15268 4356 15332
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 19380 14784 19444 14788
rect 19380 14728 19430 14784
rect 19430 14728 19444 14784
rect 19380 14724 19444 14728
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 14412 14588 14476 14652
rect 23428 14648 23492 14652
rect 23428 14592 23478 14648
rect 23478 14592 23492 14648
rect 23428 14588 23492 14592
rect 23060 14512 23124 14516
rect 23060 14456 23074 14512
rect 23074 14456 23124 14512
rect 23060 14452 23124 14456
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 7972 13772 8036 13836
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 23612 13500 23676 13564
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 3004 13016 3068 13020
rect 3004 12960 3018 13016
rect 3018 12960 3068 13016
rect 3004 12956 3068 12960
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 13860 12820 13924 12884
rect 20484 12684 20548 12748
rect 23796 12548 23860 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 3924 12276 3988 12340
rect 23796 12276 23860 12340
rect 23980 12140 24044 12204
rect 3004 12064 3068 12068
rect 3004 12008 3054 12064
rect 3054 12008 3068 12064
rect 3004 12004 3068 12008
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 2084 11520 2148 11524
rect 2084 11464 2134 11520
rect 2134 11464 2148 11520
rect 2084 11460 2148 11464
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 19380 10780 19444 10844
rect 20484 10780 20548 10844
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 23980 10644 24044 10708
rect 11100 10432 11164 10436
rect 11100 10376 11150 10432
rect 11150 10376 11164 10432
rect 11100 10372 11164 10376
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 4292 10236 4356 10300
rect 13860 10236 13924 10300
rect 19334 10236 19398 10300
rect 6132 9964 6196 10028
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 13308 9284 13372 9348
rect 14228 9284 14292 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 3740 9148 3804 9212
rect 23060 9012 23124 9076
rect 9812 8876 9876 8940
rect 23980 8876 24044 8940
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 7972 8740 8036 8804
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 4844 8256 4908 8260
rect 4844 8200 4858 8256
rect 4858 8200 4908 8256
rect 4844 8196 4908 8200
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 2636 7788 2700 7852
rect 20300 7848 20364 7852
rect 20300 7792 20350 7848
rect 20350 7792 20364 7848
rect 20300 7788 20364 7792
rect 10916 7652 10980 7716
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 16068 7516 16132 7580
rect 6684 7108 6748 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 6316 6760 6380 6764
rect 6316 6704 6330 6760
rect 6330 6704 6380 6760
rect 6316 6700 6380 6704
rect 13308 6564 13372 6628
rect 13676 6564 13740 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 3740 6428 3804 6492
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 8708 6428 8772 6492
rect 14412 6428 14476 6492
rect 23980 6292 24044 6356
rect 14596 6156 14660 6220
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 23980 5884 24044 5948
rect 9812 5612 9876 5676
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 3372 5340 3436 5404
rect 15516 5340 15580 5404
rect 23612 5340 23676 5404
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 12756 4448 12820 4452
rect 12756 4392 12806 4448
rect 12806 4392 12820 4448
rect 12756 4388 12820 4392
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 5212 4252 5276 4316
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 23428 4448 23492 4452
rect 23428 4392 23478 4448
rect 23478 4392 23492 4448
rect 23428 4388 23492 4392
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 16620 3980 16684 4044
rect 8340 3904 8404 3908
rect 8340 3848 8354 3904
rect 8354 3848 8404 3904
rect 8340 3844 8404 3848
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 16068 3708 16132 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 1164 3164 1228 3228
rect 16620 3088 16684 3092
rect 16620 3032 16634 3088
rect 16634 3032 16684 3088
rect 16620 3028 16684 3032
rect 17356 2756 17420 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 4844 2680 4908 2684
rect 4844 2624 4894 2680
rect 4894 2624 4908 2680
rect 4844 2620 4908 2624
rect 9812 2348 9876 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 14412 1260 14476 1324
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 2083 16556 2149 16557
rect 2083 16492 2084 16556
rect 2148 16492 2149 16556
rect 2083 16491 2149 16492
rect 2086 11525 2146 16491
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 4291 15332 4357 15333
rect 4291 15268 4292 15332
rect 4356 15268 4357 15332
rect 4291 15267 4357 15268
rect 3003 13020 3069 13021
rect 3003 12956 3004 13020
rect 3068 12956 3069 13020
rect 3003 12955 3069 12956
rect 3006 12069 3066 12955
rect 3923 12340 3989 12341
rect 3923 12276 3924 12340
rect 3988 12276 3989 12340
rect 3923 12275 3989 12276
rect 3003 12068 3069 12069
rect 3003 12004 3004 12068
rect 3068 12004 3069 12068
rect 3926 12018 3986 12275
rect 3003 12003 3069 12004
rect 2083 11524 2149 11525
rect 2083 11460 2084 11524
rect 2148 11460 2149 11524
rect 2083 11459 2149 11460
rect 4294 10301 4354 15267
rect 5610 15264 5931 16288
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 6499 16012 6565 16013
rect 6499 15948 6500 16012
rect 6564 15948 6565 16012
rect 6499 15947 6565 15948
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 4291 10300 4357 10301
rect 4291 10236 4292 10300
rect 4356 10236 4357 10300
rect 4291 10235 4357 10236
rect 5610 9824 5931 10848
rect 6134 10029 6194 12462
rect 6131 10028 6197 10029
rect 6131 9964 6132 10028
rect 6196 9964 6197 10028
rect 6131 9963 6197 9964
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 4843 8260 4909 8261
rect 4843 8196 4844 8260
rect 4908 8196 4909 8260
rect 4843 8195 4909 8196
rect 3739 6492 3805 6493
rect 3739 6428 3740 6492
rect 3804 6428 3805 6492
rect 3739 6427 3805 6428
rect 3371 5404 3437 5405
rect 3371 5340 3372 5404
rect 3436 5340 3437 5404
rect 3371 5339 3437 5340
rect 3374 4538 3434 5339
rect 1166 3229 1226 3622
rect 1163 3228 1229 3229
rect 1163 3164 1164 3228
rect 1228 3164 1229 3228
rect 1163 3163 1229 3164
rect 3742 2498 3802 6427
rect 4846 2685 4906 8195
rect 5610 7648 5931 8672
rect 6502 7850 6562 15947
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 7971 13836 8037 13837
rect 7971 13772 7972 13836
rect 8036 13772 8037 13836
rect 7971 13771 8037 13772
rect 7974 8805 8034 13771
rect 10277 13632 10597 14656
rect 14411 14652 14477 14653
rect 14411 14588 14412 14652
rect 14476 14588 14477 14652
rect 14411 14587 14477 14588
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 11102 10437 11162 14502
rect 13859 12884 13925 12885
rect 13859 12820 13860 12884
rect 13924 12820 13925 12884
rect 13859 12819 13925 12820
rect 11099 10436 11165 10437
rect 11099 10372 11100 10436
rect 11164 10372 11165 10436
rect 11099 10371 11165 10372
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 13862 10301 13922 12819
rect 14414 12698 14474 14587
rect 14944 14176 15264 15200
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19379 14788 19445 14789
rect 19379 14724 19380 14788
rect 19444 14724 19445 14788
rect 19379 14723 19445 14724
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 13859 10300 13925 10301
rect 13859 10236 13860 10300
rect 13924 10236 13925 10300
rect 13859 10235 13925 10236
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 9811 8940 9877 8941
rect 9811 8876 9812 8940
rect 9876 8876 9877 8940
rect 9811 8875 9877 8876
rect 7971 8804 8037 8805
rect 7971 8740 7972 8804
rect 8036 8740 8037 8804
rect 7971 8739 8037 8740
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 6318 7790 6562 7850
rect 6318 6765 6378 7790
rect 6315 6764 6381 6765
rect 6315 6700 6316 6764
rect 6380 6700 6381 6764
rect 6315 6699 6381 6700
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 9814 5677 9874 8875
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10918 7717 10978 9742
rect 13307 9348 13373 9349
rect 13307 9284 13308 9348
rect 13372 9284 13373 9348
rect 14227 9348 14293 9349
rect 14227 9298 14228 9348
rect 14292 9298 14293 9348
rect 13307 9283 13373 9284
rect 10915 7716 10981 7717
rect 10915 7652 10916 7716
rect 10980 7652 10981 7716
rect 10915 7651 10981 7652
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 13310 6629 13370 9283
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 13307 6628 13373 6629
rect 13307 6564 13308 6628
rect 13372 6564 13373 6628
rect 13307 6563 13373 6564
rect 13675 6628 13741 6629
rect 13675 6564 13676 6628
rect 13740 6564 13741 6628
rect 13675 6563 13741 6564
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 9811 5676 9877 5677
rect 9811 5612 9812 5676
rect 9876 5612 9877 5676
rect 9811 5611 9877 5612
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5214 4317 5274 4982
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5211 4316 5277 4317
rect 5211 4252 5212 4316
rect 5276 4252 5277 4316
rect 5211 4251 5277 4252
rect 5610 3296 5931 4320
rect 8339 3908 8405 3909
rect 8339 3844 8340 3908
rect 8404 3844 8405 3908
rect 8339 3843 8405 3844
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 4843 2684 4909 2685
rect 4843 2620 4844 2684
rect 4908 2620 4909 2684
rect 4843 2619 4909 2620
rect 5610 2208 5931 3232
rect 8342 3178 8402 3843
rect 9814 2413 9874 5611
rect 10277 4928 10597 5952
rect 13678 5898 13738 6563
rect 14411 6492 14477 6493
rect 14411 6428 14412 6492
rect 14476 6428 14477 6492
rect 14411 6427 14477 6428
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 12755 4452 12821 4453
rect 12755 4388 12756 4452
rect 12820 4388 12821 4452
rect 12755 4387 12821 4388
rect 12758 3858 12818 4387
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 9811 2412 9877 2413
rect 9811 2348 9812 2412
rect 9876 2348 9877 2412
rect 9811 2347 9877 2348
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2128 10597 2688
rect 14414 1325 14474 6427
rect 14598 6221 14658 7022
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14595 6220 14661 6221
rect 14595 6156 14596 6220
rect 14660 6156 14661 6220
rect 14595 6155 14661 6156
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 15518 5405 15578 11782
rect 16070 7581 16130 11102
rect 19382 10845 19442 14723
rect 19610 14720 19930 15744
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 23059 14516 23125 14517
rect 23059 14452 23060 14516
rect 23124 14452 23125 14516
rect 23059 14451 23125 14452
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 20483 12748 20549 12749
rect 20483 12684 20484 12748
rect 20548 12684 20549 12748
rect 20483 12683 20549 12684
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19379 10844 19445 10845
rect 19379 10780 19380 10844
rect 19444 10780 19445 10844
rect 19379 10779 19445 10780
rect 19382 10570 19442 10779
rect 19336 10510 19442 10570
rect 19336 10301 19396 10510
rect 19610 10368 19930 11392
rect 20486 10845 20546 12683
rect 20483 10844 20549 10845
rect 20483 10780 20484 10844
rect 20548 10780 20549 10844
rect 20483 10779 20549 10780
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19333 10300 19399 10301
rect 19333 10236 19334 10300
rect 19398 10236 19399 10300
rect 19333 10235 19399 10236
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 16067 7580 16133 7581
rect 16067 7516 16068 7580
rect 16132 7516 16133 7580
rect 16067 7515 16133 7516
rect 15515 5404 15581 5405
rect 15515 5340 15516 5404
rect 15580 5340 15581 5404
rect 15515 5339 15581 5340
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 16070 3773 16130 7515
rect 16438 5218 16498 9062
rect 19610 8192 19930 9216
rect 23062 9077 23122 14451
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23611 13564 23677 13565
rect 23611 13500 23612 13564
rect 23676 13500 23677 13564
rect 23611 13499 23677 13500
rect 23059 9076 23125 9077
rect 23059 9012 23060 9076
rect 23124 9012 23125 9076
rect 23059 9011 23125 9012
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 23614 5405 23674 13499
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23795 12612 23861 12613
rect 23795 12548 23796 12612
rect 23860 12548 23861 12612
rect 23795 12547 23861 12548
rect 23798 12341 23858 12547
rect 23795 12340 23861 12341
rect 23795 12276 23796 12340
rect 23860 12276 23861 12340
rect 23795 12275 23861 12276
rect 23979 12204 24045 12205
rect 23979 12140 23980 12204
rect 24044 12140 24045 12204
rect 23979 12139 24045 12140
rect 23982 11338 24042 12139
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23979 10708 24045 10709
rect 23979 10644 23980 10708
rect 24044 10644 24045 10708
rect 23979 10643 24045 10644
rect 23982 9978 24042 10643
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 23982 8941 24042 9062
rect 23979 8940 24045 8941
rect 23979 8876 23980 8940
rect 24044 8876 24045 8940
rect 23979 8875 24045 8876
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 23979 6292 23980 6342
rect 24044 6292 24045 6342
rect 23979 6291 24045 6292
rect 23979 5948 24045 5949
rect 23979 5898 23980 5948
rect 24044 5898 24045 5948
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23611 5404 23677 5405
rect 23611 5340 23612 5404
rect 23676 5340 23677 5404
rect 23611 5339 23677 5340
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 16619 4044 16685 4045
rect 16619 3980 16620 4044
rect 16684 3980 16685 4044
rect 16619 3979 16685 3980
rect 16622 3858 16682 3979
rect 16067 3772 16133 3773
rect 16067 3708 16068 3772
rect 16132 3708 16133 3772
rect 16067 3707 16133 3708
rect 19610 3840 19930 4864
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 17355 2820 17421 2821
rect 17355 2756 17356 2820
rect 17420 2756 17421 2820
rect 17355 2755 17421 2756
rect 17358 2498 17418 2755
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2128 19930 2688
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 14411 1324 14477 1325
rect 14411 1260 14412 1324
rect 14476 1260 14477 1324
rect 14411 1259 14477 1260
<< via4 >>
rect 3838 11782 4074 12018
rect 6046 12462 6282 12698
rect 3654 9212 3890 9298
rect 3654 9148 3740 9212
rect 3740 9148 3804 9212
rect 3804 9148 3890 9212
rect 3654 9062 3890 9148
rect 2550 7852 2786 7938
rect 2550 7788 2636 7852
rect 2636 7788 2700 7852
rect 2700 7788 2786 7852
rect 2550 7702 2786 7788
rect 3286 4302 3522 4538
rect 1078 3622 1314 3858
rect 11014 14502 11250 14738
rect 14326 12462 14562 12698
rect 15430 11782 15666 12018
rect 10830 9742 11066 9978
rect 6598 7172 6834 7258
rect 6598 7108 6684 7172
rect 6684 7108 6748 7172
rect 6748 7108 6834 7172
rect 6598 7022 6834 7108
rect 8622 6492 8858 6578
rect 8622 6428 8708 6492
rect 8708 6428 8772 6492
rect 8772 6428 8858 6492
rect 8622 6342 8858 6428
rect 14142 9284 14228 9298
rect 14228 9284 14292 9298
rect 14292 9284 14378 9298
rect 14142 9062 14378 9284
rect 14510 7022 14746 7258
rect 5126 4982 5362 5218
rect 3654 2262 3890 2498
rect 8254 2942 8490 3178
rect 13590 5662 13826 5898
rect 12670 3622 12906 3858
rect 15982 11102 16218 11338
rect 23342 14652 23578 14738
rect 23342 14588 23428 14652
rect 23428 14588 23492 14652
rect 23492 14588 23578 14652
rect 23342 14502 23578 14588
rect 16350 9062 16586 9298
rect 20214 7852 20450 7938
rect 20214 7788 20300 7852
rect 20300 7788 20364 7852
rect 20364 7788 20450 7852
rect 20214 7702 20450 7788
rect 16350 4982 16586 5218
rect 23894 11102 24130 11338
rect 23894 9742 24130 9978
rect 23894 9062 24130 9298
rect 23894 6356 24130 6578
rect 23894 6342 23980 6356
rect 23980 6342 24044 6356
rect 24044 6342 24130 6356
rect 23894 5884 23980 5898
rect 23980 5884 24044 5898
rect 24044 5884 24130 5898
rect 23894 5662 24130 5884
rect 16534 3622 16770 3858
rect 23342 4452 23578 4538
rect 23342 4388 23428 4452
rect 23428 4388 23492 4452
rect 23492 4388 23578 4452
rect 23342 4302 23578 4388
rect 16534 3092 16770 3178
rect 16534 3028 16620 3092
rect 16620 3028 16684 3092
rect 16684 3028 16770 3092
rect 16534 2942 16770 3028
rect 17270 2262 17506 2498
<< metal5 >>
rect 10972 14738 23620 14780
rect 10972 14502 11014 14738
rect 11250 14502 23342 14738
rect 23578 14502 23620 14738
rect 10972 14460 23620 14502
rect 6004 12698 14604 12740
rect 6004 12462 6046 12698
rect 6282 12462 14326 12698
rect 14562 12462 14604 12698
rect 6004 12420 14604 12462
rect 3796 12018 15708 12060
rect 3796 11782 3838 12018
rect 4074 11782 15430 12018
rect 15666 11782 15708 12018
rect 3796 11740 15708 11782
rect 15940 11338 24172 11380
rect 15940 11102 15982 11338
rect 16218 11102 23894 11338
rect 24130 11102 24172 11338
rect 15940 11060 24172 11102
rect 10788 9978 24172 10020
rect 10788 9742 10830 9978
rect 11066 9742 23894 9978
rect 24130 9742 24172 9978
rect 10788 9700 24172 9742
rect 3612 9298 14420 9340
rect 3612 9062 3654 9298
rect 3890 9062 14142 9298
rect 14378 9062 14420 9298
rect 3612 9020 14420 9062
rect 16308 9298 24172 9340
rect 16308 9062 16350 9298
rect 16586 9062 23894 9298
rect 24130 9062 24172 9298
rect 16308 9020 24172 9062
rect 2508 7938 20492 7980
rect 2508 7702 2550 7938
rect 2786 7702 20214 7938
rect 20450 7702 20492 7938
rect 2508 7660 20492 7702
rect 6556 7258 14788 7300
rect 6556 7022 6598 7258
rect 6834 7022 14510 7258
rect 14746 7022 14788 7258
rect 6556 6980 14788 7022
rect 8580 6578 24172 6620
rect 8580 6342 8622 6578
rect 8858 6342 23894 6578
rect 24130 6342 24172 6578
rect 8580 6300 24172 6342
rect 13548 5898 24172 5940
rect 13548 5662 13590 5898
rect 13826 5662 23894 5898
rect 24130 5662 24172 5898
rect 13548 5620 24172 5662
rect 5084 5218 16628 5260
rect 5084 4982 5126 5218
rect 5362 4982 16350 5218
rect 16586 4982 16628 5218
rect 5084 4940 16628 4982
rect 3244 4538 23620 4580
rect 3244 4302 3286 4538
rect 3522 4302 23342 4538
rect 23578 4302 23620 4538
rect 3244 4260 23620 4302
rect 1036 3858 16812 3900
rect 1036 3622 1078 3858
rect 1314 3622 12670 3858
rect 12906 3622 16534 3858
rect 16770 3622 16812 3858
rect 1036 3580 16812 3622
rect 8212 3178 16812 3220
rect 8212 2942 8254 3178
rect 8490 2942 16534 3178
rect 16770 2942 16812 3178
rect 8212 2900 16812 2942
rect 3612 2498 17548 2540
rect 3612 2262 3654 2498
rect 3890 2262 17270 2498
rect 17506 2262 17548 2498
rect 3612 2220 17548 2262
use sky130_fd_sc_hd__decap_3  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1604681595
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1604681595
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_1_47
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_43
timestamp 1604681595
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_52
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_71
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1604681595
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_80
timestamp 1604681595
transform 1 0 8464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_103
timestamp 1604681595
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1604681595
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1604681595
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1604681595
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1604681595
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_156
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16192 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1604681595
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_204
timestamp 1604681595
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18400 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_228
timestamp 1604681595
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 20608 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_236
timestamp 1604681595
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_235
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_261
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_273
timestamp 1604681595
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1472 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1604681595
transform 1 0 2300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_17
timestamp 1604681595
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_21
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1604681595
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_83
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1604681595
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1604681595
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_114
timestamp 1604681595
transform 1 0 11592 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1604681595
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1604681595
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_194
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21804 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_223
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604681595
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604681595
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1472 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_21
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1604681595
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_87
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_108
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_112
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_153
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_156
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_207
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_272
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_14
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1604681595
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_25
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_22
timestamp 1604681595
transform 1 0 3128 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1604681595
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_173
timestamp 1604681595
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1604681595
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1604681595
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_228
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_33
timestamp 1604681595
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1604681595
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1604681595
transform 1 0 8464 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_103
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1604681595
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_192
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_213
timestamp 1604681595
transform 1 0 20700 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23276 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_235
timestamp 1604681595
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_239
timestamp 1604681595
transform 1 0 23092 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604681595
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_261
timestamp 1604681595
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_265
timestamp 1604681595
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_273
timestamp 1604681595
transform 1 0 26220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1656 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1604681595
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1604681595
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_22
timestamp 1604681595
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_33
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1604681595
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1604681595
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_83
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 1604681595
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_126
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_154
timestamp 1604681595
transform 1 0 15272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1604681595
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1604681595
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 1604681595
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1604681595
transform 1 0 20148 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_211
timestamp 1604681595
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_227
timestamp 1604681595
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_223
timestamp 1604681595
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1604681595
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23092 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 22356 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1604681595
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_254
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_258
timestamp 1604681595
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1604681595
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_272
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1656 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_35
timestamp 1604681595
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 1604681595
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9936 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1604681595
transform 1 0 15824 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_164
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_189
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1604681595
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_235
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_255
timestamp 1604681595
transform 1 0 24564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp 1604681595
transform 1 0 24932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1604681595
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_10
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6900 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_72
timestamp 1604681595
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_80
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1604681595
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 16100 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp 1604681595
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_217
timestamp 1604681595
transform 1 0 21068 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_251
timestamp 1604681595
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1604681595
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_268
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_272
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1604681595
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 5888 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1604681595
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_103
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1604681595
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 18676 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1604681595
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21804 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1604681595
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_222
timestamp 1604681595
transform 1 0 21528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1604681595
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_238
timestamp 1604681595
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 24932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_257
timestamp 1604681595
transform 1 0 24748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1604681595
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1604681595
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1604681595
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_73
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1604681595
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_151
timestamp 1604681595
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1604681595
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 20976 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_261
timestamp 1604681595
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_265
timestamp 1604681595
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_273
timestamp 1604681595
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604681595
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4140 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604681595
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1604681595
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_96
timestamp 1604681595
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1604681595
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1604681595
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21344 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1604681595
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_229
timestamp 1604681595
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_233
timestamp 1604681595
transform 1 0 22540 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_238
timestamp 1604681595
transform 1 0 23000 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 25024 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_252
timestamp 1604681595
transform 1 0 24288 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_256
timestamp 1604681595
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_264
timestamp 1604681595
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_268 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_18
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_14
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1656 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_31
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1604681595
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1604681595
transform 1 0 6348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_144
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 21252 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22816 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_249
timestamp 1604681595
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1604681595
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23736 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_262
timestamp 1604681595
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_266
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_262
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_270
timestamp 1604681595
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_270
timestamp 1604681595
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_274
timestamp 1604681595
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4508 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1604681595
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 12604 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_218
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_223
timestamp 1604681595
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23920 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604681595
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_272
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1604681595
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_20
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_24
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_81
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_101
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_96
timestamp 1604681595
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_120
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_133
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_147
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_196
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 21804 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1604681595
transform 1 0 21252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_234
timestamp 1604681595
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_238
timestamp 1604681595
transform 1 0 23000 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_252
timestamp 1604681595
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_256
timestamp 1604681595
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_264
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_268
timestamp 1604681595
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_55
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_205
timestamp 1604681595
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1604681595
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_229
timestamp 1604681595
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23920 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1604681595
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1604681595
transform 1 0 22908 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_268
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_272
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1604681595
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_24
timestamp 1604681595
transform 1 0 3312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_86
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_125
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_148
timestamp 1604681595
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1604681595
transform 1 0 16008 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1604681595
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1604681595
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_225
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_229
timestamp 1604681595
transform 1 0 22172 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_243
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_57
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_79
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_108
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1604681595
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1604681595
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_160
timestamp 1604681595
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1604681595
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_192
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_207
timestamp 1604681595
transform 1 0 20148 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1604681595
transform 1 0 19780 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21344 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_237
timestamp 1604681595
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_233
timestamp 1604681595
transform 1 0 22540 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22724 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_255
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1604681595
transform 1 0 24840 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_262
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_52
timestamp 1604681595
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_56
timestamp 1604681595
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_115
timestamp 1604681595
transform 1 0 11684 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15548 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_153
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_166
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_170
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1604681595
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_234
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_262
timestamp 1604681595
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_266
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_274
timestamp 1604681595
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_49
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1604681595
transform 1 0 5980 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_63
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_87
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1604681595
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_120
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1604681595
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_180
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_184
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1604681595
transform 1 0 18492 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21160 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23368 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1604681595
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_262
timestamp 1604681595
transform 1 0 25208 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4508 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_46
timestamp 1604681595
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_55
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 8096 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1604681595
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1604681595
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1604681595
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_91
timestamp 1604681595
transform 1 0 9476 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_160
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17664 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_173
timestamp 1604681595
transform 1 0 17020 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1604681595
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19872 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1604681595
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_226
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_272
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1604681595
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1604681595
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1604681595
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604681595
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1604681595
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_167
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1604681595
transform 1 0 17296 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1604681595
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23276 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22724 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_233
timestamp 1604681595
transform 1 0 22540 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1604681595
transform 1 0 22908 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1604681595
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_254
timestamp 1604681595
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_264
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1604681595
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 3036 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_52
timestamp 1604681595
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_44
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604681595
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_56
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_105
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 15548 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_187
timestamp 1604681595
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_198
timestamp 1604681595
transform 1 0 19320 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_270
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 1472 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 1564 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_19
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_14
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_13
timestamp 1604681595
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604681595
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_60
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_48
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_72
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12696 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_138
timestamp 1604681595
transform 1 0 13800 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1604681595
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_150
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_162
timestamp 1604681595
transform 1 0 16008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_176
timestamp 1604681595
transform 1 0 17296 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_195
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 18768 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_188
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20976 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1604681595
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_229
timestamp 1604681595
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1604681595
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1604681595
transform 1 0 24012 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_255
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604681595
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1604681595
transform 1 0 2300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_25
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_60
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_131
timestamp 1604681595
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17112 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_192
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1604681595
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21068 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_223
timestamp 1604681595
transform 1 0 21620 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 23460 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 22356 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_235
timestamp 1604681595
transform 1 0 22724 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_23
timestamp 1604681595
transform 1 0 3220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_46
timestamp 1604681595
transform 1 0 5336 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_188
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_200
timestamp 1604681595
transform 1 0 19504 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_212
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_224
timestamp 1604681595
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1604681595
transform 1 0 24012 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1604681595
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_263
timestamp 1604681595
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_275
timestamp 1604681595
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_19
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_38
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_50
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_74
timestamp 1604681595
transform 1 0 7912 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_188
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_200
timestamp 1604681595
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_231
timestamp 1604681595
transform 1 0 22356 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_259
timestamp 1604681595
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1604681595
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_19
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_259
timestamp 1604681595
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1604681595
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_13
timestamp 1604681595
transform 1 0 2300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_25
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_217
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_221
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_221
timestamp 1604681595
transform 1 0 21436 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 21528 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_226
timestamp 1604681595
transform 1 0 21896 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_224
timestamp 1604681595
transform 1 0 21712 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_35
timestamp 1604681595
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_47
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604681595
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_11
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_23
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_35
timestamp 1604681595
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_47
timestamp 1604681595
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1604681595
transform 1 0 24196 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1604681595
transform 1 0 25668 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_275
timestamp 1604681595
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604681595
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 24490 27520 24546 28000 6 SC_IN_BOT
port 0 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27066 0 27122 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3606 0 3662 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 4158 0 4214 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 ccff_head
port 12 nsew default input
rlabel metal2 s 17498 27520 17554 28000 6 ccff_tail
port 13 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[0]
port 14 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[10]
port 15 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[11]
port 16 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[12]
port 17 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[13]
port 18 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[14]
port 19 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[15]
port 20 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[16]
port 21 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[17]
port 22 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chanx_left_in[18]
port 23 nsew default input
rlabel metal3 s 0 15648 480 15768 6 chanx_left_in[19]
port 24 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[1]
port 25 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 26 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[3]
port 27 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[4]
port 28 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[5]
port 29 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[6]
port 30 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[7]
port 31 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[8]
port 32 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[9]
port 33 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[0]
port 34 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[10]
port 35 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[11]
port 36 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[12]
port 37 nsew default tristate
rlabel metal3 s 0 23672 480 23792 6 chanx_left_out[13]
port 38 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[14]
port 39 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[15]
port 40 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[16]
port 41 nsew default tristate
rlabel metal3 s 0 25984 480 26104 6 chanx_left_out[17]
port 42 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[18]
port 43 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[19]
port 44 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[1]
port 45 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[2]
port 46 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[3]
port 47 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 48 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 49 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[6]
port 50 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 51 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[8]
port 52 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[9]
port 53 nsew default tristate
rlabel metal3 s 27520 4632 28000 4752 6 chanx_right_in[0]
port 54 nsew default input
rlabel metal3 s 27520 10344 28000 10464 6 chanx_right_in[10]
port 55 nsew default input
rlabel metal3 s 27520 10888 28000 11008 6 chanx_right_in[11]
port 56 nsew default input
rlabel metal3 s 27520 11432 28000 11552 6 chanx_right_in[12]
port 57 nsew default input
rlabel metal3 s 27520 11976 28000 12096 6 chanx_right_in[13]
port 58 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[14]
port 59 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[15]
port 60 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[16]
port 61 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[17]
port 62 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[18]
port 63 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[19]
port 64 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 65 nsew default input
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_in[2]
port 66 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[3]
port 67 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[4]
port 68 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_in[5]
port 69 nsew default input
rlabel metal3 s 27520 8032 28000 8152 6 chanx_right_in[6]
port 70 nsew default input
rlabel metal3 s 27520 8576 28000 8696 6 chanx_right_in[7]
port 71 nsew default input
rlabel metal3 s 27520 9120 28000 9240 6 chanx_right_in[8]
port 72 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[9]
port 73 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[0]
port 74 nsew default tristate
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_out[10]
port 75 nsew default tristate
rlabel metal3 s 27520 22040 28000 22160 6 chanx_right_out[11]
port 76 nsew default tristate
rlabel metal3 s 27520 22584 28000 22704 6 chanx_right_out[12]
port 77 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[13]
port 78 nsew default tristate
rlabel metal3 s 27520 23808 28000 23928 6 chanx_right_out[14]
port 79 nsew default tristate
rlabel metal3 s 27520 24352 28000 24472 6 chanx_right_out[15]
port 80 nsew default tristate
rlabel metal3 s 27520 24896 28000 25016 6 chanx_right_out[16]
port 81 nsew default tristate
rlabel metal3 s 27520 25440 28000 25560 6 chanx_right_out[17]
port 82 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[18]
port 83 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[19]
port 84 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chanx_right_out[1]
port 85 nsew default tristate
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_out[2]
port 86 nsew default tristate
rlabel metal3 s 27520 17552 28000 17672 6 chanx_right_out[3]
port 87 nsew default tristate
rlabel metal3 s 27520 18096 28000 18216 6 chanx_right_out[4]
port 88 nsew default tristate
rlabel metal3 s 27520 18640 28000 18760 6 chanx_right_out[5]
port 89 nsew default tristate
rlabel metal3 s 27520 19320 28000 19440 6 chanx_right_out[6]
port 90 nsew default tristate
rlabel metal3 s 27520 19864 28000 19984 6 chanx_right_out[7]
port 91 nsew default tristate
rlabel metal3 s 27520 20408 28000 20528 6 chanx_right_out[8]
port 92 nsew default tristate
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_out[9]
port 93 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[0]
port 94 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 95 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[11]
port 96 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[12]
port 97 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[13]
port 98 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[14]
port 99 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[15]
port 100 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[16]
port 101 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[17]
port 102 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[18]
port 103 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[19]
port 104 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[1]
port 105 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[2]
port 106 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[3]
port 107 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[4]
port 108 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[5]
port 109 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[6]
port 110 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[7]
port 111 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[8]
port 112 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[9]
port 113 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[0]
port 114 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[10]
port 115 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 116 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[12]
port 117 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[13]
port 118 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[14]
port 119 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[15]
port 120 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[16]
port 121 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[17]
port 122 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[18]
port 123 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[19]
port 124 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[1]
port 125 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[2]
port 126 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[3]
port 127 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[4]
port 128 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[5]
port 129 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[6]
port 130 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[7]
port 131 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[8]
port 132 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[9]
port 133 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 134 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 135 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 136 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 137 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_38_
port 138 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 139 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 140 nsew default input
rlabel metal3 s 0 4224 480 4344 6 left_bottom_grid_pin_41_
port 141 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_1_
port 142 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 prog_clk
port 143 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 144 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 145 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 146 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 147 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 148 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 right_bottom_grid_pin_39_
port 149 nsew default input
rlabel metal3 s 27520 3544 28000 3664 6 right_bottom_grid_pin_40_
port 150 nsew default input
rlabel metal3 s 27520 4088 28000 4208 6 right_bottom_grid_pin_41_
port 151 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_1_
port 152 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 153 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 154 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
