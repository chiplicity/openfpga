magic
tech sky130A
magscale 1 2
timestamp 1608157018
<< obsli1 >>
rect 1104 1377 22235 20145
<< obsm1 >>
rect 198 1164 22618 20664
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 938 22000 994 22800
rect 1306 22000 1362 22800
rect 1674 22000 1730 22800
rect 2042 22000 2098 22800
rect 2410 22000 2466 22800
rect 2778 22000 2834 22800
rect 3238 22000 3294 22800
rect 3606 22000 3662 22800
rect 3974 22000 4030 22800
rect 4342 22000 4398 22800
rect 4710 22000 4766 22800
rect 5078 22000 5134 22800
rect 5446 22000 5502 22800
rect 5906 22000 5962 22800
rect 6274 22000 6330 22800
rect 6642 22000 6698 22800
rect 7010 22000 7066 22800
rect 7378 22000 7434 22800
rect 7746 22000 7802 22800
rect 8114 22000 8170 22800
rect 8482 22000 8538 22800
rect 8942 22000 8998 22800
rect 9310 22000 9366 22800
rect 9678 22000 9734 22800
rect 10046 22000 10102 22800
rect 10414 22000 10470 22800
rect 10782 22000 10838 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12346 22000 12402 22800
rect 12714 22000 12770 22800
rect 13082 22000 13138 22800
rect 13450 22000 13506 22800
rect 13818 22000 13874 22800
rect 14186 22000 14242 22800
rect 14646 22000 14702 22800
rect 15014 22000 15070 22800
rect 15382 22000 15438 22800
rect 15750 22000 15806 22800
rect 16118 22000 16174 22800
rect 16486 22000 16542 22800
rect 16854 22000 16910 22800
rect 17314 22000 17370 22800
rect 17682 22000 17738 22800
rect 18050 22000 18106 22800
rect 18418 22000 18474 22800
rect 18786 22000 18842 22800
rect 19154 22000 19210 22800
rect 19522 22000 19578 22800
rect 19890 22000 19946 22800
rect 20350 22000 20406 22800
rect 20718 22000 20774 22800
rect 21086 22000 21142 22800
rect 21454 22000 21510 22800
rect 21822 22000 21878 22800
rect 22190 22000 22246 22800
rect 22558 22000 22614 22800
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
<< obsm2 >>
rect 314 21944 514 22681
rect 682 21944 882 22681
rect 1050 21944 1250 22681
rect 1418 21944 1618 22681
rect 1786 21944 1986 22681
rect 2154 21944 2354 22681
rect 2522 21944 2722 22681
rect 2890 21944 3182 22681
rect 3350 21944 3550 22681
rect 3718 21944 3918 22681
rect 4086 21944 4286 22681
rect 4454 21944 4654 22681
rect 4822 21944 5022 22681
rect 5190 21944 5390 22681
rect 5558 21944 5850 22681
rect 6018 21944 6218 22681
rect 6386 21944 6586 22681
rect 6754 21944 6954 22681
rect 7122 21944 7322 22681
rect 7490 21944 7690 22681
rect 7858 21944 8058 22681
rect 8226 21944 8426 22681
rect 8594 21944 8886 22681
rect 9054 21944 9254 22681
rect 9422 21944 9622 22681
rect 9790 21944 9990 22681
rect 10158 21944 10358 22681
rect 10526 21944 10726 22681
rect 10894 21944 11094 22681
rect 11262 21944 11554 22681
rect 11722 21944 11922 22681
rect 12090 21944 12290 22681
rect 12458 21944 12658 22681
rect 12826 21944 13026 22681
rect 13194 21944 13394 22681
rect 13562 21944 13762 22681
rect 13930 21944 14130 22681
rect 14298 21944 14590 22681
rect 14758 21944 14958 22681
rect 15126 21944 15326 22681
rect 15494 21944 15694 22681
rect 15862 21944 16062 22681
rect 16230 21944 16430 22681
rect 16598 21944 16798 22681
rect 16966 21944 17258 22681
rect 17426 21944 17626 22681
rect 17794 21944 17994 22681
rect 18162 21944 18362 22681
rect 18530 21944 18730 22681
rect 18898 21944 19098 22681
rect 19266 21944 19466 22681
rect 19634 21944 19834 22681
rect 20002 21944 20294 22681
rect 20462 21944 20662 22681
rect 20830 21944 21030 22681
rect 21198 21944 21398 22681
rect 21566 21944 21766 22681
rect 21934 21944 22134 22681
rect 22302 21944 22502 22681
rect 204 856 22612 21944
rect 314 167 514 856
rect 682 167 882 856
rect 1050 167 1250 856
rect 1418 167 1618 856
rect 1786 167 1986 856
rect 2154 167 2354 856
rect 2522 167 2722 856
rect 2890 167 3090 856
rect 3258 167 3458 856
rect 3626 167 3826 856
rect 3994 167 4194 856
rect 4362 167 4562 856
rect 4730 167 4930 856
rect 5098 167 5298 856
rect 5466 167 5666 856
rect 5834 167 6126 856
rect 6294 167 6494 856
rect 6662 167 6862 856
rect 7030 167 7230 856
rect 7398 167 7598 856
rect 7766 167 7966 856
rect 8134 167 8334 856
rect 8502 167 8702 856
rect 8870 167 9070 856
rect 9238 167 9438 856
rect 9606 167 9806 856
rect 9974 167 10174 856
rect 10342 167 10542 856
rect 10710 167 10910 856
rect 11078 167 11278 856
rect 11446 167 11738 856
rect 11906 167 12106 856
rect 12274 167 12474 856
rect 12642 167 12842 856
rect 13010 167 13210 856
rect 13378 167 13578 856
rect 13746 167 13946 856
rect 14114 167 14314 856
rect 14482 167 14682 856
rect 14850 167 15050 856
rect 15218 167 15418 856
rect 15586 167 15786 856
rect 15954 167 16154 856
rect 16322 167 16522 856
rect 16690 167 16890 856
rect 17058 167 17350 856
rect 17518 167 17718 856
rect 17886 167 18086 856
rect 18254 167 18454 856
rect 18622 167 18822 856
rect 18990 167 19190 856
rect 19358 167 19558 856
rect 19726 167 19926 856
rect 20094 167 20294 856
rect 20462 167 20662 856
rect 20830 167 21030 856
rect 21198 167 21398 856
rect 21566 167 21766 856
rect 21934 167 22134 856
rect 22302 167 22502 856
<< metal3 >>
rect 0 22584 800 22704
rect 22000 22584 22800 22704
rect 0 22176 800 22296
rect 22000 22176 22800 22296
rect 0 21768 800 21888
rect 22000 21768 22800 21888
rect 0 21360 800 21480
rect 22000 21360 22800 21480
rect 0 20952 800 21072
rect 22000 20952 22800 21072
rect 0 20544 800 20664
rect 22000 20544 22800 20664
rect 0 20136 800 20256
rect 22000 20136 22800 20256
rect 0 19728 800 19848
rect 22000 19728 22800 19848
rect 0 19320 800 19440
rect 0 19048 800 19168
rect 22000 19320 22800 19440
rect 22000 19048 22800 19168
rect 0 18640 800 18760
rect 22000 18640 22800 18760
rect 0 18232 800 18352
rect 22000 18232 22800 18352
rect 0 17824 800 17944
rect 22000 17824 22800 17944
rect 0 17416 800 17536
rect 22000 17416 22800 17536
rect 0 17008 800 17128
rect 22000 17008 22800 17128
rect 0 16600 800 16720
rect 22000 16600 22800 16720
rect 0 16192 800 16312
rect 22000 16192 22800 16312
rect 0 15784 800 15904
rect 22000 15784 22800 15904
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 22000 15376 22800 15496
rect 22000 15104 22800 15224
rect 0 14696 800 14816
rect 22000 14696 22800 14816
rect 0 14288 800 14408
rect 22000 14288 22800 14408
rect 0 13880 800 14000
rect 22000 13880 22800 14000
rect 0 13472 800 13592
rect 22000 13472 22800 13592
rect 0 13064 800 13184
rect 22000 13064 22800 13184
rect 0 12656 800 12776
rect 22000 12656 22800 12776
rect 0 12248 800 12368
rect 22000 12248 22800 12368
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 22000 11840 22800 11960
rect 22000 11568 22800 11688
rect 0 11160 800 11280
rect 22000 11160 22800 11280
rect 0 10752 800 10872
rect 22000 10752 22800 10872
rect 0 10344 800 10464
rect 22000 10344 22800 10464
rect 0 9936 800 10056
rect 22000 9936 22800 10056
rect 0 9528 800 9648
rect 22000 9528 22800 9648
rect 0 9120 800 9240
rect 22000 9120 22800 9240
rect 0 8712 800 8832
rect 22000 8712 22800 8832
rect 0 8304 800 8424
rect 22000 8304 22800 8424
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 22000 7896 22800 8016
rect 22000 7624 22800 7744
rect 0 7216 800 7336
rect 22000 7216 22800 7336
rect 0 6808 800 6928
rect 22000 6808 22800 6928
rect 0 6400 800 6520
rect 22000 6400 22800 6520
rect 0 5992 800 6112
rect 22000 5992 22800 6112
rect 0 5584 800 5704
rect 22000 5584 22800 5704
rect 0 5176 800 5296
rect 22000 5176 22800 5296
rect 0 4768 800 4888
rect 22000 4768 22800 4888
rect 0 4360 800 4480
rect 22000 4360 22800 4480
rect 0 3952 800 4072
rect 0 3680 800 3800
rect 22000 3952 22800 4072
rect 22000 3680 22800 3800
rect 0 3272 800 3392
rect 22000 3272 22800 3392
rect 0 2864 800 2984
rect 22000 2864 22800 2984
rect 0 2456 800 2576
rect 22000 2456 22800 2576
rect 0 2048 800 2168
rect 22000 2048 22800 2168
rect 0 1640 800 1760
rect 22000 1640 22800 1760
rect 0 1232 800 1352
rect 22000 1232 22800 1352
rect 0 824 800 944
rect 22000 824 22800 944
rect 0 416 800 536
rect 0 144 800 264
rect 22000 416 22800 536
rect 22000 144 22800 264
<< obsm3 >>
rect 880 22504 21920 22677
rect 800 22376 22018 22504
rect 880 22096 21920 22376
rect 800 21968 22018 22096
rect 880 21688 21920 21968
rect 800 21560 22018 21688
rect 880 21280 21920 21560
rect 800 21152 22018 21280
rect 880 20872 21920 21152
rect 800 20744 22018 20872
rect 880 20464 21920 20744
rect 800 20336 22018 20464
rect 880 20056 21920 20336
rect 800 19928 22018 20056
rect 880 19648 21920 19928
rect 800 19520 22018 19648
rect 880 18968 21920 19520
rect 800 18840 22018 18968
rect 880 18560 21920 18840
rect 800 18432 22018 18560
rect 880 18152 21920 18432
rect 800 18024 22018 18152
rect 880 17744 21920 18024
rect 800 17616 22018 17744
rect 880 17336 21920 17616
rect 800 17208 22018 17336
rect 880 16928 21920 17208
rect 800 16800 22018 16928
rect 880 16520 21920 16800
rect 800 16392 22018 16520
rect 880 16112 21920 16392
rect 800 15984 22018 16112
rect 880 15704 21920 15984
rect 800 15576 22018 15704
rect 880 15024 21920 15576
rect 800 14896 22018 15024
rect 880 14616 21920 14896
rect 800 14488 22018 14616
rect 880 14208 21920 14488
rect 800 14080 22018 14208
rect 880 13800 21920 14080
rect 800 13672 22018 13800
rect 880 13392 21920 13672
rect 800 13264 22018 13392
rect 880 12984 21920 13264
rect 800 12856 22018 12984
rect 880 12576 21920 12856
rect 800 12448 22018 12576
rect 880 12168 21920 12448
rect 800 12040 22018 12168
rect 880 11488 21920 12040
rect 800 11360 22018 11488
rect 880 11080 21920 11360
rect 800 10952 22018 11080
rect 880 10672 21920 10952
rect 800 10544 22018 10672
rect 880 10264 21920 10544
rect 800 10136 22018 10264
rect 880 9856 21920 10136
rect 800 9728 22018 9856
rect 880 9448 21920 9728
rect 800 9320 22018 9448
rect 880 9040 21920 9320
rect 800 8912 22018 9040
rect 880 8632 21920 8912
rect 800 8504 22018 8632
rect 880 8224 21920 8504
rect 800 8096 22018 8224
rect 880 7544 21920 8096
rect 800 7416 22018 7544
rect 880 7136 21920 7416
rect 800 7008 22018 7136
rect 880 6728 21920 7008
rect 800 6600 22018 6728
rect 880 6320 21920 6600
rect 800 6192 22018 6320
rect 880 5912 21920 6192
rect 800 5784 22018 5912
rect 880 5504 21920 5784
rect 800 5376 22018 5504
rect 880 5096 21920 5376
rect 800 4968 22018 5096
rect 880 4688 21920 4968
rect 800 4560 22018 4688
rect 880 4280 21920 4560
rect 800 4152 22018 4280
rect 880 3600 21920 4152
rect 800 3472 22018 3600
rect 880 3192 21920 3472
rect 800 3064 22018 3192
rect 880 2784 21920 3064
rect 800 2656 22018 2784
rect 880 2376 21920 2656
rect 800 2248 22018 2376
rect 880 1968 21920 2248
rect 800 1840 22018 1968
rect 880 1560 21920 1840
rect 800 1432 22018 1560
rect 880 1152 21920 1432
rect 800 1024 22018 1152
rect 880 744 21920 1024
rect 800 616 22018 744
rect 880 171 21920 616
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 2451 2048 4296 20176
rect 4776 2048 7728 20176
rect 8208 2048 20181 20176
rect 2451 851 20181 2048
<< labels >>
rlabel metal2 s 18418 22000 18474 22800 6 Test_en_N_out
port 1 nsew default output
rlabel metal2 s 18878 0 18934 800 6 Test_en_S_in
port 2 nsew default input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 3 nsew default input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 4 nsew default input
rlabel metal2 s 938 0 994 800 6 bottom_left_grid_pin_44_
port 5 nsew default input
rlabel metal2 s 1306 0 1362 800 6 bottom_left_grid_pin_45_
port 6 nsew default input
rlabel metal2 s 1674 0 1730 800 6 bottom_left_grid_pin_46_
port 7 nsew default input
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_47_
port 8 nsew default input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_48_
port 9 nsew default input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_49_
port 10 nsew default input
rlabel metal2 s 3146 0 3202 800 6 ccff_head
port 11 nsew default input
rlabel metal2 s 3514 0 3570 800 6 ccff_tail
port 12 nsew default output
rlabel metal3 s 0 3272 800 3392 6 chanx_left_in[0]
port 13 nsew default input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[10]
port 14 nsew default input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[11]
port 15 nsew default input
rlabel metal3 s 0 7896 800 8016 6 chanx_left_in[12]
port 16 nsew default input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[13]
port 17 nsew default input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[14]
port 18 nsew default input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[15]
port 19 nsew default input
rlabel metal3 s 0 9528 800 9648 6 chanx_left_in[16]
port 20 nsew default input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[17]
port 21 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[18]
port 22 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[19]
port 23 nsew default input
rlabel metal3 s 0 3680 800 3800 6 chanx_left_in[1]
port 24 nsew default input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[2]
port 25 nsew default input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[3]
port 26 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[4]
port 27 nsew default input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[5]
port 28 nsew default input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[6]
port 29 nsew default input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[7]
port 30 nsew default input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[8]
port 31 nsew default input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[9]
port 32 nsew default input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_out[0]
port 33 nsew default output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[10]
port 34 nsew default output
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[11]
port 35 nsew default output
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[12]
port 36 nsew default output
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[13]
port 37 nsew default output
rlabel metal3 s 0 16600 800 16720 6 chanx_left_out[14]
port 38 nsew default output
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[15]
port 39 nsew default output
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[16]
port 40 nsew default output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[17]
port 41 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[18]
port 42 nsew default output
rlabel metal3 s 0 18640 800 18760 6 chanx_left_out[19]
port 43 nsew default output
rlabel metal3 s 0 11568 800 11688 6 chanx_left_out[1]
port 44 nsew default output
rlabel metal3 s 0 11840 800 11960 6 chanx_left_out[2]
port 45 nsew default output
rlabel metal3 s 0 12248 800 12368 6 chanx_left_out[3]
port 46 nsew default output
rlabel metal3 s 0 12656 800 12776 6 chanx_left_out[4]
port 47 nsew default output
rlabel metal3 s 0 13064 800 13184 6 chanx_left_out[5]
port 48 nsew default output
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[6]
port 49 nsew default output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[7]
port 50 nsew default output
rlabel metal3 s 0 14288 800 14408 6 chanx_left_out[8]
port 51 nsew default output
rlabel metal3 s 0 14696 800 14816 6 chanx_left_out[9]
port 52 nsew default output
rlabel metal3 s 22000 3272 22800 3392 6 chanx_right_in[0]
port 53 nsew default input
rlabel metal3 s 22000 7216 22800 7336 6 chanx_right_in[10]
port 54 nsew default input
rlabel metal3 s 22000 7624 22800 7744 6 chanx_right_in[11]
port 55 nsew default input
rlabel metal3 s 22000 7896 22800 8016 6 chanx_right_in[12]
port 56 nsew default input
rlabel metal3 s 22000 8304 22800 8424 6 chanx_right_in[13]
port 57 nsew default input
rlabel metal3 s 22000 8712 22800 8832 6 chanx_right_in[14]
port 58 nsew default input
rlabel metal3 s 22000 9120 22800 9240 6 chanx_right_in[15]
port 59 nsew default input
rlabel metal3 s 22000 9528 22800 9648 6 chanx_right_in[16]
port 60 nsew default input
rlabel metal3 s 22000 9936 22800 10056 6 chanx_right_in[17]
port 61 nsew default input
rlabel metal3 s 22000 10344 22800 10464 6 chanx_right_in[18]
port 62 nsew default input
rlabel metal3 s 22000 10752 22800 10872 6 chanx_right_in[19]
port 63 nsew default input
rlabel metal3 s 22000 3680 22800 3800 6 chanx_right_in[1]
port 64 nsew default input
rlabel metal3 s 22000 3952 22800 4072 6 chanx_right_in[2]
port 65 nsew default input
rlabel metal3 s 22000 4360 22800 4480 6 chanx_right_in[3]
port 66 nsew default input
rlabel metal3 s 22000 4768 22800 4888 6 chanx_right_in[4]
port 67 nsew default input
rlabel metal3 s 22000 5176 22800 5296 6 chanx_right_in[5]
port 68 nsew default input
rlabel metal3 s 22000 5584 22800 5704 6 chanx_right_in[6]
port 69 nsew default input
rlabel metal3 s 22000 5992 22800 6112 6 chanx_right_in[7]
port 70 nsew default input
rlabel metal3 s 22000 6400 22800 6520 6 chanx_right_in[8]
port 71 nsew default input
rlabel metal3 s 22000 6808 22800 6928 6 chanx_right_in[9]
port 72 nsew default input
rlabel metal3 s 22000 11160 22800 11280 6 chanx_right_out[0]
port 73 nsew default output
rlabel metal3 s 22000 15104 22800 15224 6 chanx_right_out[10]
port 74 nsew default output
rlabel metal3 s 22000 15376 22800 15496 6 chanx_right_out[11]
port 75 nsew default output
rlabel metal3 s 22000 15784 22800 15904 6 chanx_right_out[12]
port 76 nsew default output
rlabel metal3 s 22000 16192 22800 16312 6 chanx_right_out[13]
port 77 nsew default output
rlabel metal3 s 22000 16600 22800 16720 6 chanx_right_out[14]
port 78 nsew default output
rlabel metal3 s 22000 17008 22800 17128 6 chanx_right_out[15]
port 79 nsew default output
rlabel metal3 s 22000 17416 22800 17536 6 chanx_right_out[16]
port 80 nsew default output
rlabel metal3 s 22000 17824 22800 17944 6 chanx_right_out[17]
port 81 nsew default output
rlabel metal3 s 22000 18232 22800 18352 6 chanx_right_out[18]
port 82 nsew default output
rlabel metal3 s 22000 18640 22800 18760 6 chanx_right_out[19]
port 83 nsew default output
rlabel metal3 s 22000 11568 22800 11688 6 chanx_right_out[1]
port 84 nsew default output
rlabel metal3 s 22000 11840 22800 11960 6 chanx_right_out[2]
port 85 nsew default output
rlabel metal3 s 22000 12248 22800 12368 6 chanx_right_out[3]
port 86 nsew default output
rlabel metal3 s 22000 12656 22800 12776 6 chanx_right_out[4]
port 87 nsew default output
rlabel metal3 s 22000 13064 22800 13184 6 chanx_right_out[5]
port 88 nsew default output
rlabel metal3 s 22000 13472 22800 13592 6 chanx_right_out[6]
port 89 nsew default output
rlabel metal3 s 22000 13880 22800 14000 6 chanx_right_out[7]
port 90 nsew default output
rlabel metal3 s 22000 14288 22800 14408 6 chanx_right_out[8]
port 91 nsew default output
rlabel metal3 s 22000 14696 22800 14816 6 chanx_right_out[9]
port 92 nsew default output
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 93 nsew default input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[10]
port 94 nsew default input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[11]
port 95 nsew default input
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_in[12]
port 96 nsew default input
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[13]
port 97 nsew default input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[14]
port 98 nsew default input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[15]
port 99 nsew default input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[16]
port 100 nsew default input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[17]
port 101 nsew default input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[18]
port 102 nsew default input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[19]
port 103 nsew default input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[1]
port 104 nsew default input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[2]
port 105 nsew default input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[3]
port 106 nsew default input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[4]
port 107 nsew default input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[5]
port 108 nsew default input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[6]
port 109 nsew default input
rlabel metal2 s 6550 0 6606 800 6 chany_bottom_in[7]
port 110 nsew default input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[8]
port 111 nsew default input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[9]
port 112 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_out[0]
port 113 nsew default output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[10]
port 114 nsew default output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[11]
port 115 nsew default output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[12]
port 116 nsew default output
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_out[13]
port 117 nsew default output
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[14]
port 118 nsew default output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[15]
port 119 nsew default output
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[16]
port 120 nsew default output
rlabel metal2 s 17774 0 17830 800 6 chany_bottom_out[17]
port 121 nsew default output
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[18]
port 122 nsew default output
rlabel metal2 s 18510 0 18566 800 6 chany_bottom_out[19]
port 123 nsew default output
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_out[1]
port 124 nsew default output
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[2]
port 125 nsew default output
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[3]
port 126 nsew default output
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_out[4]
port 127 nsew default output
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[5]
port 128 nsew default output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[6]
port 129 nsew default output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[7]
port 130 nsew default output
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[8]
port 131 nsew default output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[9]
port 132 nsew default output
rlabel metal2 s 3238 22000 3294 22800 6 chany_top_in[0]
port 133 nsew default input
rlabel metal2 s 7010 22000 7066 22800 6 chany_top_in[10]
port 134 nsew default input
rlabel metal2 s 7378 22000 7434 22800 6 chany_top_in[11]
port 135 nsew default input
rlabel metal2 s 7746 22000 7802 22800 6 chany_top_in[12]
port 136 nsew default input
rlabel metal2 s 8114 22000 8170 22800 6 chany_top_in[13]
port 137 nsew default input
rlabel metal2 s 8482 22000 8538 22800 6 chany_top_in[14]
port 138 nsew default input
rlabel metal2 s 8942 22000 8998 22800 6 chany_top_in[15]
port 139 nsew default input
rlabel metal2 s 9310 22000 9366 22800 6 chany_top_in[16]
port 140 nsew default input
rlabel metal2 s 9678 22000 9734 22800 6 chany_top_in[17]
port 141 nsew default input
rlabel metal2 s 10046 22000 10102 22800 6 chany_top_in[18]
port 142 nsew default input
rlabel metal2 s 10414 22000 10470 22800 6 chany_top_in[19]
port 143 nsew default input
rlabel metal2 s 3606 22000 3662 22800 6 chany_top_in[1]
port 144 nsew default input
rlabel metal2 s 3974 22000 4030 22800 6 chany_top_in[2]
port 145 nsew default input
rlabel metal2 s 4342 22000 4398 22800 6 chany_top_in[3]
port 146 nsew default input
rlabel metal2 s 4710 22000 4766 22800 6 chany_top_in[4]
port 147 nsew default input
rlabel metal2 s 5078 22000 5134 22800 6 chany_top_in[5]
port 148 nsew default input
rlabel metal2 s 5446 22000 5502 22800 6 chany_top_in[6]
port 149 nsew default input
rlabel metal2 s 5906 22000 5962 22800 6 chany_top_in[7]
port 150 nsew default input
rlabel metal2 s 6274 22000 6330 22800 6 chany_top_in[8]
port 151 nsew default input
rlabel metal2 s 6642 22000 6698 22800 6 chany_top_in[9]
port 152 nsew default input
rlabel metal2 s 10782 22000 10838 22800 6 chany_top_out[0]
port 153 nsew default output
rlabel metal2 s 14646 22000 14702 22800 6 chany_top_out[10]
port 154 nsew default output
rlabel metal2 s 15014 22000 15070 22800 6 chany_top_out[11]
port 155 nsew default output
rlabel metal2 s 15382 22000 15438 22800 6 chany_top_out[12]
port 156 nsew default output
rlabel metal2 s 15750 22000 15806 22800 6 chany_top_out[13]
port 157 nsew default output
rlabel metal2 s 16118 22000 16174 22800 6 chany_top_out[14]
port 158 nsew default output
rlabel metal2 s 16486 22000 16542 22800 6 chany_top_out[15]
port 159 nsew default output
rlabel metal2 s 16854 22000 16910 22800 6 chany_top_out[16]
port 160 nsew default output
rlabel metal2 s 17314 22000 17370 22800 6 chany_top_out[17]
port 161 nsew default output
rlabel metal2 s 17682 22000 17738 22800 6 chany_top_out[18]
port 162 nsew default output
rlabel metal2 s 18050 22000 18106 22800 6 chany_top_out[19]
port 163 nsew default output
rlabel metal2 s 11150 22000 11206 22800 6 chany_top_out[1]
port 164 nsew default output
rlabel metal2 s 11610 22000 11666 22800 6 chany_top_out[2]
port 165 nsew default output
rlabel metal2 s 11978 22000 12034 22800 6 chany_top_out[3]
port 166 nsew default output
rlabel metal2 s 12346 22000 12402 22800 6 chany_top_out[4]
port 167 nsew default output
rlabel metal2 s 12714 22000 12770 22800 6 chany_top_out[5]
port 168 nsew default output
rlabel metal2 s 13082 22000 13138 22800 6 chany_top_out[6]
port 169 nsew default output
rlabel metal2 s 13450 22000 13506 22800 6 chany_top_out[7]
port 170 nsew default output
rlabel metal2 s 13818 22000 13874 22800 6 chany_top_out[8]
port 171 nsew default output
rlabel metal2 s 14186 22000 14242 22800 6 chany_top_out[9]
port 172 nsew default output
rlabel metal3 s 22000 20544 22800 20664 6 clk_1_E_out
port 173 nsew default output
rlabel metal2 s 18786 22000 18842 22800 6 clk_1_N_in
port 174 nsew default input
rlabel metal2 s 19246 0 19302 800 6 clk_1_S_in
port 175 nsew default input
rlabel metal3 s 0 19048 800 19168 6 clk_1_W_out
port 176 nsew default output
rlabel metal3 s 22000 19048 22800 19168 6 clk_2_E_in
port 177 nsew default input
rlabel metal3 s 22000 20952 22800 21072 6 clk_2_E_out
port 178 nsew default output
rlabel metal2 s 19154 22000 19210 22800 6 clk_2_N_in
port 179 nsew default input
rlabel metal2 s 21454 22000 21510 22800 6 clk_2_N_out
port 180 nsew default output
rlabel metal2 s 19614 0 19670 800 6 clk_2_S_in
port 181 nsew default input
rlabel metal2 s 20350 0 20406 800 6 clk_2_S_out
port 182 nsew default output
rlabel metal3 s 0 21360 800 21480 6 clk_2_W_in
port 183 nsew default input
rlabel metal3 s 0 19320 800 19440 6 clk_2_W_out
port 184 nsew default output
rlabel metal3 s 22000 19320 22800 19440 6 clk_3_E_in
port 185 nsew default input
rlabel metal3 s 22000 21360 22800 21480 6 clk_3_E_out
port 186 nsew default output
rlabel metal2 s 19522 22000 19578 22800 6 clk_3_N_in
port 187 nsew default input
rlabel metal2 s 21822 22000 21878 22800 6 clk_3_N_out
port 188 nsew default output
rlabel metal2 s 19982 0 20038 800 6 clk_3_S_in
port 189 nsew default input
rlabel metal2 s 20718 0 20774 800 6 clk_3_S_out
port 190 nsew default output
rlabel metal3 s 0 21768 800 21888 6 clk_3_W_in
port 191 nsew default input
rlabel metal3 s 0 19728 800 19848 6 clk_3_W_out
port 192 nsew default output
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 193 nsew default input
rlabel metal3 s 0 416 800 536 6 left_bottom_grid_pin_35_
port 194 nsew default input
rlabel metal3 s 0 824 800 944 6 left_bottom_grid_pin_36_
port 195 nsew default input
rlabel metal3 s 0 1232 800 1352 6 left_bottom_grid_pin_37_
port 196 nsew default input
rlabel metal3 s 0 1640 800 1760 6 left_bottom_grid_pin_38_
port 197 nsew default input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_39_
port 198 nsew default input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_40_
port 199 nsew default input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_41_
port 200 nsew default input
rlabel metal2 s 19890 22000 19946 22800 6 prog_clk_0_N_in
port 201 nsew default input
rlabel metal3 s 22000 21768 22800 21888 6 prog_clk_1_E_out
port 202 nsew default output
rlabel metal2 s 20350 22000 20406 22800 6 prog_clk_1_N_in
port 203 nsew default input
rlabel metal2 s 21086 0 21142 800 6 prog_clk_1_S_in
port 204 nsew default input
rlabel metal3 s 0 20136 800 20256 6 prog_clk_1_W_out
port 205 nsew default output
rlabel metal3 s 22000 19728 22800 19848 6 prog_clk_2_E_in
port 206 nsew default input
rlabel metal3 s 22000 22176 22800 22296 6 prog_clk_2_E_out
port 207 nsew default output
rlabel metal2 s 20718 22000 20774 22800 6 prog_clk_2_N_in
port 208 nsew default input
rlabel metal2 s 22190 22000 22246 22800 6 prog_clk_2_N_out
port 209 nsew default output
rlabel metal2 s 21454 0 21510 800 6 prog_clk_2_S_in
port 210 nsew default input
rlabel metal2 s 22190 0 22246 800 6 prog_clk_2_S_out
port 211 nsew default output
rlabel metal3 s 0 22176 800 22296 6 prog_clk_2_W_in
port 212 nsew default input
rlabel metal3 s 0 20544 800 20664 6 prog_clk_2_W_out
port 213 nsew default output
rlabel metal3 s 22000 20136 22800 20256 6 prog_clk_3_E_in
port 214 nsew default input
rlabel metal3 s 22000 22584 22800 22704 6 prog_clk_3_E_out
port 215 nsew default output
rlabel metal2 s 21086 22000 21142 22800 6 prog_clk_3_N_in
port 216 nsew default input
rlabel metal2 s 22558 22000 22614 22800 6 prog_clk_3_N_out
port 217 nsew default output
rlabel metal2 s 21822 0 21878 800 6 prog_clk_3_S_in
port 218 nsew default input
rlabel metal2 s 22558 0 22614 800 6 prog_clk_3_S_out
port 219 nsew default output
rlabel metal3 s 0 22584 800 22704 6 prog_clk_3_W_in
port 220 nsew default input
rlabel metal3 s 0 20952 800 21072 6 prog_clk_3_W_out
port 221 nsew default output
rlabel metal3 s 22000 144 22800 264 6 right_bottom_grid_pin_34_
port 222 nsew default input
rlabel metal3 s 22000 416 22800 536 6 right_bottom_grid_pin_35_
port 223 nsew default input
rlabel metal3 s 22000 824 22800 944 6 right_bottom_grid_pin_36_
port 224 nsew default input
rlabel metal3 s 22000 1232 22800 1352 6 right_bottom_grid_pin_37_
port 225 nsew default input
rlabel metal3 s 22000 1640 22800 1760 6 right_bottom_grid_pin_38_
port 226 nsew default input
rlabel metal3 s 22000 2048 22800 2168 6 right_bottom_grid_pin_39_
port 227 nsew default input
rlabel metal3 s 22000 2456 22800 2576 6 right_bottom_grid_pin_40_
port 228 nsew default input
rlabel metal3 s 22000 2864 22800 2984 6 right_bottom_grid_pin_41_
port 229 nsew default input
rlabel metal2 s 202 22000 258 22800 6 top_left_grid_pin_42_
port 230 nsew default input
rlabel metal2 s 570 22000 626 22800 6 top_left_grid_pin_43_
port 231 nsew default input
rlabel metal2 s 938 22000 994 22800 6 top_left_grid_pin_44_
port 232 nsew default input
rlabel metal2 s 1306 22000 1362 22800 6 top_left_grid_pin_45_
port 233 nsew default input
rlabel metal2 s 1674 22000 1730 22800 6 top_left_grid_pin_46_
port 234 nsew default input
rlabel metal2 s 2042 22000 2098 22800 6 top_left_grid_pin_47_
port 235 nsew default input
rlabel metal2 s 2410 22000 2466 22800 6 top_left_grid_pin_48_
port 236 nsew default input
rlabel metal2 s 2778 22000 2834 22800 6 top_left_grid_pin_49_
port 237 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 238 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 239 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
