magic
tech sky130A
magscale 1 2
timestamp 1608155778
<< obsli1 >>
rect 1104 2015 21775 20001
<< obsm1 >>
rect 290 1156 22526 20032
<< metal2 >>
rect 294 21856 350 22656
rect 846 21856 902 22656
rect 1398 21856 1454 22656
rect 1950 21856 2006 22656
rect 2502 21856 2558 22656
rect 3054 21856 3110 22656
rect 3606 21856 3662 22656
rect 4158 21856 4214 22656
rect 4710 21856 4766 22656
rect 5262 21856 5318 22656
rect 5814 21856 5870 22656
rect 6366 21856 6422 22656
rect 6918 21856 6974 22656
rect 7470 21856 7526 22656
rect 8022 21856 8078 22656
rect 8574 21856 8630 22656
rect 9126 21856 9182 22656
rect 9678 21856 9734 22656
rect 10230 21856 10286 22656
rect 10782 21856 10838 22656
rect 11334 21856 11390 22656
rect 11978 21856 12034 22656
rect 12530 21856 12586 22656
rect 13082 21856 13138 22656
rect 13634 21856 13690 22656
rect 14186 21856 14242 22656
rect 14738 21856 14794 22656
rect 15290 21856 15346 22656
rect 15842 21856 15898 22656
rect 16394 21856 16450 22656
rect 16946 21856 17002 22656
rect 17498 21856 17554 22656
rect 18050 21856 18106 22656
rect 18602 21856 18658 22656
rect 19154 21856 19210 22656
rect 19706 21856 19762 22656
rect 20258 21856 20314 22656
rect 20810 21856 20866 22656
rect 21362 21856 21418 22656
rect 21914 21856 21970 22656
rect 22466 21856 22522 22656
<< obsm2 >>
rect 406 21800 790 22401
rect 958 21800 1342 22401
rect 1510 21800 1894 22401
rect 2062 21800 2446 22401
rect 2614 21800 2998 22401
rect 3166 21800 3550 22401
rect 3718 21800 4102 22401
rect 4270 21800 4654 22401
rect 4822 21800 5206 22401
rect 5374 21800 5758 22401
rect 5926 21800 6310 22401
rect 6478 21800 6862 22401
rect 7030 21800 7414 22401
rect 7582 21800 7966 22401
rect 8134 21800 8518 22401
rect 8686 21800 9070 22401
rect 9238 21800 9622 22401
rect 9790 21800 10174 22401
rect 10342 21800 10726 22401
rect 10894 21800 11278 22401
rect 11446 21800 11922 22401
rect 12090 21800 12474 22401
rect 12642 21800 13026 22401
rect 13194 21800 13578 22401
rect 13746 21800 14130 22401
rect 14298 21800 14682 22401
rect 14850 21800 15234 22401
rect 15402 21800 15786 22401
rect 15954 21800 16338 22401
rect 16506 21800 16890 22401
rect 17058 21800 17442 22401
rect 17610 21800 17994 22401
rect 18162 21800 18546 22401
rect 18714 21800 19098 22401
rect 19266 21800 19650 22401
rect 19818 21800 20202 22401
rect 20370 21800 20754 22401
rect 20922 21800 21306 22401
rect 21474 21800 21858 22401
rect 22026 21800 22410 22401
rect 296 23 22520 21800
<< metal3 >>
rect 22000 22304 22800 22424
rect 22000 21896 22800 22016
rect 22000 21352 22800 21472
rect 22000 20944 22800 21064
rect 22000 20536 22800 20656
rect 22000 19992 22800 20112
rect 22000 19584 22800 19704
rect 22000 19176 22800 19296
rect 22000 18632 22800 18752
rect 22000 18224 22800 18344
rect 22000 17816 22800 17936
rect 22000 17272 22800 17392
rect 0 17000 800 17120
rect 22000 16864 22800 16984
rect 22000 16320 22800 16440
rect 22000 15912 22800 16032
rect 22000 15504 22800 15624
rect 22000 14960 22800 15080
rect 22000 14552 22800 14672
rect 22000 14144 22800 14264
rect 22000 13600 22800 13720
rect 22000 13192 22800 13312
rect 22000 12784 22800 12904
rect 22000 12240 22800 12360
rect 22000 11832 22800 11952
rect 22000 11424 22800 11544
rect 22000 10880 22800 11000
rect 22000 10472 22800 10592
rect 22000 9928 22800 10048
rect 22000 9520 22800 9640
rect 22000 9112 22800 9232
rect 22000 8568 22800 8688
rect 22000 8160 22800 8280
rect 22000 7752 22800 7872
rect 22000 7208 22800 7328
rect 22000 6800 22800 6920
rect 22000 6392 22800 6512
rect 22000 5848 22800 5968
rect 0 5576 800 5696
rect 22000 5440 22800 5560
rect 22000 4896 22800 5016
rect 22000 4488 22800 4608
rect 22000 4080 22800 4200
rect 22000 3536 22800 3656
rect 22000 3128 22800 3248
rect 22000 2720 22800 2840
rect 22000 2176 22800 2296
rect 22000 1768 22800 1888
rect 22000 1360 22800 1480
rect 22000 816 22800 936
rect 22000 408 22800 528
rect 22000 0 22800 120
<< obsm3 >>
rect 800 22224 21920 22397
rect 800 22096 22000 22224
rect 800 21816 21920 22096
rect 800 21552 22000 21816
rect 800 21272 21920 21552
rect 800 21144 22000 21272
rect 800 20864 21920 21144
rect 800 20736 22000 20864
rect 800 20456 21920 20736
rect 800 20192 22000 20456
rect 800 19912 21920 20192
rect 800 19784 22000 19912
rect 800 19504 21920 19784
rect 800 19376 22000 19504
rect 800 19096 21920 19376
rect 800 18832 22000 19096
rect 800 18552 21920 18832
rect 800 18424 22000 18552
rect 800 18144 21920 18424
rect 800 18016 22000 18144
rect 800 17736 21920 18016
rect 800 17472 22000 17736
rect 800 17200 21920 17472
rect 880 17192 21920 17200
rect 880 17064 22000 17192
rect 880 16920 21920 17064
rect 800 16784 21920 16920
rect 800 16520 22000 16784
rect 800 16240 21920 16520
rect 800 16112 22000 16240
rect 800 15832 21920 16112
rect 800 15704 22000 15832
rect 800 15424 21920 15704
rect 800 15160 22000 15424
rect 800 14880 21920 15160
rect 800 14752 22000 14880
rect 800 14472 21920 14752
rect 800 14344 22000 14472
rect 800 14064 21920 14344
rect 800 13800 22000 14064
rect 800 13520 21920 13800
rect 800 13392 22000 13520
rect 800 13112 21920 13392
rect 800 12984 22000 13112
rect 800 12704 21920 12984
rect 800 12440 22000 12704
rect 800 12160 21920 12440
rect 800 12032 22000 12160
rect 800 11752 21920 12032
rect 800 11624 22000 11752
rect 800 11344 21920 11624
rect 800 11080 22000 11344
rect 800 10800 21920 11080
rect 800 10672 22000 10800
rect 800 10392 21920 10672
rect 800 10128 22000 10392
rect 800 9848 21920 10128
rect 800 9720 22000 9848
rect 800 9440 21920 9720
rect 800 9312 22000 9440
rect 800 9032 21920 9312
rect 800 8768 22000 9032
rect 800 8488 21920 8768
rect 800 8360 22000 8488
rect 800 8080 21920 8360
rect 800 7952 22000 8080
rect 800 7672 21920 7952
rect 800 7408 22000 7672
rect 800 7128 21920 7408
rect 800 7000 22000 7128
rect 800 6720 21920 7000
rect 800 6592 22000 6720
rect 800 6312 21920 6592
rect 800 6048 22000 6312
rect 800 5776 21920 6048
rect 880 5768 21920 5776
rect 880 5640 22000 5768
rect 880 5496 21920 5640
rect 800 5360 21920 5496
rect 800 5096 22000 5360
rect 800 4816 21920 5096
rect 800 4688 22000 4816
rect 800 4408 21920 4688
rect 800 4280 22000 4408
rect 800 4000 21920 4280
rect 800 3736 22000 4000
rect 800 3456 21920 3736
rect 800 3328 22000 3456
rect 800 3048 21920 3328
rect 800 2920 22000 3048
rect 800 2640 21920 2920
rect 800 2376 22000 2640
rect 800 2096 21920 2376
rect 800 1968 22000 2096
rect 800 1688 21920 1968
rect 800 1560 22000 1688
rect 800 1280 21920 1560
rect 800 1016 22000 1280
rect 800 736 21920 1016
rect 800 608 22000 736
rect 800 328 21920 608
rect 800 200 22000 328
rect 800 27 21920 200
<< metal4 >>
rect 4376 1984 4696 20032
rect 7808 1984 8128 20032
<< obsm4 >>
rect 11240 1984 18424 20032
<< labels >>
rlabel metal3 s 0 5576 800 5696 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 17000 800 17120 6 ccff_tail
port 2 nsew default output
rlabel metal3 s 22000 4080 22800 4200 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22000 8568 22800 8688 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22000 9112 22800 9232 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22000 9520 22800 9640 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22000 9928 22800 10048 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22000 10472 22800 10592 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22000 10880 22800 11000 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22000 11424 22800 11544 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22000 11832 22800 11952 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22000 12240 22800 12360 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22000 12784 22800 12904 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22000 4488 22800 4608 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22000 4896 22800 5016 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22000 5440 22800 5560 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22000 5848 22800 5968 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22000 6392 22800 6512 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22000 6800 22800 6920 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22000 7208 22800 7328 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22000 7752 22800 7872 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22000 8160 22800 8280 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22000 13192 22800 13312 6 chanx_right_out[0]
port 23 nsew default output
rlabel metal3 s 22000 17816 22800 17936 6 chanx_right_out[10]
port 24 nsew default output
rlabel metal3 s 22000 18224 22800 18344 6 chanx_right_out[11]
port 25 nsew default output
rlabel metal3 s 22000 18632 22800 18752 6 chanx_right_out[12]
port 26 nsew default output
rlabel metal3 s 22000 19176 22800 19296 6 chanx_right_out[13]
port 27 nsew default output
rlabel metal3 s 22000 19584 22800 19704 6 chanx_right_out[14]
port 28 nsew default output
rlabel metal3 s 22000 19992 22800 20112 6 chanx_right_out[15]
port 29 nsew default output
rlabel metal3 s 22000 20536 22800 20656 6 chanx_right_out[16]
port 30 nsew default output
rlabel metal3 s 22000 20944 22800 21064 6 chanx_right_out[17]
port 31 nsew default output
rlabel metal3 s 22000 21352 22800 21472 6 chanx_right_out[18]
port 32 nsew default output
rlabel metal3 s 22000 21896 22800 22016 6 chanx_right_out[19]
port 33 nsew default output
rlabel metal3 s 22000 13600 22800 13720 6 chanx_right_out[1]
port 34 nsew default output
rlabel metal3 s 22000 14144 22800 14264 6 chanx_right_out[2]
port 35 nsew default output
rlabel metal3 s 22000 14552 22800 14672 6 chanx_right_out[3]
port 36 nsew default output
rlabel metal3 s 22000 14960 22800 15080 6 chanx_right_out[4]
port 37 nsew default output
rlabel metal3 s 22000 15504 22800 15624 6 chanx_right_out[5]
port 38 nsew default output
rlabel metal3 s 22000 15912 22800 16032 6 chanx_right_out[6]
port 39 nsew default output
rlabel metal3 s 22000 16320 22800 16440 6 chanx_right_out[7]
port 40 nsew default output
rlabel metal3 s 22000 16864 22800 16984 6 chanx_right_out[8]
port 41 nsew default output
rlabel metal3 s 22000 17272 22800 17392 6 chanx_right_out[9]
port 42 nsew default output
rlabel metal2 s 846 21856 902 22656 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 6366 21856 6422 22656 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 6918 21856 6974 22656 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 7470 21856 7526 22656 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 8022 21856 8078 22656 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 8574 21856 8630 22656 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 9126 21856 9182 22656 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 9678 21856 9734 22656 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 10230 21856 10286 22656 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 10782 21856 10838 22656 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 11334 21856 11390 22656 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 1398 21856 1454 22656 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 1950 21856 2006 22656 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 2502 21856 2558 22656 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 3054 21856 3110 22656 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 3606 21856 3662 22656 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 4158 21856 4214 22656 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 4710 21856 4766 22656 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 5262 21856 5318 22656 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 5814 21856 5870 22656 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 11978 21856 12034 22656 6 chany_top_out[0]
port 63 nsew default output
rlabel metal2 s 17498 21856 17554 22656 6 chany_top_out[10]
port 64 nsew default output
rlabel metal2 s 18050 21856 18106 22656 6 chany_top_out[11]
port 65 nsew default output
rlabel metal2 s 18602 21856 18658 22656 6 chany_top_out[12]
port 66 nsew default output
rlabel metal2 s 19154 21856 19210 22656 6 chany_top_out[13]
port 67 nsew default output
rlabel metal2 s 19706 21856 19762 22656 6 chany_top_out[14]
port 68 nsew default output
rlabel metal2 s 20258 21856 20314 22656 6 chany_top_out[15]
port 69 nsew default output
rlabel metal2 s 20810 21856 20866 22656 6 chany_top_out[16]
port 70 nsew default output
rlabel metal2 s 21362 21856 21418 22656 6 chany_top_out[17]
port 71 nsew default output
rlabel metal2 s 21914 21856 21970 22656 6 chany_top_out[18]
port 72 nsew default output
rlabel metal2 s 22466 21856 22522 22656 6 chany_top_out[19]
port 73 nsew default output
rlabel metal2 s 12530 21856 12586 22656 6 chany_top_out[1]
port 74 nsew default output
rlabel metal2 s 13082 21856 13138 22656 6 chany_top_out[2]
port 75 nsew default output
rlabel metal2 s 13634 21856 13690 22656 6 chany_top_out[3]
port 76 nsew default output
rlabel metal2 s 14186 21856 14242 22656 6 chany_top_out[4]
port 77 nsew default output
rlabel metal2 s 14738 21856 14794 22656 6 chany_top_out[5]
port 78 nsew default output
rlabel metal2 s 15290 21856 15346 22656 6 chany_top_out[6]
port 79 nsew default output
rlabel metal2 s 15842 21856 15898 22656 6 chany_top_out[7]
port 80 nsew default output
rlabel metal2 s 16394 21856 16450 22656 6 chany_top_out[8]
port 81 nsew default output
rlabel metal2 s 16946 21856 17002 22656 6 chany_top_out[9]
port 82 nsew default output
rlabel metal3 s 22000 22304 22800 22424 6 prog_clk_0_E_in
port 83 nsew default input
rlabel metal3 s 22000 2176 22800 2296 6 right_bottom_grid_pin_11_
port 84 nsew default input
rlabel metal3 s 22000 2720 22800 2840 6 right_bottom_grid_pin_13_
port 85 nsew default input
rlabel metal3 s 22000 3128 22800 3248 6 right_bottom_grid_pin_15_
port 86 nsew default input
rlabel metal3 s 22000 3536 22800 3656 6 right_bottom_grid_pin_17_
port 87 nsew default input
rlabel metal3 s 22000 0 22800 120 6 right_bottom_grid_pin_1_
port 88 nsew default input
rlabel metal3 s 22000 408 22800 528 6 right_bottom_grid_pin_3_
port 89 nsew default input
rlabel metal3 s 22000 816 22800 936 6 right_bottom_grid_pin_5_
port 90 nsew default input
rlabel metal3 s 22000 1360 22800 1480 6 right_bottom_grid_pin_7_
port 91 nsew default input
rlabel metal3 s 22000 1768 22800 1888 6 right_bottom_grid_pin_9_
port 92 nsew default input
rlabel metal2 s 294 21856 350 22656 6 top_left_grid_pin_1_
port 93 nsew default input
rlabel metal4 s 4376 1984 4696 20032 6 VPWR
port 94 nsew power input
rlabel metal4 s 7808 1984 8128 20032 6 VGND
port 95 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22656
string LEFview TRUE
<< end >>
