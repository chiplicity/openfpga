magic
tech sky130A
magscale 1 2
timestamp 1605200686
<< locali >>
rect 10517 10047 10551 10217
<< viali >>
rect 9965 20553 9999 20587
rect 12817 20553 12851 20587
rect 13921 20553 13955 20587
rect 11069 20485 11103 20519
rect 2513 20417 2547 20451
rect 2237 20349 2271 20383
rect 4077 20349 4111 20383
rect 5353 20349 5387 20383
rect 6929 20349 6963 20383
rect 8033 20349 8067 20383
rect 9781 20349 9815 20383
rect 10885 20349 10919 20383
rect 12633 20349 12667 20383
rect 13737 20349 13771 20383
rect 4353 20281 4387 20315
rect 5549 20213 5583 20247
rect 7113 20213 7147 20247
rect 8217 20213 8251 20247
rect 12633 20009 12667 20043
rect 4353 19941 4387 19975
rect 9965 19941 9999 19975
rect 11437 19941 11471 19975
rect 2145 19873 2179 19907
rect 2421 19873 2455 19907
rect 4077 19873 4111 19907
rect 5365 19873 5399 19907
rect 6653 19873 6687 19907
rect 8309 19873 8343 19907
rect 9689 19873 9723 19907
rect 11161 19873 11195 19907
rect 12449 19873 12483 19907
rect 13553 19873 13587 19907
rect 17233 19873 17267 19907
rect 5641 19805 5675 19839
rect 8585 19805 8619 19839
rect 13737 19737 13771 19771
rect 6837 19669 6871 19703
rect 9137 19465 9171 19499
rect 12449 19465 12483 19499
rect 4905 19329 4939 19363
rect 7481 19329 7515 19363
rect 9781 19329 9815 19363
rect 13093 19329 13127 19363
rect 2329 19261 2363 19295
rect 10701 19261 10735 19295
rect 20545 19261 20579 19295
rect 2605 19193 2639 19227
rect 7205 19193 7239 19227
rect 20453 19193 20487 19227
rect 4261 19125 4295 19159
rect 4629 19125 4663 19159
rect 4721 19125 4755 19159
rect 6837 19125 6871 19159
rect 7297 19125 7331 19159
rect 9505 19125 9539 19159
rect 9597 19125 9631 19159
rect 10885 19125 10919 19159
rect 12817 19125 12851 19159
rect 12909 19125 12943 19159
rect 20729 19125 20763 19159
rect 1409 18921 1443 18955
rect 6377 18921 6411 18955
rect 8585 18921 8619 18955
rect 9689 18921 9723 18955
rect 13461 18921 13495 18955
rect 2697 18853 2731 18887
rect 5242 18853 5276 18887
rect 11498 18853 11532 18887
rect 2421 18785 2455 18819
rect 7461 18785 7495 18819
rect 10057 18785 10091 18819
rect 11253 18785 11287 18819
rect 4997 18717 5031 18751
rect 7205 18717 7239 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 10609 18581 10643 18615
rect 12633 18581 12667 18615
rect 5457 18377 5491 18411
rect 11253 18377 11287 18411
rect 2513 18241 2547 18275
rect 12633 18241 12667 18275
rect 2237 18173 2271 18207
rect 4077 18173 4111 18207
rect 7021 18173 7055 18207
rect 9873 18173 9907 18207
rect 12889 18173 12923 18207
rect 4344 18105 4378 18139
rect 7288 18105 7322 18139
rect 10140 18105 10174 18139
rect 8401 18037 8435 18071
rect 14013 18037 14047 18071
rect 4905 17833 4939 17867
rect 7021 17833 7055 17867
rect 7389 17833 7423 17867
rect 8585 17833 8619 17867
rect 11069 17833 11103 17867
rect 12081 17833 12115 17867
rect 13001 17833 13035 17867
rect 6929 17765 6963 17799
rect 2226 17697 2260 17731
rect 5273 17697 5307 17731
rect 5365 17697 5399 17731
rect 7481 17697 7515 17731
rect 9689 17697 9723 17731
rect 9956 17697 9990 17731
rect 11897 17697 11931 17731
rect 2513 17629 2547 17663
rect 4813 17629 4847 17663
rect 5457 17629 5491 17663
rect 7573 17629 7607 17663
rect 5181 17289 5215 17323
rect 9505 17289 9539 17323
rect 12449 17289 12483 17323
rect 11253 17221 11287 17255
rect 8585 17153 8619 17187
rect 10149 17153 10183 17187
rect 13001 17153 13035 17187
rect 2134 17085 2168 17119
rect 3801 17085 3835 17119
rect 6837 17085 6871 17119
rect 11069 17085 11103 17119
rect 12817 17085 12851 17119
rect 2421 17017 2455 17051
rect 4068 17017 4102 17051
rect 8401 17017 8435 17051
rect 9873 17017 9907 17051
rect 7021 16949 7055 16983
rect 7941 16949 7975 16983
rect 8309 16949 8343 16983
rect 9965 16949 9999 16983
rect 12909 16949 12943 16983
rect 13277 16949 13311 16983
rect 2421 16745 2455 16779
rect 11989 16745 12023 16779
rect 5917 16677 5951 16711
rect 12817 16677 12851 16711
rect 1409 16609 1443 16643
rect 2789 16609 2823 16643
rect 4445 16609 4479 16643
rect 4537 16609 4571 16643
rect 5641 16609 5675 16643
rect 7196 16609 7230 16643
rect 10609 16609 10643 16643
rect 10876 16609 10910 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 4721 16541 4755 16575
rect 6929 16541 6963 16575
rect 4077 16473 4111 16507
rect 8309 16405 8343 16439
rect 5733 16201 5767 16235
rect 12449 16201 12483 16235
rect 11161 16133 11195 16167
rect 2513 16065 2547 16099
rect 13001 16065 13035 16099
rect 2237 15997 2271 16031
rect 4353 15997 4387 16031
rect 7389 15997 7423 16031
rect 9781 15997 9815 16031
rect 14013 15997 14047 16031
rect 4620 15929 4654 15963
rect 7656 15929 7690 15963
rect 10048 15929 10082 15963
rect 8769 15861 8803 15895
rect 12817 15861 12851 15895
rect 12909 15861 12943 15895
rect 13277 15861 13311 15895
rect 5457 15657 5491 15691
rect 6285 15657 6319 15691
rect 6653 15657 6687 15691
rect 7849 15657 7883 15691
rect 10057 15657 10091 15691
rect 13001 15657 13035 15691
rect 4344 15589 4378 15623
rect 10425 15589 10459 15623
rect 2237 15521 2271 15555
rect 4077 15521 4111 15555
rect 6193 15521 6227 15555
rect 6745 15521 6779 15555
rect 8217 15521 8251 15555
rect 8309 15521 8343 15555
rect 11888 15521 11922 15555
rect 2513 15453 2547 15487
rect 6837 15453 6871 15487
rect 7757 15453 7791 15487
rect 8401 15453 8435 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 11621 15453 11655 15487
rect 9873 15317 9907 15351
rect 3433 15113 3467 15147
rect 7021 15113 7055 15147
rect 9965 15113 9999 15147
rect 11621 15113 11655 15147
rect 13829 15113 13863 15147
rect 5181 15045 5215 15079
rect 4077 14977 4111 15011
rect 5825 14977 5859 15011
rect 8769 14977 8803 15011
rect 10609 14977 10643 15011
rect 1685 14909 1719 14943
rect 6837 14909 6871 14943
rect 7757 14909 7791 14943
rect 8585 14909 8619 14943
rect 11805 14909 11839 14943
rect 12449 14909 12483 14943
rect 1961 14841 1995 14875
rect 3801 14841 3835 14875
rect 5641 14841 5675 14875
rect 8125 14841 8159 14875
rect 12694 14841 12728 14875
rect 3893 14773 3927 14807
rect 5549 14773 5583 14807
rect 7573 14773 7607 14807
rect 8217 14773 8251 14807
rect 8677 14773 8711 14807
rect 10333 14773 10367 14807
rect 10425 14773 10459 14807
rect 7021 14569 7055 14603
rect 7849 14569 7883 14603
rect 8309 14569 8343 14603
rect 9873 14569 9907 14603
rect 12449 14569 12483 14603
rect 1409 14501 1443 14535
rect 4445 14501 4479 14535
rect 5886 14501 5920 14535
rect 2789 14433 2823 14467
rect 5641 14433 5675 14467
rect 8217 14433 8251 14467
rect 9689 14433 9723 14467
rect 11069 14433 11103 14467
rect 11336 14433 11370 14467
rect 2881 14365 2915 14399
rect 2973 14365 3007 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 8401 14365 8435 14399
rect 2421 14229 2455 14263
rect 4077 14229 4111 14263
rect 4997 14229 5031 14263
rect 5181 14025 5215 14059
rect 9229 14025 9263 14059
rect 10057 14025 10091 14059
rect 1593 13957 1627 13991
rect 2145 13889 2179 13923
rect 3801 13889 3835 13923
rect 5825 13889 5859 13923
rect 10701 13889 10735 13923
rect 2053 13821 2087 13855
rect 3617 13821 3651 13855
rect 4721 13821 4755 13855
rect 5089 13821 5123 13855
rect 5641 13821 5675 13855
rect 7849 13821 7883 13855
rect 8116 13821 8150 13855
rect 9965 13821 9999 13855
rect 12449 13753 12483 13787
rect 1961 13685 1995 13719
rect 3157 13685 3191 13719
rect 3525 13685 3559 13719
rect 4537 13685 4571 13719
rect 5549 13685 5583 13719
rect 6837 13685 6871 13719
rect 10425 13685 10459 13719
rect 10517 13685 10551 13719
rect 2421 13481 2455 13515
rect 2789 13481 2823 13515
rect 4261 13481 4295 13515
rect 6653 13481 6687 13515
rect 7481 13481 7515 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 8493 13481 8527 13515
rect 10333 13481 10367 13515
rect 12725 13481 12759 13515
rect 2881 13413 2915 13447
rect 1409 13345 1443 13379
rect 4077 13345 4111 13379
rect 5273 13345 5307 13379
rect 5540 13345 5574 13379
rect 7665 13345 7699 13379
rect 11601 13345 11635 13379
rect 3065 13277 3099 13311
rect 8677 13277 8711 13311
rect 11345 13277 11379 13311
rect 1685 12937 1719 12971
rect 3985 12937 4019 12971
rect 10517 12937 10551 12971
rect 12081 12937 12115 12971
rect 5733 12801 5767 12835
rect 11161 12801 11195 12835
rect 1501 12733 1535 12767
rect 2605 12733 2639 12767
rect 7757 12733 7791 12767
rect 8013 12733 8047 12767
rect 12265 12733 12299 12767
rect 2872 12665 2906 12699
rect 5549 12665 5583 12699
rect 10885 12665 10919 12699
rect 12449 12665 12483 12699
rect 5181 12597 5215 12631
rect 5641 12597 5675 12631
rect 9137 12597 9171 12631
rect 10977 12597 11011 12631
rect 1409 12393 1443 12427
rect 6929 12393 6963 12427
rect 7849 12393 7883 12427
rect 11069 12393 11103 12427
rect 4353 12325 4387 12359
rect 12142 12325 12176 12359
rect 2789 12257 2823 12291
rect 4077 12257 4111 12291
rect 5549 12257 5583 12291
rect 5805 12257 5839 12291
rect 8217 12257 8251 12291
rect 9689 12257 9723 12291
rect 9945 12257 9979 12291
rect 11897 12257 11931 12291
rect 19717 12257 19751 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 2421 12121 2455 12155
rect 13277 12053 13311 12087
rect 19901 12053 19935 12087
rect 3341 11849 3375 11883
rect 7021 11849 7055 11883
rect 9689 11849 9723 11883
rect 9873 11849 9907 11883
rect 10701 11849 10735 11883
rect 8309 11713 8343 11747
rect 10425 11713 10459 11747
rect 11253 11713 11287 11747
rect 1961 11645 1995 11679
rect 4537 11645 4571 11679
rect 4804 11645 4838 11679
rect 6837 11645 6871 11679
rect 8576 11645 8610 11679
rect 11069 11645 11103 11679
rect 19625 11645 19659 11679
rect 2228 11577 2262 11611
rect 5917 11509 5951 11543
rect 10241 11509 10275 11543
rect 10333 11509 10367 11543
rect 11161 11509 11195 11543
rect 13277 11509 13311 11543
rect 19809 11509 19843 11543
rect 2421 11305 2455 11339
rect 2789 11305 2823 11339
rect 6929 11305 6963 11339
rect 8033 11305 8067 11339
rect 8401 11305 8435 11339
rect 12265 11305 12299 11339
rect 5794 11237 5828 11271
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 7941 11169 7975 11203
rect 8493 11169 8527 11203
rect 10425 11169 10459 11203
rect 12541 11169 12575 11203
rect 12808 11169 12842 11203
rect 19073 11169 19107 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 5549 11101 5583 11135
rect 8585 11101 8619 11135
rect 15853 11101 15887 11135
rect 7757 11033 7791 11067
rect 11713 11033 11747 11067
rect 19257 11033 19291 11067
rect 13921 10965 13955 10999
rect 2053 10761 2087 10795
rect 4997 10761 5031 10795
rect 10149 10761 10183 10795
rect 12081 10761 12115 10795
rect 8217 10693 8251 10727
rect 13829 10693 13863 10727
rect 14657 10693 14691 10727
rect 2605 10625 2639 10659
rect 3617 10625 3651 10659
rect 7113 10625 7147 10659
rect 8861 10625 8895 10659
rect 10793 10625 10827 10659
rect 15209 10625 15243 10659
rect 2421 10557 2455 10591
rect 2513 10557 2547 10591
rect 3884 10557 3918 10591
rect 6929 10557 6963 10591
rect 8677 10557 8711 10591
rect 12265 10557 12299 10591
rect 12449 10557 12483 10591
rect 18521 10557 18555 10591
rect 12716 10489 12750 10523
rect 15025 10489 15059 10523
rect 8585 10421 8619 10455
rect 10517 10421 10551 10455
rect 10609 10421 10643 10455
rect 15117 10421 15151 10455
rect 16221 10421 16255 10455
rect 18705 10421 18739 10455
rect 2789 10217 2823 10251
rect 4261 10217 4295 10251
rect 7021 10217 7055 10251
rect 8033 10217 8067 10251
rect 10517 10217 10551 10251
rect 8493 10149 8527 10183
rect 1676 10081 1710 10115
rect 4077 10081 4111 10115
rect 5825 10081 5859 10115
rect 8401 10081 8435 10115
rect 10854 10149 10888 10183
rect 13277 10081 13311 10115
rect 15568 10081 15602 10115
rect 17509 10081 17543 10115
rect 1409 10013 1443 10047
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 8677 10013 8711 10047
rect 10517 10013 10551 10047
rect 10609 10013 10643 10047
rect 13369 10013 13403 10047
rect 13553 10013 13587 10047
rect 15301 10013 15335 10047
rect 17785 10013 17819 10047
rect 5457 9877 5491 9911
rect 11989 9877 12023 9911
rect 12909 9877 12943 9911
rect 16681 9877 16715 9911
rect 16221 9673 16255 9707
rect 3341 9605 3375 9639
rect 4721 9605 4755 9639
rect 10609 9605 10643 9639
rect 5365 9537 5399 9571
rect 11161 9537 11195 9571
rect 13553 9537 13587 9571
rect 13737 9537 13771 9571
rect 1961 9469 1995 9503
rect 5089 9469 5123 9503
rect 6653 9469 6687 9503
rect 7481 9469 7515 9503
rect 7748 9469 7782 9503
rect 11069 9469 11103 9503
rect 14841 9469 14875 9503
rect 18061 9469 18095 9503
rect 2228 9401 2262 9435
rect 15108 9401 15142 9435
rect 18337 9401 18371 9435
rect 5181 9333 5215 9367
rect 6469 9333 6503 9367
rect 8861 9333 8895 9367
rect 10977 9333 11011 9367
rect 13093 9333 13127 9367
rect 13461 9333 13495 9367
rect 1409 9129 1443 9163
rect 2789 9129 2823 9163
rect 8493 9129 8527 9163
rect 9689 9129 9723 9163
rect 13185 9129 13219 9163
rect 13461 9129 13495 9163
rect 15577 9129 15611 9163
rect 15945 9129 15979 9163
rect 18797 9129 18831 9163
rect 5172 9061 5206 9095
rect 7358 9061 7392 9095
rect 2881 8993 2915 9027
rect 10793 8993 10827 9027
rect 11060 8993 11094 9027
rect 13369 8993 13403 9027
rect 15117 8993 15151 9027
rect 16037 8993 16071 9027
rect 17684 8993 17718 9027
rect 3065 8925 3099 8959
rect 4905 8925 4939 8959
rect 7113 8925 7147 8959
rect 16129 8925 16163 8959
rect 17417 8925 17451 8959
rect 19625 8925 19659 8959
rect 2421 8789 2455 8823
rect 6285 8789 6319 8823
rect 12173 8789 12207 8823
rect 14933 8789 14967 8823
rect 1869 8585 1903 8619
rect 3433 8585 3467 8619
rect 5089 8585 5123 8619
rect 9137 8585 9171 8619
rect 9965 8585 9999 8619
rect 11713 8585 11747 8619
rect 19349 8585 19383 8619
rect 18245 8517 18279 8551
rect 2513 8449 2547 8483
rect 4077 8449 4111 8483
rect 5733 8449 5767 8483
rect 10609 8449 10643 8483
rect 13185 8449 13219 8483
rect 15761 8449 15795 8483
rect 2237 8381 2271 8415
rect 2329 8381 2363 8415
rect 5549 8381 5583 8415
rect 7757 8381 7791 8415
rect 8024 8381 8058 8415
rect 10333 8381 10367 8415
rect 11897 8381 11931 8415
rect 15485 8381 15519 8415
rect 16773 8381 16807 8415
rect 18061 8381 18095 8415
rect 19165 8381 19199 8415
rect 5457 8313 5491 8347
rect 10425 8313 10459 8347
rect 13452 8313 13486 8347
rect 20269 8313 20303 8347
rect 3801 8245 3835 8279
rect 3893 8245 3927 8279
rect 14565 8245 14599 8279
rect 16957 8245 16991 8279
rect 2053 8041 2087 8075
rect 4997 8041 5031 8075
rect 6653 8041 6687 8075
rect 18889 8041 18923 8075
rect 12234 7973 12268 8007
rect 15546 7973 15580 8007
rect 2421 7905 2455 7939
rect 5181 7905 5215 7939
rect 5540 7905 5574 7939
rect 7665 7905 7699 7939
rect 8401 7905 8435 7939
rect 9956 7905 9990 7939
rect 11989 7905 12023 7939
rect 17509 7905 17543 7939
rect 17776 7905 17810 7939
rect 19717 7905 19751 7939
rect 2513 7837 2547 7871
rect 2697 7837 2731 7871
rect 5273 7837 5307 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 9689 7837 9723 7871
rect 14197 7837 14231 7871
rect 15301 7837 15335 7871
rect 7481 7701 7515 7735
rect 8033 7701 8067 7735
rect 11069 7701 11103 7735
rect 13369 7701 13403 7735
rect 16681 7701 16715 7735
rect 19901 7701 19935 7735
rect 6929 7497 6963 7531
rect 10701 7497 10735 7531
rect 16865 7497 16899 7531
rect 1409 7361 1443 7395
rect 7481 7361 7515 7395
rect 11253 7361 11287 7395
rect 13001 7361 13035 7395
rect 18705 7361 18739 7395
rect 3617 7293 3651 7327
rect 7389 7293 7423 7327
rect 8493 7293 8527 7327
rect 12909 7293 12943 7327
rect 14013 7293 14047 7327
rect 15485 7293 15519 7327
rect 15752 7293 15786 7327
rect 19625 7293 19659 7327
rect 1676 7225 1710 7259
rect 3862 7225 3896 7259
rect 8738 7225 8772 7259
rect 14289 7225 14323 7259
rect 2789 7157 2823 7191
rect 4997 7157 5031 7191
rect 7297 7157 7331 7191
rect 9873 7157 9907 7191
rect 11069 7157 11103 7191
rect 11161 7157 11195 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 18061 7157 18095 7191
rect 18429 7157 18463 7191
rect 18521 7157 18555 7191
rect 19809 7157 19843 7191
rect 2237 6953 2271 6987
rect 13277 6953 13311 6987
rect 15669 6953 15703 6987
rect 19257 6953 19291 6987
rect 19625 6953 19659 6987
rect 2605 6885 2639 6919
rect 4322 6885 4356 6919
rect 11621 6885 11655 6919
rect 13369 6885 13403 6919
rect 18061 6885 18095 6919
rect 4077 6817 4111 6851
rect 6285 6817 6319 6851
rect 7389 6817 7423 6851
rect 7656 6817 7690 6851
rect 10057 6817 10091 6851
rect 14657 6817 14691 6851
rect 17509 6817 17543 6851
rect 18153 6817 18187 6851
rect 19717 6817 19751 6851
rect 2697 6749 2731 6783
rect 2789 6749 2823 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 13461 6749 13495 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 18245 6749 18279 6783
rect 19809 6749 19843 6783
rect 9689 6681 9723 6715
rect 12909 6681 12943 6715
rect 14473 6681 14507 6715
rect 15301 6681 15335 6715
rect 17693 6681 17727 6715
rect 5457 6613 5491 6647
rect 8769 6613 8803 6647
rect 11253 6613 11287 6647
rect 1685 6409 1719 6443
rect 5181 6409 5215 6443
rect 8217 6409 8251 6443
rect 13829 6409 13863 6443
rect 20453 6409 20487 6443
rect 3249 6341 3283 6375
rect 2329 6273 2363 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 5733 6273 5767 6307
rect 9137 6273 9171 6307
rect 10149 6273 10183 6307
rect 14289 6273 14323 6307
rect 14473 6273 14507 6307
rect 16313 6273 16347 6307
rect 2053 6205 2087 6239
rect 3617 6205 3651 6239
rect 5641 6205 5675 6239
rect 6837 6205 6871 6239
rect 10405 6205 10439 6239
rect 12541 6205 12575 6239
rect 14197 6205 14231 6239
rect 19073 6205 19107 6239
rect 7104 6137 7138 6171
rect 12817 6137 12851 6171
rect 16037 6137 16071 6171
rect 18061 6137 18095 6171
rect 19340 6137 19374 6171
rect 2145 6069 2179 6103
rect 5549 6069 5583 6103
rect 11529 6069 11563 6103
rect 15669 6069 15703 6103
rect 16129 6069 16163 6103
rect 4077 5865 4111 5899
rect 8493 5865 8527 5899
rect 9781 5865 9815 5899
rect 13645 5865 13679 5899
rect 4445 5797 4479 5831
rect 10149 5797 10183 5831
rect 11590 5797 11624 5831
rect 14105 5797 14139 5831
rect 2697 5729 2731 5763
rect 5641 5729 5675 5763
rect 5908 5729 5942 5763
rect 8401 5729 8435 5763
rect 11345 5729 11379 5763
rect 14013 5729 14047 5763
rect 15557 5729 15591 5763
rect 18696 5729 18730 5763
rect 2789 5661 2823 5695
rect 2973 5661 3007 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 8677 5661 8711 5695
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 14289 5661 14323 5695
rect 15301 5661 15335 5695
rect 18429 5661 18463 5695
rect 8033 5593 8067 5627
rect 2329 5525 2363 5559
rect 7021 5525 7055 5559
rect 12725 5525 12759 5559
rect 16681 5525 16715 5559
rect 19809 5525 19843 5559
rect 1777 5321 1811 5355
rect 6837 5321 6871 5355
rect 8401 5321 8435 5355
rect 12633 5321 12667 5355
rect 14933 5321 14967 5355
rect 4629 5253 4663 5287
rect 10793 5253 10827 5287
rect 2421 5185 2455 5219
rect 3341 5185 3375 5219
rect 5181 5185 5215 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 8953 5185 8987 5219
rect 11345 5185 11379 5219
rect 4997 5117 5031 5151
rect 12449 5117 12483 5151
rect 13553 5117 13587 5151
rect 15761 5117 15795 5151
rect 16028 5117 16062 5151
rect 18061 5117 18095 5151
rect 20269 5117 20303 5151
rect 2145 5049 2179 5083
rect 7205 5049 7239 5083
rect 8769 5049 8803 5083
rect 11253 5049 11287 5083
rect 13820 5049 13854 5083
rect 18306 5049 18340 5083
rect 2237 4981 2271 5015
rect 5089 4981 5123 5015
rect 8861 4981 8895 5015
rect 11161 4981 11195 5015
rect 17141 4981 17175 5015
rect 19441 4981 19475 5015
rect 20453 4981 20487 5015
rect 3157 4777 3191 4811
rect 4077 4777 4111 4811
rect 6837 4777 6871 4811
rect 19073 4777 19107 4811
rect 12786 4709 12820 4743
rect 16672 4709 16706 4743
rect 1777 4641 1811 4675
rect 2044 4641 2078 4675
rect 5457 4641 5491 4675
rect 5724 4641 5758 4675
rect 8033 4641 8067 4675
rect 10057 4641 10091 4675
rect 11437 4641 11471 4675
rect 15301 4641 15335 4675
rect 16405 4641 16439 4675
rect 8125 4573 8159 4607
rect 8217 4573 8251 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 12541 4573 12575 4607
rect 19165 4573 19199 4607
rect 19349 4573 19383 4607
rect 9689 4505 9723 4539
rect 7665 4437 7699 4471
rect 11621 4437 11655 4471
rect 13921 4437 13955 4471
rect 15485 4437 15519 4471
rect 17785 4437 17819 4471
rect 18705 4437 18739 4471
rect 6837 4233 6871 4267
rect 9321 4233 9355 4267
rect 4813 4165 4847 4199
rect 11437 4165 11471 4199
rect 2513 4097 2547 4131
rect 3433 4097 3467 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 9965 4097 9999 4131
rect 13001 4097 13035 4131
rect 14565 4097 14599 4131
rect 16497 4097 16531 4131
rect 18337 4097 18371 4131
rect 3689 4029 3723 4063
rect 11253 4029 11287 4063
rect 12909 4029 12943 4063
rect 14381 4029 14415 4063
rect 16313 4029 16347 4063
rect 18061 4029 18095 4063
rect 19441 4029 19475 4063
rect 19708 4029 19742 4063
rect 5733 3961 5767 3995
rect 7205 3961 7239 3995
rect 9689 3961 9723 3995
rect 14473 3961 14507 3995
rect 1869 3893 1903 3927
rect 2237 3893 2271 3927
rect 2329 3893 2363 3927
rect 9781 3893 9815 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 14013 3893 14047 3927
rect 15853 3893 15887 3927
rect 16221 3893 16255 3927
rect 20821 3893 20855 3927
rect 2421 3689 2455 3723
rect 7205 3689 7239 3723
rect 8401 3689 8435 3723
rect 11069 3689 11103 3723
rect 16957 3689 16991 3723
rect 18061 3689 18095 3723
rect 2881 3621 2915 3655
rect 12265 3621 12299 3655
rect 2789 3553 2823 3587
rect 4629 3553 4663 3587
rect 4896 3553 4930 3587
rect 9689 3553 9723 3587
rect 9956 3553 9990 3587
rect 12357 3553 12391 3587
rect 13461 3553 13495 3587
rect 13737 3553 13771 3587
rect 15301 3553 15335 3587
rect 16865 3553 16899 3587
rect 18429 3553 18463 3587
rect 18889 3553 18923 3587
rect 19717 3553 19751 3587
rect 3065 3485 3099 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 12541 3485 12575 3519
rect 17141 3485 17175 3519
rect 18521 3485 18555 3519
rect 18705 3485 18739 3519
rect 6009 3417 6043 3451
rect 17969 3417 18003 3451
rect 6837 3349 6871 3383
rect 11897 3349 11931 3383
rect 15485 3349 15519 3383
rect 16497 3349 16531 3383
rect 19901 3349 19935 3383
rect 2881 3145 2915 3179
rect 5549 3145 5583 3179
rect 12449 3145 12483 3179
rect 1501 3009 1535 3043
rect 7757 3009 7791 3043
rect 7941 3009 7975 3043
rect 8861 3009 8895 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 14565 3009 14599 3043
rect 15853 3009 15887 3043
rect 16957 3009 16991 3043
rect 19533 3009 19567 3043
rect 4169 2941 4203 2975
rect 7665 2941 7699 2975
rect 11069 2941 11103 2975
rect 14391 2941 14425 2975
rect 15669 2941 15703 2975
rect 18061 2941 18095 2975
rect 19349 2941 19383 2975
rect 20821 2941 20855 2975
rect 1768 2873 1802 2907
rect 4436 2873 4470 2907
rect 9128 2873 9162 2907
rect 11345 2873 11379 2907
rect 18337 2873 18371 2907
rect 7297 2805 7331 2839
rect 10241 2805 10275 2839
rect 12817 2805 12851 2839
rect 2421 2601 2455 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8677 2601 8711 2635
rect 11161 2601 11195 2635
rect 12633 2601 12667 2635
rect 17233 2601 17267 2635
rect 19625 2601 19659 2635
rect 2881 2533 2915 2567
rect 4537 2533 4571 2567
rect 11253 2533 11287 2567
rect 13001 2533 13035 2567
rect 16037 2533 16071 2567
rect 2789 2465 2823 2499
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 7297 2465 7331 2499
rect 9781 2465 9815 2499
rect 14197 2465 14231 2499
rect 15761 2465 15795 2499
rect 17049 2465 17083 2499
rect 18337 2465 18371 2499
rect 19441 2465 19475 2499
rect 3065 2397 3099 2431
rect 5825 2397 5859 2431
rect 7573 2397 7607 2431
rect 11345 2397 11379 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 10793 2329 10827 2363
rect 14381 2261 14415 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 12802 20992 12808 21004
rect 4120 20964 12808 20992
rect 4120 20952 4126 20964
rect 12802 20952 12808 20964
rect 12860 20952 12866 21004
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 12526 20924 12532 20936
rect 4028 20896 12532 20924
rect 4028 20884 4034 20896
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 13906 20856 13912 20868
rect 3844 20828 13912 20856
rect 3844 20816 3850 20828
rect 13906 20816 13912 20828
rect 13964 20816 13970 20868
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 13630 20788 13636 20800
rect 3936 20760 13636 20788
rect 3936 20748 3942 20760
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 4028 20556 9965 20584
rect 4028 20544 4034 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 12802 20584 12808 20596
rect 12763 20556 12808 20584
rect 9953 20547 10011 20553
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 13906 20584 13912 20596
rect 13867 20556 13912 20584
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 4062 20476 4068 20528
rect 4120 20516 4126 20528
rect 11057 20519 11115 20525
rect 11057 20516 11069 20519
rect 4120 20488 11069 20516
rect 4120 20476 4126 20488
rect 11057 20485 11069 20488
rect 11103 20485 11115 20519
rect 11057 20479 11115 20485
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20448 2559 20451
rect 7098 20448 7104 20460
rect 2547 20420 5304 20448
rect 2547 20417 2559 20420
rect 2501 20411 2559 20417
rect 2222 20380 2228 20392
rect 2183 20352 2228 20380
rect 2222 20340 2228 20352
rect 2280 20340 2286 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 5166 20380 5172 20392
rect 4111 20352 5172 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 5276 20380 5304 20420
rect 6932 20420 7104 20448
rect 6932 20389 6960 20420
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 5341 20383 5399 20389
rect 5341 20380 5353 20383
rect 5276 20352 5353 20380
rect 5341 20349 5353 20352
rect 5387 20349 5399 20383
rect 5341 20343 5399 20349
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20349 6975 20383
rect 6917 20343 6975 20349
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7064 20352 8033 20380
rect 7064 20340 7070 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 9766 20380 9772 20392
rect 9727 20352 9772 20380
rect 8021 20343 8079 20349
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 10870 20380 10876 20392
rect 10831 20352 10876 20380
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 12618 20380 12624 20392
rect 12579 20352 12624 20380
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 13722 20380 13728 20392
rect 13683 20352 13728 20380
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 4341 20315 4399 20321
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 11238 20312 11244 20324
rect 4387 20284 11244 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 3510 20204 3516 20256
rect 3568 20244 3574 20256
rect 5537 20247 5595 20253
rect 5537 20244 5549 20247
rect 3568 20216 5549 20244
rect 3568 20204 3574 20216
rect 5537 20213 5549 20216
rect 5583 20213 5595 20247
rect 5537 20207 5595 20213
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 7064 20216 7113 20244
rect 7064 20204 7070 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 7101 20207 7159 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 10870 20040 10876 20052
rect 4356 20012 10876 20040
rect 4356 19981 4384 20012
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12621 20043 12679 20049
rect 12621 20040 12633 20043
rect 12584 20012 12633 20040
rect 12584 20000 12590 20012
rect 12621 20009 12633 20012
rect 12667 20009 12679 20043
rect 12621 20003 12679 20009
rect 4341 19975 4399 19981
rect 4341 19941 4353 19975
rect 4387 19941 4399 19975
rect 8202 19972 8208 19984
rect 4341 19935 4399 19941
rect 4448 19944 8208 19972
rect 2130 19904 2136 19916
rect 2091 19876 2136 19904
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 2406 19904 2412 19916
rect 2367 19876 2412 19904
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4080 19836 4108 19867
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 4448 19904 4476 19944
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 9766 19932 9772 19984
rect 9824 19972 9830 19984
rect 9953 19975 10011 19981
rect 9953 19972 9965 19975
rect 9824 19944 9965 19972
rect 9824 19932 9830 19944
rect 9953 19941 9965 19944
rect 9999 19941 10011 19975
rect 9953 19935 10011 19941
rect 11425 19975 11483 19981
rect 11425 19941 11437 19975
rect 11471 19972 11483 19975
rect 13722 19972 13728 19984
rect 11471 19944 13728 19972
rect 11471 19941 11483 19944
rect 11425 19935 11483 19941
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 5350 19904 5356 19916
rect 4212 19876 4476 19904
rect 5311 19876 5356 19904
rect 4212 19864 4218 19876
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 6638 19904 6644 19916
rect 5460 19876 6500 19904
rect 6599 19876 6644 19904
rect 5460 19836 5488 19876
rect 5626 19836 5632 19848
rect 4080 19808 5488 19836
rect 5587 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 6472 19836 6500 19876
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 8294 19904 8300 19916
rect 8255 19876 8300 19904
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8754 19904 8760 19916
rect 8404 19876 8760 19904
rect 8404 19836 8432 19876
rect 8754 19864 8760 19876
rect 8812 19864 8818 19916
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 10502 19904 10508 19916
rect 9723 19876 10508 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19873 11207 19907
rect 11149 19867 11207 19873
rect 8570 19836 8576 19848
rect 6472 19808 8432 19836
rect 8531 19808 8576 19836
rect 8570 19796 8576 19808
rect 8628 19796 8634 19848
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 10962 19836 10968 19848
rect 8720 19808 10968 19836
rect 8720 19796 8726 19808
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 8754 19728 8760 19780
rect 8812 19768 8818 19780
rect 10042 19768 10048 19780
rect 8812 19740 10048 19768
rect 8812 19728 8818 19740
rect 10042 19728 10048 19740
rect 10100 19728 10106 19780
rect 11164 19768 11192 19867
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 11296 19876 12449 19904
rect 11296 19864 11302 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19873 13599 19907
rect 17218 19904 17224 19916
rect 17179 19876 17224 19904
rect 13541 19867 13599 19873
rect 12434 19768 12440 19780
rect 11164 19740 12440 19768
rect 12434 19728 12440 19740
rect 12492 19728 12498 19780
rect 13556 19768 13584 19867
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 12544 19740 13584 19768
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 6825 19703 6883 19709
rect 6825 19700 6837 19703
rect 3936 19672 6837 19700
rect 3936 19660 3942 19672
rect 6825 19669 6837 19672
rect 6871 19669 6883 19703
rect 6825 19663 6883 19669
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 12544 19700 12572 19740
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 13725 19771 13783 19777
rect 13725 19768 13737 19771
rect 13688 19740 13737 19768
rect 13688 19728 13694 19740
rect 13725 19737 13737 19740
rect 13771 19737 13783 19771
rect 13725 19731 13783 19737
rect 8628 19672 12572 19700
rect 8628 19660 8634 19672
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 7650 19496 7656 19508
rect 2280 19468 7656 19496
rect 2280 19456 2286 19468
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 9125 19499 9183 19505
rect 9125 19496 9137 19499
rect 8352 19468 9137 19496
rect 8352 19456 8358 19468
rect 9125 19465 9137 19468
rect 9171 19465 9183 19499
rect 12434 19496 12440 19508
rect 12395 19468 12440 19496
rect 9125 19459 9183 19465
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 5626 19388 5632 19440
rect 5684 19428 5690 19440
rect 12618 19428 12624 19440
rect 5684 19400 12624 19428
rect 5684 19388 5690 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19360 4951 19363
rect 5166 19360 5172 19372
rect 4939 19332 5172 19360
rect 4939 19329 4951 19332
rect 4893 19323 4951 19329
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 7466 19360 7472 19372
rect 7427 19332 7472 19360
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 11422 19360 11428 19372
rect 9815 19332 11428 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13998 19360 14004 19372
rect 13127 19332 14004 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2363 19264 6868 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2593 19227 2651 19233
rect 2593 19193 2605 19227
rect 2639 19224 2651 19227
rect 6730 19224 6736 19236
rect 2639 19196 6736 19224
rect 2639 19193 2651 19196
rect 2593 19187 2651 19193
rect 6730 19184 6736 19196
rect 6788 19184 6794 19236
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 4249 19159 4307 19165
rect 4249 19156 4261 19159
rect 2464 19128 4261 19156
rect 2464 19116 2470 19128
rect 4249 19125 4261 19128
rect 4295 19125 4307 19159
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4249 19119 4307 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 4890 19156 4896 19168
rect 4755 19128 4896 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 6840 19165 6868 19264
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 8536 19264 10701 19292
rect 8536 19252 8542 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 20579 19264 20613 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 7193 19227 7251 19233
rect 7193 19193 7205 19227
rect 7239 19224 7251 19227
rect 12986 19224 12992 19236
rect 7239 19196 12992 19224
rect 7239 19193 7251 19196
rect 7193 19187 7251 19193
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 20441 19227 20499 19233
rect 20441 19193 20453 19227
rect 20487 19224 20499 19227
rect 20548 19224 20576 19255
rect 20898 19224 20904 19236
rect 20487 19196 20904 19224
rect 20487 19193 20499 19196
rect 20441 19187 20499 19193
rect 20898 19184 20904 19196
rect 20956 19184 20962 19236
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 9490 19156 9496 19168
rect 7340 19128 7385 19156
rect 9451 19128 9496 19156
rect 7340 19116 7346 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9585 19159 9643 19165
rect 9585 19125 9597 19159
rect 9631 19156 9643 19159
rect 9674 19156 9680 19168
rect 9631 19128 9680 19156
rect 9631 19125 9643 19128
rect 9585 19119 9643 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 9824 19128 10885 19156
rect 9824 19116 9830 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 12802 19156 12808 19168
rect 12763 19128 12808 19156
rect 10873 19119 10931 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 20714 19156 20720 19168
rect 12952 19128 12997 19156
rect 20675 19128 20720 19156
rect 12952 19116 12958 19128
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1397 18955 1455 18961
rect 1397 18921 1409 18955
rect 1443 18952 1455 18955
rect 4614 18952 4620 18964
rect 1443 18924 4620 18952
rect 1443 18921 1455 18924
rect 1397 18915 1455 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 6365 18955 6423 18961
rect 4816 18924 6132 18952
rect 2685 18887 2743 18893
rect 2685 18853 2697 18887
rect 2731 18884 2743 18887
rect 4816 18884 4844 18924
rect 2731 18856 4844 18884
rect 2731 18853 2743 18856
rect 2685 18847 2743 18853
rect 5166 18844 5172 18896
rect 5224 18893 5230 18896
rect 5224 18887 5288 18893
rect 5224 18853 5242 18887
rect 5276 18853 5288 18887
rect 5224 18847 5288 18853
rect 5224 18844 5230 18847
rect 2406 18816 2412 18828
rect 2367 18788 2412 18816
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4985 18751 5043 18757
rect 4985 18748 4997 18751
rect 3844 18720 4997 18748
rect 3844 18708 3850 18720
rect 4985 18717 4997 18720
rect 5031 18717 5043 18751
rect 6104 18748 6132 18924
rect 6365 18921 6377 18955
rect 6411 18921 6423 18955
rect 6365 18915 6423 18921
rect 6380 18816 6408 18915
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 7524 18924 8585 18952
rect 7524 18912 7530 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 9674 18952 9680 18964
rect 9635 18924 9680 18952
rect 8573 18915 8631 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 12860 18924 13461 18952
rect 12860 18912 12866 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 13449 18915 13507 18921
rect 7558 18884 7564 18896
rect 7484 18856 7564 18884
rect 7484 18825 7512 18856
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 11422 18844 11428 18896
rect 11480 18893 11486 18896
rect 11480 18887 11544 18893
rect 11480 18853 11498 18887
rect 11532 18853 11544 18887
rect 11480 18847 11544 18853
rect 11480 18844 11486 18847
rect 7449 18819 7512 18825
rect 7449 18816 7461 18819
rect 6380 18788 7461 18816
rect 7449 18785 7461 18788
rect 7495 18788 7512 18819
rect 7495 18785 7507 18788
rect 7449 18779 7507 18785
rect 8938 18776 8944 18828
rect 8996 18816 9002 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 8996 18788 10057 18816
rect 8996 18776 9002 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 11241 18819 11299 18825
rect 11241 18816 11253 18819
rect 10652 18788 11253 18816
rect 10652 18776 10658 18788
rect 11241 18785 11253 18788
rect 11287 18816 11299 18819
rect 12618 18816 12624 18828
rect 11287 18788 12624 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 7098 18748 7104 18760
rect 6104 18720 7104 18748
rect 4985 18711 5043 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 7190 18708 7196 18760
rect 7248 18748 7254 18760
rect 10137 18751 10195 18757
rect 7248 18720 7293 18748
rect 7248 18708 7254 18720
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 11054 18748 11060 18760
rect 10367 18720 11060 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10152 18680 10180 18711
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 10152 18652 10640 18680
rect 4062 18572 4068 18624
rect 4120 18612 4126 18624
rect 9766 18612 9772 18624
rect 4120 18584 9772 18612
rect 4120 18572 4126 18584
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 10612 18621 10640 18652
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 11974 18612 11980 18624
rect 10643 18584 11980 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 12710 18612 12716 18624
rect 12667 18584 12716 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 5166 18368 5172 18420
rect 5224 18408 5230 18420
rect 5445 18411 5503 18417
rect 5445 18408 5457 18411
rect 5224 18380 5457 18408
rect 5224 18368 5230 18380
rect 5445 18377 5457 18380
rect 5491 18377 5503 18411
rect 5445 18371 5503 18377
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 11238 18408 11244 18420
rect 5776 18380 11100 18408
rect 11199 18380 11244 18408
rect 5776 18368 5782 18380
rect 11072 18340 11100 18380
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 20714 18408 20720 18420
rect 11501 18380 20720 18408
rect 11501 18340 11529 18380
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 11072 18312 11529 18340
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 12618 18272 12624 18284
rect 2547 18244 4200 18272
rect 12579 18244 12624 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 3418 18204 3424 18216
rect 2271 18176 3424 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4065 18207 4123 18213
rect 4065 18204 4077 18207
rect 3844 18176 4077 18204
rect 3844 18164 3850 18176
rect 4065 18173 4077 18176
rect 4111 18173 4123 18207
rect 4172 18204 4200 18244
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 6638 18204 6644 18216
rect 4172 18176 6644 18204
rect 4065 18167 4123 18173
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7098 18204 7104 18216
rect 7055 18176 7104 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9824 18176 9873 18204
rect 9824 18164 9830 18176
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 9861 18167 9919 18173
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 12877 18207 12935 18213
rect 12877 18204 12889 18207
rect 12768 18176 12889 18204
rect 12768 18164 12774 18176
rect 12877 18173 12889 18176
rect 12923 18173 12935 18207
rect 12877 18167 12935 18173
rect 4332 18139 4390 18145
rect 4332 18105 4344 18139
rect 4378 18136 4390 18139
rect 5442 18136 5448 18148
rect 4378 18108 5448 18136
rect 4378 18105 4390 18108
rect 4332 18099 4390 18105
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 7276 18139 7334 18145
rect 7276 18105 7288 18139
rect 7322 18136 7334 18139
rect 7466 18136 7472 18148
rect 7322 18108 7472 18136
rect 7322 18105 7334 18108
rect 7276 18099 7334 18105
rect 7466 18096 7472 18108
rect 7524 18096 7530 18148
rect 8294 18136 8300 18148
rect 7576 18108 8300 18136
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 7576 18068 7604 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 10128 18139 10186 18145
rect 10128 18105 10140 18139
rect 10174 18136 10186 18139
rect 11054 18136 11060 18148
rect 10174 18108 11060 18136
rect 10174 18105 10186 18108
rect 10128 18099 10186 18105
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 8386 18068 8392 18080
rect 4120 18040 7604 18068
rect 8347 18040 8392 18068
rect 4120 18028 4126 18040
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 13998 18068 14004 18080
rect 13911 18040 14004 18068
rect 13998 18028 14004 18040
rect 14056 18068 14062 18080
rect 19242 18068 19248 18080
rect 14056 18040 19248 18068
rect 14056 18028 14062 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 4890 17864 4896 17876
rect 4851 17836 4896 17864
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7282 17864 7288 17876
rect 7055 17836 7288 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 8573 17867 8631 17873
rect 7423 17836 8248 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 6917 17799 6975 17805
rect 6917 17765 6929 17799
rect 6963 17796 6975 17799
rect 6963 17768 7512 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 7484 17740 7512 17768
rect 2214 17731 2272 17737
rect 2214 17697 2226 17731
rect 2260 17697 2272 17731
rect 2214 17691 2272 17697
rect 2231 17660 2259 17691
rect 4338 17688 4344 17740
rect 4396 17728 4402 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 4396 17700 5273 17728
rect 4396 17688 4402 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 6178 17728 6184 17740
rect 5399 17700 6184 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 2406 17660 2412 17672
rect 2231 17632 2412 17660
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 2501 17663 2559 17669
rect 2501 17629 2513 17663
rect 2547 17629 2559 17663
rect 2501 17623 2559 17629
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 5368 17660 5396 17691
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 7466 17728 7472 17740
rect 7427 17700 7472 17728
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 8220 17728 8248 17836
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 9490 17864 9496 17876
rect 8619 17836 9496 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17833 12127 17867
rect 12986 17864 12992 17876
rect 12947 17836 12992 17864
rect 12069 17827 12127 17833
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 12084 17796 12112 17827
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 8352 17768 12112 17796
rect 8352 17756 8358 17768
rect 8938 17728 8944 17740
rect 8220 17700 8944 17728
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 9766 17728 9772 17740
rect 9723 17700 9772 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 9944 17731 10002 17737
rect 9944 17697 9956 17731
rect 9990 17728 10002 17731
rect 10686 17728 10692 17740
rect 9990 17700 10692 17728
rect 9990 17697 10002 17700
rect 9944 17691 10002 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 11885 17731 11943 17737
rect 11885 17728 11897 17731
rect 11204 17700 11897 17728
rect 11204 17688 11210 17700
rect 11885 17697 11897 17700
rect 11931 17697 11943 17731
rect 11885 17691 11943 17697
rect 4847 17632 5396 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 2516 17592 2544 17623
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 7558 17660 7564 17672
rect 5500 17632 5545 17660
rect 7519 17632 7564 17660
rect 5500 17620 5506 17632
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 8478 17592 8484 17604
rect 2516 17564 8484 17592
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 7006 17524 7012 17536
rect 4120 17496 7012 17524
rect 4120 17484 4126 17496
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 5169 17323 5227 17329
rect 4120 17292 4752 17320
rect 4120 17280 4126 17292
rect 4724 17252 4752 17292
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5442 17320 5448 17332
rect 5215 17292 5448 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 9493 17323 9551 17329
rect 9493 17320 9505 17323
rect 5592 17292 9505 17320
rect 5592 17280 5598 17292
rect 9493 17289 9505 17292
rect 9539 17289 9551 17323
rect 9493 17283 9551 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10686 17320 10692 17332
rect 9824 17292 10692 17320
rect 9824 17280 9830 17292
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12894 17320 12900 17332
rect 12483 17292 12900 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 11241 17255 11299 17261
rect 11241 17252 11253 17255
rect 4724 17224 9987 17252
rect 8573 17187 8631 17193
rect 2056 17156 3924 17184
rect 2056 17116 2084 17156
rect 2122 17119 2180 17125
rect 2122 17116 2134 17119
rect 2056 17088 2134 17116
rect 2122 17085 2134 17088
rect 2168 17085 2180 17119
rect 3786 17116 3792 17128
rect 3747 17088 3792 17116
rect 2122 17079 2180 17085
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 3896 17116 3924 17156
rect 8573 17153 8585 17187
rect 8619 17184 8631 17187
rect 9766 17184 9772 17196
rect 8619 17156 9772 17184
rect 8619 17153 8631 17156
rect 8573 17147 8631 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 9959 17184 9987 17224
rect 10051 17224 11253 17252
rect 10051 17184 10079 17224
rect 11241 17221 11253 17224
rect 11287 17221 11299 17255
rect 11241 17215 11299 17221
rect 9959 17156 10079 17184
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10318 17184 10324 17196
rect 10183 17156 10324 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12768 17156 13001 17184
rect 12768 17144 12774 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 5166 17116 5172 17128
rect 3896 17088 5172 17116
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 6972 17088 11069 17116
rect 6972 17076 6978 17088
rect 11057 17085 11069 17088
rect 11103 17085 11115 17119
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 11057 17079 11115 17085
rect 11808 17088 12817 17116
rect 2409 17051 2467 17057
rect 2409 17017 2421 17051
rect 2455 17048 2467 17051
rect 3694 17048 3700 17060
rect 2455 17020 3700 17048
rect 2455 17017 2467 17020
rect 2409 17011 2467 17017
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 4056 17051 4114 17057
rect 4056 17017 4068 17051
rect 4102 17048 4114 17051
rect 4982 17048 4988 17060
rect 4102 17020 4988 17048
rect 4102 17017 4114 17020
rect 4056 17011 4114 17017
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 8389 17051 8447 17057
rect 5408 17020 7972 17048
rect 5408 17008 5414 17020
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 7944 16989 7972 17020
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 9766 17048 9772 17060
rect 8435 17020 9772 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 9861 17051 9919 17057
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 11698 17048 11704 17060
rect 9907 17020 11704 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 4212 16952 7021 16980
rect 4212 16940 4218 16952
rect 7009 16949 7021 16952
rect 7055 16949 7067 16983
rect 7009 16943 7067 16949
rect 7929 16983 7987 16989
rect 7929 16949 7941 16983
rect 7975 16949 7987 16983
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 7929 16943 7987 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10008 16952 10053 16980
rect 10008 16940 10014 16952
rect 10410 16940 10416 16992
rect 10468 16980 10474 16992
rect 11808 16980 11836 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 12894 16980 12900 16992
rect 10468 16952 11836 16980
rect 12855 16952 12900 16980
rect 10468 16940 10474 16952
rect 12894 16940 12900 16952
rect 12952 16980 12958 16992
rect 13265 16983 13323 16989
rect 13265 16980 13277 16983
rect 12952 16952 13277 16980
rect 12952 16940 12958 16952
rect 13265 16949 13277 16952
rect 13311 16949 13323 16983
rect 13265 16943 13323 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 2188 16748 2421 16776
rect 2188 16736 2194 16748
rect 2409 16745 2421 16748
rect 2455 16745 2467 16779
rect 2409 16739 2467 16745
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 9674 16776 9680 16788
rect 3752 16748 9680 16776
rect 3752 16736 3758 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 11977 16779 12035 16785
rect 11977 16776 11989 16779
rect 10744 16748 11989 16776
rect 10744 16736 10750 16748
rect 11977 16745 11989 16748
rect 12023 16745 12035 16779
rect 11977 16739 12035 16745
rect 5905 16711 5963 16717
rect 4172 16680 5672 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 1443 16612 2789 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 4172 16640 4200 16680
rect 2777 16603 2835 16609
rect 4080 16612 4200 16640
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3068 16436 3096 16535
rect 4080 16513 4108 16612
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4304 16612 4445 16640
rect 4304 16600 4310 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 5534 16640 5540 16652
rect 4571 16612 5540 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5644 16649 5672 16680
rect 5905 16677 5917 16711
rect 5951 16708 5963 16711
rect 6914 16708 6920 16720
rect 5951 16680 6920 16708
rect 5951 16677 5963 16680
rect 5905 16671 5963 16677
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 8352 16680 12817 16708
rect 8352 16668 8358 16680
rect 12805 16677 12817 16680
rect 12851 16677 12863 16711
rect 12805 16671 12863 16677
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 7184 16643 7242 16649
rect 7184 16609 7196 16643
rect 7230 16640 7242 16643
rect 8386 16640 8392 16652
rect 7230 16612 8392 16640
rect 7230 16609 7242 16612
rect 7184 16603 7242 16609
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 10410 16640 10416 16652
rect 8496 16612 10416 16640
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4982 16572 4988 16584
rect 4755 16544 4988 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 6914 16572 6920 16584
rect 6875 16544 6920 16572
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 8496 16572 8524 16612
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10864 16643 10922 16649
rect 10864 16609 10876 16643
rect 10910 16640 10922 16643
rect 11146 16640 11152 16652
rect 10910 16612 11152 16640
rect 10910 16609 10922 16612
rect 10864 16603 10922 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 8260 16544 8524 16572
rect 8260 16532 8266 16544
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 8294 16436 8300 16448
rect 3068 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 4338 16232 4344 16244
rect 3660 16204 4344 16232
rect 3660 16192 3666 16204
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5040 16204 5733 16232
rect 5040 16192 5046 16204
rect 5721 16201 5733 16204
rect 5767 16201 5779 16235
rect 5721 16195 5779 16201
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 9824 16204 12449 16232
rect 9824 16192 9830 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 12437 16195 12495 16201
rect 11146 16164 11152 16176
rect 11059 16136 11152 16164
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 11164 16096 11192 16124
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 2547 16068 4476 16096
rect 11164 16068 13001 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 2314 16028 2320 16040
rect 2271 16000 2320 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 4028 16000 4353 16028
rect 4028 15988 4034 16000
rect 4341 15997 4353 16000
rect 4387 15997 4399 16031
rect 4448 16028 4476 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 6822 16028 6828 16040
rect 4448 16000 6828 16028
rect 4341 15991 4399 15997
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 6972 16000 7389 16028
rect 6972 15988 6978 16000
rect 7377 15997 7389 16000
rect 7423 16028 7435 16031
rect 9582 16028 9588 16040
rect 7423 16000 9588 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 9582 15988 9588 16000
rect 9640 16028 9646 16040
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9640 16000 9781 16028
rect 9640 15988 9646 16000
rect 9769 15997 9781 16000
rect 9815 16028 9827 16031
rect 9858 16028 9864 16040
rect 9815 16000 9864 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 11698 15988 11704 16040
rect 11756 16028 11762 16040
rect 14001 16031 14059 16037
rect 14001 16028 14013 16031
rect 11756 16000 14013 16028
rect 11756 15988 11762 16000
rect 14001 15997 14013 16000
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 4608 15963 4666 15969
rect 4608 15929 4620 15963
rect 4654 15960 4666 15963
rect 5442 15960 5448 15972
rect 4654 15932 5448 15960
rect 4654 15929 4666 15932
rect 4608 15923 4666 15929
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 7644 15963 7702 15969
rect 7644 15929 7656 15963
rect 7690 15960 7702 15963
rect 8294 15960 8300 15972
rect 7690 15932 8300 15960
rect 7690 15929 7702 15932
rect 7644 15923 7702 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 10036 15963 10094 15969
rect 10036 15929 10048 15963
rect 10082 15960 10094 15963
rect 10134 15960 10140 15972
rect 10082 15932 10140 15960
rect 10082 15929 10094 15932
rect 10036 15923 10094 15929
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 8478 15892 8484 15904
rect 4120 15864 8484 15892
rect 4120 15852 4126 15864
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 8754 15892 8760 15904
rect 8715 15864 8760 15892
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 8904 15864 12817 15892
rect 8904 15852 8910 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13170 15892 13176 15904
rect 12943 15864 13176 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13170 15852 13176 15864
rect 13228 15892 13234 15904
rect 13265 15895 13323 15901
rect 13265 15892 13277 15895
rect 13228 15864 13277 15892
rect 13228 15852 13234 15864
rect 13265 15861 13277 15864
rect 13311 15861 13323 15895
rect 13265 15855 13323 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 5258 15688 5264 15700
rect 4488 15660 5264 15688
rect 4488 15648 4494 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 5592 15660 6285 15688
rect 5592 15648 5598 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 6641 15691 6699 15697
rect 6641 15657 6653 15691
rect 6687 15688 6699 15691
rect 6687 15660 7696 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 4332 15623 4390 15629
rect 4332 15589 4344 15623
rect 4378 15620 4390 15623
rect 4798 15620 4804 15632
rect 4378 15592 4804 15620
rect 4378 15589 4390 15592
rect 4332 15583 4390 15589
rect 4798 15580 4804 15592
rect 4856 15580 4862 15632
rect 7668 15620 7696 15660
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7800 15660 7849 15688
rect 7800 15648 7806 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 10008 15660 10057 15688
rect 10008 15648 10014 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 10192 15660 13001 15688
rect 10192 15648 10198 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 10413 15623 10471 15629
rect 10413 15620 10425 15623
rect 5920 15592 6868 15620
rect 7668 15592 10425 15620
rect 2222 15552 2228 15564
rect 2183 15524 2228 15552
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 4028 15524 4077 15552
rect 4028 15512 4034 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 5920 15552 5948 15592
rect 4065 15515 4123 15521
rect 4172 15524 5948 15552
rect 6181 15555 6239 15561
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2516 15348 2544 15447
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 4172 15484 4200 15524
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6730 15552 6736 15564
rect 6227 15524 6736 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 6840 15552 6868 15592
rect 10413 15589 10425 15592
rect 10459 15620 10471 15623
rect 10686 15620 10692 15632
rect 10459 15592 10692 15620
rect 10459 15589 10471 15592
rect 10413 15583 10471 15589
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 8202 15552 8208 15564
rect 6840 15524 8208 15552
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 9214 15552 9220 15564
rect 8343 15524 9220 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 2924 15456 4200 15484
rect 2924 15444 2930 15456
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 6825 15487 6883 15493
rect 5500 15456 6500 15484
rect 5500 15444 5506 15456
rect 5258 15376 5264 15428
rect 5316 15416 5322 15428
rect 6472 15416 6500 15456
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15484 7803 15487
rect 8312 15484 8340 15515
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 11882 15561 11888 15564
rect 11876 15552 11888 15561
rect 10704 15524 11888 15552
rect 7791 15456 8340 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 6840 15416 6868 15447
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 10704 15493 10732 15524
rect 11876 15515 11888 15524
rect 11882 15512 11888 15515
rect 11940 15512 11946 15564
rect 10505 15487 10563 15493
rect 8444 15456 8489 15484
rect 8444 15444 8450 15456
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 5316 15388 6132 15416
rect 6472 15388 6868 15416
rect 5316 15376 5322 15388
rect 5534 15348 5540 15360
rect 2516 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6104 15348 6132 15388
rect 8846 15348 8852 15360
rect 6104 15320 8852 15348
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 9861 15351 9919 15357
rect 9861 15348 9873 15351
rect 9824 15320 9873 15348
rect 9824 15308 9830 15320
rect 9861 15317 9873 15320
rect 9907 15348 9919 15351
rect 10520 15348 10548 15447
rect 10594 15376 10600 15428
rect 10652 15416 10658 15428
rect 11238 15416 11244 15428
rect 10652 15388 11244 15416
rect 10652 15376 10658 15388
rect 11238 15376 11244 15388
rect 11296 15416 11302 15428
rect 11624 15416 11652 15447
rect 11296 15388 11652 15416
rect 11296 15376 11302 15388
rect 9907 15320 10548 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 7009 15147 7067 15153
rect 7009 15144 7021 15147
rect 4120 15116 7021 15144
rect 4120 15104 4126 15116
rect 7009 15113 7021 15116
rect 7055 15113 7067 15147
rect 7009 15107 7067 15113
rect 9953 15147 10011 15153
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10042 15144 10048 15156
rect 9999 15116 10048 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11296 15116 11621 15144
rect 11296 15104 11302 15116
rect 11609 15113 11621 15116
rect 11655 15113 11667 15147
rect 11609 15107 11667 15113
rect 3970 15036 3976 15088
rect 4028 15076 4034 15088
rect 4338 15076 4344 15088
rect 4028 15048 4344 15076
rect 4028 15036 4034 15048
rect 4338 15036 4344 15048
rect 4396 15036 4402 15088
rect 4890 15036 4896 15088
rect 4948 15036 4954 15088
rect 5166 15076 5172 15088
rect 5127 15048 5172 15076
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 11624 15076 11652 15107
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 11940 15116 13829 15144
rect 11940 15104 11946 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 12434 15076 12440 15088
rect 5736 15048 7880 15076
rect 11624 15048 12440 15076
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4706 15008 4712 15020
rect 4111 14980 4712 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 4908 15008 4936 15036
rect 5736 15008 5764 15048
rect 4908 14980 5764 15008
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 7006 15008 7012 15020
rect 5859 14980 7012 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 1670 14940 1676 14952
rect 1631 14912 1676 14940
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 2648 14912 3924 14940
rect 2648 14900 2654 14912
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 3418 14872 3424 14884
rect 1995 14844 3424 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 3418 14832 3424 14844
rect 3476 14832 3482 14884
rect 3786 14872 3792 14884
rect 3747 14844 3792 14872
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 3896 14872 3924 14912
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 5592 14912 6837 14940
rect 5592 14900 5598 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7374 14900 7380 14952
rect 7432 14940 7438 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 7432 14912 7757 14940
rect 7432 14900 7438 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 7852 14940 7880 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 8754 15008 8760 15020
rect 8715 14980 8760 15008
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 7852 14912 8585 14940
rect 7745 14903 7803 14909
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 5629 14875 5687 14881
rect 5629 14872 5641 14875
rect 3896 14844 5641 14872
rect 5629 14841 5641 14844
rect 5675 14841 5687 14875
rect 5629 14835 5687 14841
rect 8113 14875 8171 14881
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 10612 14872 10640 14971
rect 11790 14940 11796 14952
rect 11751 14912 11796 14940
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12492 14912 12537 14940
rect 12492 14900 12498 14912
rect 12342 14872 12348 14884
rect 8159 14844 8708 14872
rect 10612 14844 12348 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 8680 14816 8708 14844
rect 12342 14832 12348 14844
rect 12400 14872 12406 14884
rect 12682 14875 12740 14881
rect 12682 14872 12694 14875
rect 12400 14844 12694 14872
rect 12400 14832 12406 14844
rect 12682 14841 12694 14844
rect 12728 14841 12740 14875
rect 12682 14835 12740 14841
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 4890 14804 4896 14816
rect 4488 14776 4896 14804
rect 4488 14764 4494 14776
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 7282 14804 7288 14816
rect 5583 14776 7288 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7558 14804 7564 14816
rect 7519 14776 7564 14804
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8662 14804 8668 14816
rect 8623 14776 8668 14804
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 10318 14804 10324 14816
rect 10279 14776 10324 14804
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10468 14776 10513 14804
rect 10468 14764 10474 14776
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4028 14572 4660 14600
rect 4028 14560 4034 14572
rect 1397 14535 1455 14541
rect 1397 14501 1409 14535
rect 1443 14532 1455 14535
rect 4246 14532 4252 14544
rect 1443 14504 4252 14532
rect 1443 14501 1455 14504
rect 1397 14495 1455 14501
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 4430 14532 4436 14544
rect 4391 14504 4436 14532
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 1544 14436 2789 14464
rect 1544 14424 1550 14436
rect 2777 14433 2789 14436
rect 2823 14433 2835 14467
rect 2777 14427 2835 14433
rect 2866 14396 2872 14408
rect 2827 14368 2872 14396
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 4632 14405 4660 14572
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 4764 14572 7021 14600
rect 4764 14560 4770 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7800 14572 7849 14600
rect 7800 14560 7806 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 7837 14563 7895 14569
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 8260 14572 8309 14600
rect 8260 14560 8266 14572
rect 8297 14569 8309 14572
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 8536 14572 9873 14600
rect 8536 14560 8542 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12400 14572 12449 14600
rect 12400 14560 12406 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 5810 14492 5816 14544
rect 5868 14541 5874 14544
rect 5868 14535 5932 14541
rect 5868 14501 5886 14535
rect 5920 14501 5932 14535
rect 5868 14495 5932 14501
rect 5868 14492 5874 14495
rect 11238 14492 11244 14544
rect 11296 14492 11302 14544
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 7558 14464 7564 14476
rect 5675 14436 7564 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 11256 14464 11284 14492
rect 11103 14436 11284 14464
rect 11324 14467 11382 14473
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 11324 14433 11336 14467
rect 11370 14464 11382 14467
rect 11698 14464 11704 14476
rect 11370 14436 11704 14464
rect 11370 14433 11382 14436
rect 11324 14427 11382 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 1762 14288 1768 14340
rect 1820 14328 1826 14340
rect 2976 14328 3004 14359
rect 1820 14300 3004 14328
rect 1820 14288 1826 14300
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 2924 14232 4077 14260
rect 2924 14220 2930 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 4540 14260 4568 14359
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 7800 14368 8401 14396
rect 7800 14356 7806 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7190 14328 7196 14340
rect 6788 14300 7196 14328
rect 6788 14288 6794 14300
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 8478 14328 8484 14340
rect 7760 14300 8484 14328
rect 4985 14263 5043 14269
rect 4985 14260 4997 14263
rect 4540 14232 4997 14260
rect 4065 14223 4123 14229
rect 4985 14229 4997 14232
rect 5031 14260 5043 14263
rect 5258 14260 5264 14272
rect 5031 14232 5264 14260
rect 5031 14229 5043 14232
rect 4985 14223 5043 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 7760 14260 7788 14300
rect 8478 14288 8484 14300
rect 8536 14288 8542 14340
rect 5592 14232 7788 14260
rect 5592 14220 5598 14232
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 3936 14028 5181 14056
rect 3936 14016 3942 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 7800 14028 9229 14056
rect 7800 14016 7806 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 10045 14059 10103 14065
rect 10045 14025 10057 14059
rect 10091 14056 10103 14059
rect 10410 14056 10416 14068
rect 10091 14028 10416 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 2498 13988 2504 14000
rect 1627 13960 2504 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 2498 13948 2504 13960
rect 2556 13948 2562 14000
rect 7374 13988 7380 14000
rect 4724 13960 7380 13988
rect 1762 13880 1768 13932
rect 1820 13920 1826 13932
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 1820 13892 2145 13920
rect 1820 13880 1826 13892
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 2133 13883 2191 13889
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3384 13892 3801 13920
rect 3384 13880 3390 13892
rect 3789 13889 3801 13892
rect 3835 13920 3847 13923
rect 3970 13920 3976 13932
rect 3835 13892 3976 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 3050 13852 3056 13864
rect 2087 13824 3056 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4724 13861 4752 13960
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 5534 13920 5540 13932
rect 4816 13892 5540 13920
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 4709 13855 4767 13861
rect 3651 13824 4660 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 4632 13784 4660 13824
rect 4709 13821 4721 13855
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 4816 13784 4844 13892
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5810 13920 5816 13932
rect 5771 13892 5816 13920
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 11698 13920 11704 13932
rect 10735 13892 11704 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5123 13824 5641 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 5718 13852 5724 13864
rect 5675 13824 5724 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 7837 13855 7895 13861
rect 7837 13852 7849 13855
rect 6748 13824 7849 13852
rect 6748 13784 6776 13824
rect 7837 13821 7849 13824
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 8104 13855 8162 13861
rect 8104 13821 8116 13855
rect 8150 13852 8162 13855
rect 9953 13855 10011 13861
rect 8150 13824 8800 13852
rect 8150 13821 8162 13824
rect 8104 13815 8162 13821
rect 8772 13796 8800 13824
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10594 13852 10600 13864
rect 9999 13824 10600 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 4632 13756 4844 13784
rect 5460 13756 6776 13784
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 3142 13716 3148 13728
rect 3103 13688 3148 13716
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3292 13688 3525 13716
rect 3292 13676 3298 13688
rect 3513 13685 3525 13688
rect 3559 13685 3571 13719
rect 3513 13679 3571 13685
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 4525 13719 4583 13725
rect 4525 13716 4537 13719
rect 4396 13688 4537 13716
rect 4396 13676 4402 13688
rect 4525 13685 4537 13688
rect 4571 13716 4583 13719
rect 5460 13716 5488 13756
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7340 13756 8708 13784
rect 7340 13744 7346 13756
rect 4571 13688 5488 13716
rect 5537 13719 5595 13725
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 5626 13716 5632 13728
rect 5583 13688 5632 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13716 6883 13719
rect 8386 13716 8392 13728
rect 6871 13688 8392 13716
rect 6871 13685 6883 13688
rect 6825 13679 6883 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 8680 13716 8708 13756
rect 8754 13744 8760 13796
rect 8812 13744 8818 13796
rect 12437 13787 12495 13793
rect 12437 13784 12449 13787
rect 8956 13756 12449 13784
rect 8956 13716 8984 13756
rect 12437 13753 12449 13756
rect 12483 13753 12495 13787
rect 12437 13747 12495 13753
rect 10410 13716 10416 13728
rect 8680 13688 8984 13716
rect 10371 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10594 13716 10600 13728
rect 10551 13688 10600 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2280 13484 2421 13512
rect 2280 13472 2286 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 3142 13512 3148 13524
rect 2823 13484 3148 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4212 13484 4261 13512
rect 4212 13472 4218 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4249 13475 4307 13481
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 5868 13484 6653 13512
rect 5868 13472 5874 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 7432 13484 7481 13512
rect 7432 13472 7438 13484
rect 7469 13481 7481 13484
rect 7515 13481 7527 13515
rect 7469 13475 7527 13481
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8202 13512 8208 13524
rect 8067 13484 8208 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 10318 13512 10324 13524
rect 8536 13484 8581 13512
rect 10279 13484 10324 13512
rect 8536 13472 8542 13484
rect 10318 13472 10324 13484
rect 10376 13472 10382 13524
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 11756 13484 12725 13512
rect 11756 13472 11762 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 2866 13444 2872 13456
rect 2827 13416 2872 13444
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 5626 13444 5632 13456
rect 3476 13416 4108 13444
rect 3476 13404 3482 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 3786 13376 3792 13388
rect 1443 13348 3792 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 4080 13385 4108 13416
rect 4264 13416 5632 13444
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3970 13308 3976 13320
rect 3099 13280 3976 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 2958 13200 2964 13252
rect 3016 13240 3022 13252
rect 4264 13240 4292 13416
rect 5626 13404 5632 13416
rect 5684 13444 5690 13456
rect 10410 13444 10416 13456
rect 5684 13416 10416 13444
rect 5684 13404 5690 13416
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 4396 13348 5273 13376
rect 4396 13336 4402 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 5261 13339 5319 13345
rect 5528 13379 5586 13385
rect 5528 13345 5540 13379
rect 5574 13376 5586 13379
rect 7006 13376 7012 13388
rect 5574 13348 7012 13376
rect 5574 13345 5586 13348
rect 5528 13339 5586 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7650 13376 7656 13388
rect 7611 13348 7656 13376
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11589 13379 11647 13385
rect 11589 13376 11601 13379
rect 11204 13348 11601 13376
rect 11204 13336 11210 13348
rect 11589 13345 11601 13348
rect 11635 13345 11647 13379
rect 11589 13339 11647 13345
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8754 13308 8760 13320
rect 8711 13280 8760 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11296 13280 11345 13308
rect 11296 13268 11302 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 3016 13212 4292 13240
rect 3016 13200 3022 13212
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 6270 13172 6276 13184
rect 3568 13144 6276 13172
rect 3568 13132 3574 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 1673 12971 1731 12977
rect 1673 12968 1685 12971
rect 1636 12940 1685 12968
rect 1636 12928 1642 12940
rect 1673 12937 1685 12940
rect 1719 12937 1731 12971
rect 3970 12968 3976 12980
rect 3931 12940 3976 12968
rect 1673 12931 1731 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 10502 12968 10508 12980
rect 10463 12940 10508 12968
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 11848 12940 12081 12968
rect 11848 12928 11854 12940
rect 12069 12937 12081 12940
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 4856 12804 5733 12832
rect 4856 12792 4862 12804
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 5721 12795 5779 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12733 1547 12767
rect 1489 12727 1547 12733
rect 1504 12696 1532 12727
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2096 12736 2605 12764
rect 2096 12724 2102 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 4430 12764 4436 12776
rect 2593 12727 2651 12733
rect 2700 12736 4436 12764
rect 2700 12696 2728 12736
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7616 12736 7757 12764
rect 7616 12724 7622 12736
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 1504 12668 2728 12696
rect 2860 12699 2918 12705
rect 2860 12665 2872 12699
rect 2906 12696 2918 12699
rect 3326 12696 3332 12708
rect 2906 12668 3332 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 5537 12699 5595 12705
rect 5537 12665 5549 12699
rect 5583 12696 5595 12699
rect 6546 12696 6552 12708
rect 5583 12668 6552 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 7760 12696 7788 12727
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8001 12767 8059 12773
rect 8001 12764 8013 12767
rect 7892 12736 8013 12764
rect 7892 12724 7898 12736
rect 8001 12733 8013 12736
rect 8047 12733 8059 12767
rect 12250 12764 12256 12776
rect 12211 12736 12256 12764
rect 8001 12727 8059 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 8202 12696 8208 12708
rect 7760 12668 8208 12696
rect 8202 12656 8208 12668
rect 8260 12696 8266 12708
rect 9582 12696 9588 12708
rect 8260 12668 9588 12696
rect 8260 12656 8266 12668
rect 9582 12656 9588 12668
rect 9640 12696 9646 12708
rect 9674 12696 9680 12708
rect 9640 12668 9680 12696
rect 9640 12656 9646 12668
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10873 12699 10931 12705
rect 10873 12665 10885 12699
rect 10919 12696 10931 12699
rect 12437 12699 12495 12705
rect 12437 12696 12449 12699
rect 10919 12668 12449 12696
rect 10919 12665 10931 12668
rect 10873 12659 10931 12665
rect 12437 12665 12449 12668
rect 12483 12665 12495 12699
rect 12437 12659 12495 12665
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 9122 12628 9128 12640
rect 5684 12600 5729 12628
rect 9083 12600 9128 12628
rect 5684 12588 5690 12600
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 11020 12600 11065 12628
rect 11020 12588 11026 12600
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 3234 12424 3240 12436
rect 1443 12396 3240 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7432 12396 7849 12424
rect 7432 12384 7438 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12393 11115 12427
rect 11057 12387 11115 12393
rect 4341 12359 4399 12365
rect 4341 12325 4353 12359
rect 4387 12356 4399 12359
rect 4430 12356 4436 12368
rect 4387 12328 4436 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 11072 12356 11100 12387
rect 11238 12356 11244 12368
rect 11072 12328 11244 12356
rect 11238 12316 11244 12328
rect 11296 12356 11302 12368
rect 12130 12359 12188 12365
rect 12130 12356 12142 12359
rect 11296 12328 12142 12356
rect 11296 12316 11302 12328
rect 12130 12325 12142 12328
rect 12176 12325 12188 12359
rect 12130 12319 12188 12325
rect 2774 12288 2780 12300
rect 2735 12260 2780 12288
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4154 12288 4160 12300
rect 4111 12260 4160 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 4304 12260 5549 12288
rect 4304 12248 4310 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5793 12291 5851 12297
rect 5793 12288 5805 12291
rect 5537 12251 5595 12257
rect 5644 12260 5805 12288
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 5644 12220 5672 12260
rect 5793 12257 5805 12260
rect 5839 12288 5851 12291
rect 6914 12288 6920 12300
rect 5839 12260 6920 12288
rect 5839 12257 5851 12260
rect 5793 12251 5851 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 9490 12288 9496 12300
rect 8251 12260 9496 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 9933 12291 9991 12297
rect 9933 12288 9945 12291
rect 9784 12260 9945 12288
rect 8294 12220 8300 12232
rect 3099 12192 5672 12220
rect 8255 12192 8300 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 2590 12152 2596 12164
rect 2455 12124 2596 12152
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 2590 12112 2596 12124
rect 2648 12112 2654 12164
rect 2884 12152 2912 12183
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12220 8539 12223
rect 9784 12220 9812 12260
rect 9933 12257 9945 12260
rect 9979 12257 9991 12291
rect 9933 12251 9991 12257
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11756 12260 11897 12288
rect 11756 12248 11762 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 11885 12251 11943 12257
rect 11992 12260 19717 12288
rect 11992 12220 12020 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 8527 12192 9812 12220
rect 10704 12192 12020 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 9692 12164 9720 12192
rect 5534 12152 5540 12164
rect 2884 12124 5540 12152
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 9674 12112 9680 12164
rect 9732 12112 9738 12164
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 10704 12084 10732 12192
rect 3476 12056 10732 12084
rect 3476 12044 3482 12056
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 11204 12056 13277 12084
rect 11204 12044 11210 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20622 12084 20628 12096
rect 19935 12056 20628 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 3326 11880 3332 11892
rect 3287 11852 3332 11880
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6328 11852 7021 11880
rect 6328 11840 6334 11852
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 7009 11843 7067 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 10962 11880 10968 11892
rect 10735 11852 10968 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12894 11880 12900 11892
rect 12124 11852 12900 11880
rect 12124 11840 12130 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8260 11716 8309 11744
rect 8260 11704 8266 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 9456 11716 10425 11744
rect 9456 11704 9462 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 10413 11707 10471 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2038 11676 2044 11688
rect 1995 11648 2044 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2038 11636 2044 11648
rect 2096 11676 2102 11688
rect 4338 11676 4344 11688
rect 2096 11648 4344 11676
rect 2096 11636 2102 11648
rect 4338 11636 4344 11648
rect 4396 11676 4402 11688
rect 4798 11685 4804 11688
rect 4525 11679 4583 11685
rect 4525 11676 4537 11679
rect 4396 11648 4537 11676
rect 4396 11636 4402 11648
rect 4525 11645 4537 11648
rect 4571 11645 4583 11679
rect 4792 11676 4804 11685
rect 4759 11648 4804 11676
rect 4525 11639 4583 11645
rect 4792 11639 4804 11648
rect 4798 11636 4804 11639
rect 4856 11636 4862 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5810 11676 5816 11688
rect 5592 11648 5816 11676
rect 5592 11636 5598 11648
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7098 11676 7104 11688
rect 6871 11648 7104 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 8570 11685 8576 11688
rect 8564 11676 8576 11685
rect 8483 11648 8576 11676
rect 8564 11639 8576 11648
rect 8628 11676 8634 11688
rect 9122 11676 9128 11688
rect 8628 11648 9128 11676
rect 8570 11636 8576 11639
rect 8628 11636 8634 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 11054 11676 11060 11688
rect 9232 11648 11060 11676
rect 2216 11611 2274 11617
rect 2216 11577 2228 11611
rect 2262 11608 2274 11611
rect 2590 11608 2596 11620
rect 2262 11580 2596 11608
rect 2262 11577 2274 11580
rect 2216 11571 2274 11577
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 9232 11608 9260 11648
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 11204 11648 19625 11676
rect 11204 11636 11210 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 2832 11580 9260 11608
rect 2832 11568 2838 11580
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6546 11500 6552 11552
rect 6604 11540 6610 11552
rect 8386 11540 8392 11552
rect 6604 11512 8392 11540
rect 6604 11500 6610 11512
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 10042 11540 10048 11552
rect 8812 11512 10048 11540
rect 8812 11500 8818 11512
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10226 11540 10232 11552
rect 10187 11512 10232 11540
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10594 11540 10600 11552
rect 10367 11512 10600 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 13262 11540 13268 11552
rect 11204 11512 11249 11540
rect 13223 11512 13268 11540
rect 11204 11500 11210 11512
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 20438 11540 20444 11552
rect 19843 11512 20444 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2372 11308 2421 11336
rect 2372 11296 2378 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 6822 11336 6828 11348
rect 2823 11308 6828 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 8021 11339 8079 11345
rect 6972 11308 7017 11336
rect 6972 11296 6978 11308
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8294 11336 8300 11348
rect 8067 11308 8300 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8444 11308 8489 11336
rect 8444 11296 8450 11308
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 9548 11308 12265 11336
rect 9548 11296 9554 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 5782 11271 5840 11277
rect 5782 11268 5794 11271
rect 3068 11240 5794 11268
rect 3068 11141 3096 11240
rect 5782 11237 5794 11240
rect 5828 11268 5840 11271
rect 5902 11268 5908 11280
rect 5828 11240 5908 11268
rect 5828 11237 5840 11240
rect 5782 11231 5840 11237
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 5994 11228 6000 11280
rect 6052 11268 6058 11280
rect 6052 11240 19104 11268
rect 6052 11228 6058 11240
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3476 11172 4077 11200
rect 3476 11160 3482 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4430 11200 4436 11212
rect 4387 11172 4436 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11200 7987 11203
rect 8481 11203 8539 11209
rect 7975 11172 8340 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 2884 11064 2912 11095
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 4982 11132 4988 11144
rect 3568 11104 4988 11132
rect 3568 11092 3574 11104
rect 4982 11092 4988 11104
rect 5040 11132 5046 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5040 11104 5549 11132
rect 5040 11092 5046 11104
rect 5537 11101 5549 11104
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5166 11064 5172 11076
rect 2884 11036 5172 11064
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 7650 11064 7656 11076
rect 7432 11036 7656 11064
rect 7432 11024 7438 11036
rect 7650 11024 7656 11036
rect 7708 11064 7714 11076
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 7708 11036 7757 11064
rect 7708 11024 7714 11036
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 8312 11064 8340 11172
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9214 11200 9220 11212
rect 8527 11172 9220 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10870 11200 10876 11212
rect 10459 11172 10876 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 12342 11200 12348 11212
rect 11756 11172 12348 11200
rect 11756 11160 11762 11172
rect 12342 11160 12348 11172
rect 12400 11200 12406 11212
rect 12802 11209 12808 11212
rect 12529 11203 12587 11209
rect 12529 11200 12541 11203
rect 12400 11172 12541 11200
rect 12400 11160 12406 11172
rect 12529 11169 12541 11172
rect 12575 11169 12587 11203
rect 12796 11200 12808 11209
rect 12763 11172 12808 11200
rect 12529 11163 12587 11169
rect 12796 11163 12808 11172
rect 12802 11160 12808 11163
rect 12860 11160 12866 11212
rect 19076 11209 19104 11240
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11169 19119 11203
rect 19061 11163 19119 11169
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 15838 11132 15844 11144
rect 8628 11104 8673 11132
rect 15799 11104 15844 11132
rect 8628 11092 8634 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 11698 11064 11704 11076
rect 8312 11036 11704 11064
rect 7745 11027 7803 11033
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 19245 11067 19303 11073
rect 13740 11036 14044 11064
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 13740 10996 13768 11036
rect 13906 10996 13912 11008
rect 3752 10968 13768 10996
rect 13867 10968 13912 10996
rect 3752 10956 3758 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14016 10996 14044 11036
rect 19245 11033 19257 11067
rect 19291 11064 19303 11067
rect 19978 11064 19984 11076
rect 19291 11036 19984 11064
rect 19291 11033 19303 11036
rect 19245 11027 19303 11033
rect 19978 11024 19984 11036
rect 20036 11024 20042 11076
rect 17402 10996 17408 11008
rect 14016 10968 17408 10996
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1728 10764 2053 10792
rect 1728 10752 1734 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4028 10764 4568 10792
rect 4028 10752 4034 10764
rect 4540 10724 4568 10764
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4856 10764 4997 10792
rect 4856 10752 4862 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 10137 10795 10195 10801
rect 4985 10755 5043 10761
rect 5092 10764 9996 10792
rect 5092 10724 5120 10764
rect 4540 10696 5120 10724
rect 8205 10727 8263 10733
rect 8205 10693 8217 10727
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 2590 10656 2596 10668
rect 2551 10628 2596 10656
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3568 10628 3617 10656
rect 3568 10616 3574 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 3605 10619 3663 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 3878 10597 3884 10600
rect 2556 10560 2601 10588
rect 2556 10548 2562 10560
rect 3872 10551 3884 10597
rect 3936 10588 3942 10600
rect 6917 10591 6975 10597
rect 3936 10560 3972 10588
rect 3878 10548 3884 10551
rect 3936 10548 3942 10560
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 8220 10588 8248 10687
rect 8846 10656 8852 10668
rect 8807 10628 8852 10656
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 6963 10560 8248 10588
rect 8665 10591 8723 10597
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9858 10588 9864 10600
rect 8711 10560 9864 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 9968 10588 9996 10764
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10226 10792 10232 10804
rect 10183 10764 10232 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12250 10792 12256 10804
rect 12115 10764 12256 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 13814 10724 13820 10736
rect 13775 10696 13820 10724
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14645 10727 14703 10733
rect 14645 10693 14657 10727
rect 14691 10724 14703 10727
rect 16022 10724 16028 10736
rect 14691 10696 16028 10724
rect 14691 10693 14703 10696
rect 14645 10687 14703 10693
rect 16022 10684 16028 10696
rect 16080 10684 16086 10736
rect 10778 10656 10784 10668
rect 10739 10628 10784 10656
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 10888 10628 12572 10656
rect 10888 10588 10916 10628
rect 9968 10560 10916 10588
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11756 10560 12265 10588
rect 11756 10548 11762 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 12400 10560 12449 10588
rect 12400 10548 12406 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12544 10588 12572 10628
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 14792 10628 15209 10656
rect 14792 10616 14798 10628
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 12544 10560 18521 10588
rect 12437 10551 12495 10557
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 12704 10523 12762 10529
rect 9732 10492 12173 10520
rect 9732 10480 9738 10492
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 10502 10452 10508 10464
rect 10463 10424 10508 10452
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10452 10655 10455
rect 11054 10452 11060 10464
rect 10643 10424 11060 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 11054 10412 11060 10424
rect 11112 10452 11118 10464
rect 11974 10452 11980 10464
rect 11112 10424 11980 10452
rect 11112 10412 11118 10424
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12145 10452 12173 10492
rect 12704 10489 12716 10523
rect 12750 10520 12762 10523
rect 13538 10520 13544 10532
rect 12750 10492 13544 10520
rect 12750 10489 12762 10492
rect 12704 10483 12762 10489
rect 13538 10480 13544 10492
rect 13596 10480 13602 10532
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 13648 10492 15025 10520
rect 13648 10452 13676 10492
rect 15013 10489 15025 10492
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 12145 10424 13676 10452
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 13780 10424 15117 10452
rect 13780 10412 13786 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 15105 10415 15163 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 18693 10455 18751 10461
rect 18693 10421 18705 10455
rect 18739 10452 18751 10455
rect 19426 10452 19432 10464
rect 18739 10424 19432 10452
rect 18739 10421 18751 10424
rect 18693 10415 18751 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2648 10220 2789 10248
rect 2648 10208 2654 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 4120 10220 4261 10248
rect 4120 10208 4126 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6880 10220 7021 10248
rect 6880 10208 6886 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8570 10248 8576 10260
rect 8067 10220 8576 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 11054 10248 11060 10260
rect 10551 10220 11060 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 11054 10208 11060 10220
rect 11112 10248 11118 10260
rect 12342 10248 12348 10260
rect 11112 10220 12348 10248
rect 11112 10208 11118 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 9950 10180 9956 10192
rect 8527 10152 9956 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 10778 10140 10784 10192
rect 10836 10189 10842 10192
rect 10836 10183 10900 10189
rect 10836 10149 10854 10183
rect 10888 10149 10900 10183
rect 10836 10143 10900 10149
rect 10836 10140 10842 10143
rect 1670 10121 1676 10124
rect 1664 10112 1676 10121
rect 1631 10084 1676 10112
rect 1664 10075 1676 10084
rect 1670 10072 1676 10075
rect 1728 10072 1734 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4246 10112 4252 10124
rect 4111 10084 4252 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10112 5871 10115
rect 6270 10112 6276 10124
rect 5859 10084 6276 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 9674 10112 9680 10124
rect 8435 10084 9680 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12492 10084 13277 10112
rect 12492 10072 12498 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 15556 10115 15614 10121
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 16114 10112 16120 10124
rect 15602 10084 16120 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 17494 10112 17500 10124
rect 17455 10084 17500 10112
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5132 10016 5917 10044
rect 5132 10004 5138 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6052 10016 6097 10044
rect 6052 10004 6058 10016
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8628 10016 8677 10044
rect 8628 10004 8634 10016
rect 8665 10013 8677 10016
rect 8711 10044 8723 10047
rect 9398 10044 9404 10056
rect 8711 10016 9404 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10551 10016 10609 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 10597 10007 10655 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 3786 9936 3792 9988
rect 3844 9976 3850 9988
rect 10410 9976 10416 9988
rect 3844 9948 10416 9976
rect 3844 9936 3850 9948
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 13556 9976 13584 10007
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15252 10016 15301 10044
rect 15252 10004 15258 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 18046 10044 18052 10056
rect 17819 10016 18052 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 12860 9948 13584 9976
rect 12860 9936 12866 9948
rect 5442 9908 5448 9920
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 9456 9880 11989 9908
rect 9456 9868 9462 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 12894 9908 12900 9920
rect 12855 9880 12900 9908
rect 11977 9871 12035 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13556 9908 13584 9948
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 13556 9880 16681 9908
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 1728 9676 2903 9704
rect 1728 9664 1734 9676
rect 2875 9636 2903 9676
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 5776 9676 6132 9704
rect 5776 9664 5782 9676
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2875 9608 3341 9636
rect 3329 9605 3341 9608
rect 3375 9605 3387 9639
rect 3329 9599 3387 9605
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4212 9608 4721 9636
rect 4212 9596 4218 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 4709 9599 4767 9605
rect 5350 9568 5356 9580
rect 5311 9540 5356 9568
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1452 9472 1961 9500
rect 1452 9460 1458 9472
rect 1949 9469 1961 9472
rect 1995 9500 2007 9503
rect 3510 9500 3516 9512
rect 1995 9472 3516 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5442 9500 5448 9512
rect 5123 9472 5448 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6104 9500 6132 9676
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 16172 9676 16221 9704
rect 16172 9664 16178 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 16209 9667 16267 9673
rect 10594 9636 10600 9648
rect 10555 9608 10600 9636
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 11882 9596 11888 9648
rect 11940 9596 11946 9648
rect 12066 9596 12072 9648
rect 12124 9636 12130 9648
rect 12158 9636 12164 9648
rect 12124 9608 12164 9636
rect 12124 9596 12130 9608
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19886 9636 19892 9648
rect 19484 9608 19892 9636
rect 19484 9596 19490 9608
rect 19886 9596 19892 9608
rect 19944 9596 19950 9648
rect 6472 9540 7604 9568
rect 6362 9500 6368 9512
rect 6104 9472 6368 9500
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 2216 9435 2274 9441
rect 2216 9401 2228 9435
rect 2262 9432 2274 9435
rect 2498 9432 2504 9444
rect 2262 9404 2504 9432
rect 2262 9401 2274 9404
rect 2216 9395 2274 9401
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 2866 9432 2872 9444
rect 2648 9404 2872 9432
rect 2648 9392 2654 9404
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 6472 9432 6500 9540
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7374 9500 7380 9512
rect 6687 9472 7380 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 7484 9432 7512 9463
rect 4948 9404 6500 9432
rect 7392 9404 7512 9432
rect 7576 9432 7604 9540
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10836 9540 11161 9568
rect 10836 9528 10842 9540
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11900 9568 11928 9596
rect 12342 9568 12348 9580
rect 11900 9540 12348 9568
rect 11149 9531 11207 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 12952 9540 13553 9568
rect 12952 9528 12958 9540
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 13906 9568 13912 9580
rect 13771 9540 13912 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 7736 9503 7794 9509
rect 7736 9469 7748 9503
rect 7782 9500 7794 9503
rect 8570 9500 8576 9512
rect 7782 9472 8576 9500
rect 7782 9469 7794 9472
rect 7736 9463 7794 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 11020 9472 11069 9500
rect 11020 9460 11026 9472
rect 11057 9469 11069 9472
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 14918 9500 14924 9512
rect 14875 9472 14924 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 15028 9472 18061 9500
rect 15028 9432 15056 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 7576 9404 11008 9432
rect 4948 9392 4954 9404
rect 7392 9376 7420 9404
rect 5166 9324 5172 9376
rect 5224 9364 5230 9376
rect 6454 9364 6460 9376
rect 5224 9336 5269 9364
rect 6415 9336 6460 9364
rect 5224 9324 5230 9336
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7374 9324 7380 9376
rect 7432 9324 7438 9376
rect 8846 9364 8852 9376
rect 8807 9336 8852 9364
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 10980 9373 11008 9404
rect 13096 9404 15056 9432
rect 15096 9435 15154 9441
rect 13096 9373 13124 9404
rect 15096 9401 15108 9435
rect 15142 9432 15154 9435
rect 16298 9432 16304 9444
rect 15142 9404 16304 9432
rect 15142 9401 15154 9404
rect 15096 9395 15154 9401
rect 10965 9367 11023 9373
rect 10965 9333 10977 9367
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 13081 9367 13139 9373
rect 13081 9333 13093 9367
rect 13127 9333 13139 9367
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13081 9327 13139 9333
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 15120 9364 15148 9395
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 18325 9435 18383 9441
rect 18325 9401 18337 9435
rect 18371 9432 18383 9435
rect 19610 9432 19616 9444
rect 18371 9404 19616 9432
rect 18371 9401 18383 9404
rect 18325 9395 18383 9401
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 14792 9336 15148 9364
rect 14792 9324 14798 9336
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1486 9160 1492 9172
rect 1443 9132 1492 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 4890 9160 4896 9172
rect 2823 9132 4896 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 5920 9132 8493 9160
rect 5160 9095 5218 9101
rect 5160 9061 5172 9095
rect 5206 9092 5218 9095
rect 5350 9092 5356 9104
rect 5206 9064 5356 9092
rect 5206 9061 5218 9064
rect 5160 9055 5218 9061
rect 5350 9052 5356 9064
rect 5408 9092 5414 9104
rect 5920 9092 5948 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 8481 9123 8539 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11054 9160 11060 9172
rect 10796 9132 11060 9160
rect 5408 9064 5948 9092
rect 5408 9052 5414 9064
rect 5994 9052 6000 9104
rect 6052 9092 6058 9104
rect 7346 9095 7404 9101
rect 7346 9092 7358 9095
rect 6052 9064 7358 9092
rect 6052 9052 6058 9064
rect 7346 9061 7358 9064
rect 7392 9061 7404 9095
rect 7346 9055 7404 9061
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 4338 9024 4344 9036
rect 2915 8996 4344 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 5534 9024 5540 9036
rect 4816 8996 5540 9024
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 4816 8956 4844 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 10796 9033 10824 9132
rect 11054 9120 11060 9132
rect 11112 9160 11118 9172
rect 11698 9160 11704 9172
rect 11112 9132 11704 9160
rect 11112 9120 11118 9132
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9129 13231 9163
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13173 9123 13231 9129
rect 13188 9092 13216 9123
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9129 15623 9163
rect 15565 9123 15623 9129
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16206 9160 16212 9172
rect 15979 9132 16212 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 14642 9092 14648 9104
rect 13188 9064 14648 9092
rect 14642 9052 14648 9064
rect 14700 9092 14706 9104
rect 15580 9092 15608 9123
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 16356 9132 18797 9160
rect 16356 9120 16362 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 18785 9123 18843 9129
rect 17494 9092 17500 9104
rect 14700 9064 15148 9092
rect 15580 9064 17500 9092
rect 14700 9052 14706 9064
rect 11054 9033 11060 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 11048 9024 11060 9033
rect 11015 8996 11060 9024
rect 10781 8987 10839 8993
rect 11048 8987 11060 8996
rect 11054 8984 11060 8987
rect 11112 8984 11118 9036
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 15120 9033 15148 9064
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 12308 8996 13369 9024
rect 12308 8984 12314 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 8993 15163 9027
rect 16022 9024 16028 9036
rect 15983 8996 16028 9024
rect 15105 8987 15163 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 17672 9027 17730 9033
rect 17672 8993 17684 9027
rect 17718 9024 17730 9027
rect 18874 9024 18880 9036
rect 17718 8996 18880 9024
rect 17718 8993 17730 8996
rect 17672 8987 17730 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 4897 8965 4903 8968
rect 3099 8928 4844 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 4893 8919 4903 8965
rect 4955 8956 4961 8968
rect 7101 8959 7159 8965
rect 4955 8928 4993 8956
rect 4897 8916 4903 8919
rect 4955 8916 4961 8928
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 3878 8820 3884 8832
rect 2455 8792 3884 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 6273 8823 6331 8829
rect 6273 8820 6285 8823
rect 4120 8792 6285 8820
rect 4120 8780 4126 8792
rect 6273 8789 6285 8792
rect 6319 8789 6331 8823
rect 7116 8820 7144 8919
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16172 8928 16217 8956
rect 16172 8916 16178 8928
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 16540 8928 17417 8956
rect 16540 8916 16546 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19613 8959 19671 8965
rect 19613 8956 19625 8959
rect 19392 8928 19625 8956
rect 19392 8916 19398 8928
rect 19613 8925 19625 8928
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 7374 8820 7380 8832
rect 7116 8792 7380 8820
rect 6273 8783 6331 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 9398 8820 9404 8832
rect 8536 8792 9404 8820
rect 8536 8780 8542 8792
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 12158 8820 12164 8832
rect 12119 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15194 8820 15200 8832
rect 14967 8792 15200 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 1946 8616 1952 8628
rect 1903 8588 1952 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 3108 8588 3433 8616
rect 3108 8576 3114 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5166 8616 5172 8628
rect 5123 8588 5172 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 5408 8588 9137 8616
rect 5408 8576 5414 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9950 8616 9956 8628
rect 9364 8588 9812 8616
rect 9911 8588 9956 8616
rect 9364 8576 9370 8588
rect 3602 8548 3608 8560
rect 2240 8520 3608 8548
rect 2240 8421 2268 8520
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 6546 8548 6552 8560
rect 3844 8520 6552 8548
rect 3844 8508 3850 8520
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 9784 8548 9812 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10410 8616 10416 8628
rect 10192 8588 10416 8616
rect 10192 8576 10198 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 14458 8616 14464 8628
rect 13188 8588 14464 8616
rect 9784 8520 10916 8548
rect 2498 8480 2504 8492
rect 2411 8452 2504 8480
rect 2498 8440 2504 8452
rect 2556 8480 2562 8492
rect 4062 8480 4068 8492
rect 2556 8452 4068 8480
rect 2556 8440 2562 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 5994 8480 6000 8492
rect 5767 8452 6000 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 10597 8483 10655 8489
rect 9456 8452 10364 8480
rect 9456 8440 9462 8452
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 2958 8412 2964 8424
rect 2363 8384 2964 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 3936 8384 5549 8412
rect 3936 8372 3942 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7432 8384 7757 8412
rect 7432 8372 7438 8384
rect 7745 8381 7757 8384
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 8012 8415 8070 8421
rect 8012 8381 8024 8415
rect 8058 8412 8070 8415
rect 8846 8412 8852 8424
rect 8058 8384 8852 8412
rect 8058 8381 8070 8384
rect 8012 8375 8070 8381
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 10336 8421 10364 8452
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10778 8480 10784 8492
rect 10643 8452 10784 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10888 8480 10916 8520
rect 13078 8480 13084 8492
rect 10888 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13188 8489 13216 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 17920 8588 19349 8616
rect 17920 8576 17926 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18598 8548 18604 8560
rect 18279 8520 18604 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8480 15807 8483
rect 20162 8480 20168 8492
rect 15795 8452 20168 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 10321 8415 10379 8421
rect 8996 8384 9536 8412
rect 8996 8372 9002 8384
rect 9508 8356 9536 8384
rect 10321 8381 10333 8415
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11848 8384 11897 8412
rect 11848 8372 11854 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 15344 8384 15485 8412
rect 15344 8372 15350 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 16758 8412 16764 8424
rect 16719 8384 16764 8412
rect 15473 8375 15531 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8412 19211 8415
rect 19518 8412 19524 8424
rect 19199 8384 19524 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 19518 8372 19524 8384
rect 19576 8372 19582 8424
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 3050 8344 3056 8356
rect 2832 8316 3056 8344
rect 2832 8304 2838 8316
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 4798 8344 4804 8356
rect 3896 8316 4804 8344
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 3896 8285 3924 8316
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5445 8347 5503 8353
rect 5445 8313 5457 8347
rect 5491 8344 5503 8347
rect 6822 8344 6828 8356
rect 5491 8316 6828 8344
rect 5491 8313 5503 8316
rect 5445 8307 5503 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 13446 8353 13452 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 9548 8316 10425 8344
rect 9548 8304 9554 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 13440 8344 13452 8353
rect 13407 8316 13452 8344
rect 10413 8307 10471 8313
rect 13440 8307 13452 8316
rect 13446 8304 13452 8307
rect 13504 8304 13510 8356
rect 19058 8304 19064 8356
rect 19116 8344 19122 8356
rect 20257 8347 20315 8353
rect 20257 8344 20269 8347
rect 19116 8316 20269 8344
rect 19116 8304 19122 8316
rect 20257 8313 20269 8316
rect 20303 8313 20315 8347
rect 20257 8307 20315 8313
rect 3881 8279 3939 8285
rect 3881 8245 3893 8279
rect 3927 8245 3939 8279
rect 3881 8239 3939 8245
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 9030 8276 9036 8288
rect 4120 8248 9036 8276
rect 4120 8236 4126 8248
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 14550 8276 14556 8288
rect 14511 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 16942 8276 16948 8288
rect 16903 8248 16948 8276
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 3418 8072 3424 8084
rect 2087 8044 3424 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4948 8044 4997 8072
rect 4948 8032 4954 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 4985 8035 5043 8041
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6052 8044 6653 8072
rect 6052 8032 6058 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 11238 8072 11244 8084
rect 6788 8044 11244 8072
rect 6788 8032 6794 8044
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 18874 8072 18880 8084
rect 11348 8044 16068 8072
rect 18835 8044 18880 8072
rect 6454 8004 6460 8016
rect 5184 7976 6460 8004
rect 2222 7896 2228 7948
rect 2280 7936 2286 7948
rect 5184 7945 5212 7976
rect 6454 7964 6460 7976
rect 6512 8004 6518 8016
rect 6512 7976 7696 8004
rect 6512 7964 6518 7976
rect 5534 7945 5540 7948
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 2280 7908 2421 7936
rect 2280 7896 2286 7908
rect 2409 7905 2421 7908
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5528 7936 5540 7945
rect 5447 7908 5540 7936
rect 5169 7899 5227 7905
rect 5528 7899 5540 7908
rect 5592 7936 5598 7948
rect 6730 7936 6736 7948
rect 5592 7908 6736 7936
rect 5534 7896 5540 7899
rect 5592 7896 5598 7908
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 7668 7945 7696 7976
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 11348 8004 11376 8044
rect 9640 7976 11376 8004
rect 9640 7964 9646 7976
rect 12158 7964 12164 8016
rect 12216 8013 12222 8016
rect 12216 8007 12280 8013
rect 12216 7973 12234 8007
rect 12268 7973 12280 8007
rect 12216 7967 12280 7973
rect 12216 7964 12222 7967
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 15534 8007 15592 8013
rect 15534 8004 15546 8007
rect 14608 7976 15546 8004
rect 14608 7964 14614 7976
rect 15534 7973 15546 7976
rect 15580 7973 15592 8007
rect 16040 8004 16068 8044
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 19794 8004 19800 8016
rect 16040 7976 19800 8004
rect 15534 7967 15592 7973
rect 19794 7964 19800 7976
rect 19852 7964 19858 8016
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 7800 7908 8401 7936
rect 7800 7896 7806 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 9944 7939 10002 7945
rect 9944 7905 9956 7939
rect 9990 7936 10002 7939
rect 10226 7936 10232 7948
rect 9990 7908 10232 7936
rect 9990 7905 10002 7908
rect 9944 7899 10002 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11756 7908 11989 7936
rect 11756 7896 11762 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 16482 7936 16488 7948
rect 11977 7899 12035 7905
rect 15304 7908 16488 7936
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 4246 7868 4252 7880
rect 2731 7840 4252 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 8478 7868 8484 7880
rect 8439 7840 8484 7868
rect 5261 7831 5319 7837
rect 5276 7732 5304 7831
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9677 7871 9735 7877
rect 8628 7840 8673 7868
rect 8628 7828 8634 7840
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 14182 7868 14188 7880
rect 14143 7840 14188 7868
rect 9677 7831 9735 7837
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 9122 7800 9128 7812
rect 8352 7772 9128 7800
rect 8352 7760 8358 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 7374 7732 7380 7744
rect 5276 7704 7380 7732
rect 7374 7692 7380 7704
rect 7432 7732 7438 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7432 7704 7481 7732
rect 7432 7692 7438 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7469 7695 7527 7701
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8386 7732 8392 7744
rect 8067 7704 8392 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9692 7732 9720 7831
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15304 7877 15332 7908
rect 16482 7896 16488 7908
rect 16540 7936 16546 7948
rect 17770 7945 17776 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 16540 7908 17509 7936
rect 16540 7896 16546 7908
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 17764 7899 17776 7945
rect 17828 7936 17834 7948
rect 17828 7908 17864 7936
rect 17770 7896 17776 7899
rect 17828 7896 17834 7908
rect 18782 7896 18788 7948
rect 18840 7936 18846 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 18840 7908 19717 7936
rect 18840 7896 18846 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15252 7840 15301 7868
rect 15252 7828 15258 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 10042 7732 10048 7744
rect 9692 7704 10048 7732
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 11054 7732 11060 7744
rect 10967 7704 11060 7732
rect 11054 7692 11060 7704
rect 11112 7732 11118 7744
rect 11882 7732 11888 7744
rect 11112 7704 11888 7732
rect 11112 7692 11118 7704
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 13357 7735 13415 7741
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13446 7732 13452 7744
rect 13403 7704 13452 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 16080 7704 16681 7732
rect 16080 7692 16086 7704
rect 16669 7701 16681 7704
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19024 7704 19901 7732
rect 19024 7692 19030 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 19889 7695 19947 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7742 7528 7748 7540
rect 6963 7500 7748 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 8128 7500 10701 7528
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 8128 7460 8156 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 10689 7491 10747 7497
rect 10796 7500 16865 7528
rect 6880 7432 8156 7460
rect 6880 7420 6886 7432
rect 10410 7420 10416 7472
rect 10468 7460 10474 7472
rect 10796 7460 10824 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 22278 7528 22284 7540
rect 20956 7500 22284 7528
rect 20956 7488 20962 7500
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 10468 7432 10824 7460
rect 10468 7420 10474 7432
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7156 7364 7481 7392
rect 7156 7352 7162 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 7469 7355 7527 7361
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12216 7364 13001 7392
rect 12216 7352 12222 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 18874 7392 18880 7404
rect 18739 7364 18880 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 1412 7324 1440 7352
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 1412 7296 3617 7324
rect 3605 7293 3617 7296
rect 3651 7324 3663 7327
rect 3694 7324 3700 7336
rect 3651 7296 3700 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6972 7296 7389 7324
rect 6972 7284 6978 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 8202 7324 8208 7336
rect 7616 7296 8208 7324
rect 7616 7284 7622 7296
rect 8202 7284 8208 7296
rect 8260 7324 8266 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8260 7296 8493 7324
rect 8260 7284 8266 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 12710 7324 12716 7336
rect 9088 7296 12716 7324
rect 9088 7284 9094 7296
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 12894 7324 12900 7336
rect 12807 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7324 12958 7336
rect 13722 7324 13728 7336
rect 12952 7296 13728 7324
rect 12952 7284 12958 7296
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 13998 7324 14004 7336
rect 13959 7296 14004 7324
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 14516 7296 15485 7324
rect 14516 7284 14522 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 15740 7327 15798 7333
rect 15740 7293 15752 7327
rect 15786 7324 15798 7327
rect 16022 7324 16028 7336
rect 15786 7296 16028 7324
rect 15786 7293 15798 7296
rect 15740 7287 15798 7293
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 19610 7324 19616 7336
rect 19571 7296 19616 7324
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 1670 7265 1676 7268
rect 1664 7256 1676 7265
rect 1631 7228 1676 7256
rect 1664 7219 1676 7228
rect 1670 7216 1676 7219
rect 1728 7216 1734 7268
rect 3850 7259 3908 7265
rect 3850 7256 3862 7259
rect 2792 7228 3862 7256
rect 2792 7200 2820 7228
rect 3850 7225 3862 7228
rect 3896 7225 3908 7259
rect 3850 7219 3908 7225
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 4120 7228 7512 7256
rect 4120 7216 4126 7228
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2832 7160 2925 7188
rect 2832 7148 2838 7160
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4304 7160 4997 7188
rect 4304 7148 4310 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 7064 7160 7297 7188
rect 7064 7148 7070 7160
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 7484 7188 7512 7228
rect 8662 7216 8668 7268
rect 8720 7265 8726 7268
rect 8720 7259 8784 7265
rect 8720 7225 8738 7259
rect 8772 7225 8784 7259
rect 13906 7256 13912 7268
rect 8720 7219 8784 7225
rect 8864 7228 13912 7256
rect 8720 7216 8726 7219
rect 8864 7188 8892 7228
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 14277 7259 14335 7265
rect 14277 7225 14289 7259
rect 14323 7256 14335 7259
rect 14366 7256 14372 7268
rect 14323 7228 14372 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 7484 7160 8892 7188
rect 9861 7191 9919 7197
rect 7285 7151 7343 7157
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10226 7188 10232 7200
rect 9907 7160 10232 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 10652 7160 11069 7188
rect 10652 7148 10658 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11974 7188 11980 7200
rect 11195 7160 11980 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 12805 7151 12863 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18414 7188 18420 7200
rect 18375 7160 18420 7188
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18506 7148 18512 7200
rect 18564 7188 18570 7200
rect 18564 7160 18609 7188
rect 18564 7148 18570 7160
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 19208 7160 19809 7188
rect 19208 7148 19214 7160
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2222 6984 2228 6996
rect 2183 6956 2228 6984
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 13262 6984 13268 6996
rect 4212 6956 9628 6984
rect 13223 6956 13268 6984
rect 4212 6944 4218 6956
rect 2593 6919 2651 6925
rect 2593 6885 2605 6919
rect 2639 6916 2651 6919
rect 3326 6916 3332 6928
rect 2639 6888 3332 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 4028 6888 4200 6916
rect 4028 6876 4034 6888
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3752 6820 4077 6848
rect 3752 6808 3758 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4172 6848 4200 6888
rect 4246 6876 4252 6928
rect 4304 6925 4310 6928
rect 4304 6919 4368 6925
rect 4304 6885 4322 6919
rect 4356 6885 4368 6919
rect 8846 6916 8852 6928
rect 4304 6879 4368 6885
rect 4448 6888 8852 6916
rect 4304 6876 4310 6879
rect 4448 6848 4476 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 6270 6848 6276 6860
rect 4172 6820 4476 6848
rect 6231 6820 6276 6848
rect 4065 6811 4123 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7466 6848 7472 6860
rect 7423 6820 7472 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7644 6851 7702 6857
rect 7644 6817 7656 6851
rect 7690 6848 7702 6851
rect 8570 6848 8576 6860
rect 7690 6820 8576 6848
rect 7690 6817 7702 6820
rect 7644 6811 7702 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9600 6848 9628 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 15657 6987 15715 6993
rect 15657 6953 15669 6987
rect 15703 6984 15715 6987
rect 15838 6984 15844 6996
rect 15703 6956 15844 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18564 6956 19257 6984
rect 18564 6944 18570 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19613 6987 19671 6993
rect 19613 6953 19625 6987
rect 19659 6984 19671 6987
rect 19794 6984 19800 6996
rect 19659 6956 19800 6984
rect 19659 6953 19671 6956
rect 19613 6947 19671 6953
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 11609 6919 11667 6925
rect 11609 6916 11621 6919
rect 9732 6888 11621 6916
rect 9732 6876 9738 6888
rect 11609 6885 11621 6888
rect 11655 6885 11667 6919
rect 11609 6879 11667 6885
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 13357 6919 13415 6925
rect 13357 6916 13369 6919
rect 12492 6888 13369 6916
rect 12492 6876 12498 6888
rect 13357 6885 13369 6888
rect 13403 6885 13415 6919
rect 13357 6879 13415 6885
rect 18049 6919 18107 6925
rect 18049 6885 18061 6919
rect 18095 6916 18107 6919
rect 19334 6916 19340 6928
rect 18095 6888 19340 6916
rect 18095 6885 18107 6888
rect 18049 6879 18107 6885
rect 19334 6876 19340 6888
rect 19392 6876 19398 6928
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9600 6820 10057 6848
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 14642 6848 14648 6860
rect 14603 6820 14648 6848
rect 10045 6811 10103 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17460 6820 17509 6848
rect 17460 6808 17466 6820
rect 17497 6817 17509 6820
rect 17543 6848 17555 6851
rect 18141 6851 18199 6857
rect 18141 6848 18153 6851
rect 17543 6820 18153 6848
rect 17543 6817 17555 6820
rect 17497 6811 17555 6817
rect 18141 6817 18153 6820
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19668 6820 19717 6848
rect 19668 6808 19674 6820
rect 19705 6817 19717 6820
rect 19751 6817 19763 6851
rect 19705 6811 19763 6817
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2648 6752 2697 6780
rect 2648 6740 2654 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 2832 6752 2877 6780
rect 2832 6740 2838 6752
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9916 6752 10149 6780
rect 9916 6740 9922 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 10284 6752 10329 6780
rect 10704 6752 11713 6780
rect 10284 6740 10290 6752
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 3878 6712 3884 6724
rect 1728 6684 3884 6712
rect 1728 6672 1734 6684
rect 3878 6672 3884 6684
rect 3936 6672 3942 6724
rect 9677 6715 9735 6721
rect 5000 6684 5580 6712
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5000 6644 5028 6684
rect 5442 6644 5448 6656
rect 4120 6616 5028 6644
rect 5403 6616 5448 6644
rect 4120 6604 4126 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5552 6644 5580 6684
rect 8312 6684 8892 6712
rect 8312 6644 8340 6684
rect 5552 6616 8340 6644
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8720 6616 8769 6644
rect 8720 6604 8726 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8864 6644 8892 6684
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 10704 6712 10732 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11882 6780 11888 6792
rect 11843 6752 11888 6780
rect 11701 6743 11759 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12618 6780 12624 6792
rect 11992 6752 12624 6780
rect 11992 6712 12020 6752
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13504 6752 13549 6780
rect 13504 6740 13510 6752
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 13872 6752 15761 6780
rect 13872 6740 13878 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17828 6752 18245 6780
rect 17828 6740 17834 6752
rect 18233 6749 18245 6752
rect 18279 6780 18291 6783
rect 19794 6780 19800 6792
rect 18279 6752 19800 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 9723 6684 10732 6712
rect 11164 6684 12020 6712
rect 12897 6715 12955 6721
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 11164 6644 11192 6684
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13998 6712 14004 6724
rect 12943 6684 14004 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14458 6712 14464 6724
rect 14419 6684 14464 6712
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 15286 6712 15292 6724
rect 15247 6684 15292 6712
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 17681 6715 17739 6721
rect 17681 6681 17693 6715
rect 17727 6712 17739 6715
rect 18414 6712 18420 6724
rect 17727 6684 18420 6712
rect 17727 6681 17739 6684
rect 17681 6675 17739 6681
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 8864 6616 11192 6644
rect 11241 6647 11299 6653
rect 8757 6607 8815 6613
rect 11241 6613 11253 6647
rect 11287 6644 11299 6647
rect 12526 6644 12532 6656
rect 11287 6616 12532 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 2498 6440 2504 6452
rect 1719 6412 2504 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5169 6443 5227 6449
rect 5169 6440 5181 6443
rect 5132 6412 5181 6440
rect 5132 6400 5138 6412
rect 5169 6409 5181 6412
rect 5215 6409 5227 6443
rect 8205 6443 8263 6449
rect 5169 6403 5227 6409
rect 5460 6412 8156 6440
rect 3237 6375 3295 6381
rect 3237 6372 3249 6375
rect 2056 6344 3249 6372
rect 2056 6245 2084 6344
rect 3237 6341 3249 6344
rect 3283 6341 3295 6375
rect 3237 6335 3295 6341
rect 3418 6332 3424 6384
rect 3476 6372 3482 6384
rect 5460 6372 5488 6412
rect 3476 6344 5488 6372
rect 8128 6372 8156 6412
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8570 6440 8576 6452
rect 8251 6412 8576 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 19794 6400 19800 6452
rect 19852 6440 19858 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 19852 6412 20453 6440
rect 19852 6400 19858 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 9490 6372 9496 6384
rect 8128 6344 9496 6372
rect 3476 6332 3482 6344
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2774 6304 2780 6316
rect 2363 6276 2780 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3694 6304 3700 6316
rect 3016 6276 3700 6304
rect 3016 6264 3022 6276
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 3878 6304 3884 6316
rect 3791 6276 3884 6304
rect 3878 6264 3884 6276
rect 3936 6304 3942 6316
rect 5350 6304 5356 6316
rect 3936 6276 5356 6304
rect 3936 6264 3942 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 3602 6236 3608 6248
rect 3563 6208 3608 6236
rect 2041 6199 2099 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 5460 6236 5488 6344
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 12308 6344 13400 6372
rect 12308 6332 12314 6344
rect 13372 6316 13400 6344
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5592 6276 5733 6304
rect 5592 6264 5598 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9674 6304 9680 6316
rect 9171 6276 9680 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10100 6276 10149 6304
rect 10100 6264 10106 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13412 6276 14289 6304
rect 13412 6264 13418 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 14550 6304 14556 6316
rect 14507 6276 14556 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16482 6304 16488 6316
rect 16347 6276 16488 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5460 6208 5641 6236
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6052 6208 6837 6236
rect 6052 6196 6058 6208
rect 6825 6205 6837 6208
rect 6871 6236 6883 6239
rect 7466 6236 7472 6248
rect 6871 6208 7472 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 10410 6245 10416 6248
rect 10393 6239 10416 6245
rect 10393 6205 10405 6239
rect 10393 6199 10416 6205
rect 10410 6196 10416 6199
rect 10468 6196 10474 6248
rect 12526 6236 12532 6248
rect 12487 6208 12532 6236
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13964 6208 14197 6236
rect 13964 6196 13970 6208
rect 14185 6205 14197 6208
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18196 6208 19073 6236
rect 18196 6196 18202 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 6914 6168 6920 6180
rect 3568 6140 6920 6168
rect 3568 6128 3574 6140
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7098 6177 7104 6180
rect 7092 6168 7104 6177
rect 7059 6140 7104 6168
rect 7092 6131 7104 6140
rect 7098 6128 7104 6131
rect 7156 6128 7162 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 14734 6168 14740 6180
rect 12851 6140 14740 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 19334 6177 19340 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 16071 6140 18061 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 18049 6137 18061 6140
rect 18095 6137 18107 6171
rect 19328 6168 19340 6177
rect 19295 6140 19340 6168
rect 18049 6131 18107 6137
rect 19328 6131 19340 6140
rect 19334 6128 19340 6131
rect 19392 6128 19398 6180
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 5534 6100 5540 6112
rect 4028 6072 5540 6100
rect 4028 6060 4034 6072
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 6932 6100 6960 6128
rect 11330 6100 11336 6112
rect 6932 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11514 6100 11520 6112
rect 11475 6072 11520 6100
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 12342 6100 12348 6112
rect 11756 6072 12348 6100
rect 11756 6060 11762 6072
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15746 6100 15752 6112
rect 15703 6072 15752 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2188 5868 4077 5896
rect 2188 5856 2194 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 8340 5896
rect 5592 5856 5598 5868
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 3786 5828 3792 5840
rect 2372 5800 3792 5828
rect 2372 5788 2378 5800
rect 3786 5788 3792 5800
rect 3844 5828 3850 5840
rect 4433 5831 4491 5837
rect 4433 5828 4445 5831
rect 3844 5800 4445 5828
rect 3844 5788 3850 5800
rect 4433 5797 4445 5800
rect 4479 5797 4491 5831
rect 5994 5828 6000 5840
rect 4433 5791 4491 5797
rect 5644 5800 6000 5828
rect 2682 5760 2688 5772
rect 2643 5732 2688 5760
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 5644 5769 5672 5800
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 8312 5828 8340 5868
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8444 5868 8493 5896
rect 8444 5856 8450 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 9398 5896 9404 5908
rect 8481 5859 8539 5865
rect 8772 5868 9404 5896
rect 8772 5828 8800 5868
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 9769 5899 9827 5905
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 11054 5896 11060 5908
rect 9815 5868 11060 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 13633 5899 13691 5905
rect 11388 5868 11744 5896
rect 11388 5856 11394 5868
rect 8312 5800 8800 5828
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 8904 5800 10149 5828
rect 8904 5788 8910 5800
rect 10137 5797 10149 5800
rect 10183 5797 10195 5831
rect 10137 5791 10195 5797
rect 11238 5788 11244 5840
rect 11296 5828 11302 5840
rect 11514 5828 11520 5840
rect 11296 5800 11520 5828
rect 11296 5788 11302 5800
rect 11514 5788 11520 5800
rect 11572 5837 11578 5840
rect 11572 5831 11636 5837
rect 11572 5797 11590 5831
rect 11624 5797 11636 5831
rect 11716 5828 11744 5868
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 16114 5896 16120 5908
rect 13679 5868 16120 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 11716 5800 14105 5828
rect 11572 5791 11636 5797
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 11572 5788 11578 5791
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 5896 5763 5954 5769
rect 5896 5729 5908 5763
rect 5942 5760 5954 5763
rect 6822 5760 6828 5772
rect 5942 5732 6828 5760
rect 5942 5729 5954 5732
rect 5896 5723 5954 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 6972 5732 8401 5760
rect 6972 5720 6978 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 8389 5723 8447 5729
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 10042 5760 10048 5772
rect 9732 5732 10048 5760
rect 9732 5720 9738 5732
rect 10042 5720 10048 5732
rect 10100 5760 10106 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10100 5732 11345 5760
rect 10100 5720 10106 5732
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 12342 5760 12348 5772
rect 11379 5732 12348 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 14001 5763 14059 5769
rect 14001 5760 14013 5763
rect 13136 5732 14013 5760
rect 13136 5720 13142 5732
rect 14001 5729 14013 5732
rect 14047 5729 14059 5763
rect 14918 5760 14924 5772
rect 14001 5723 14059 5729
rect 14292 5732 14924 5760
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 1912 5664 2789 5692
rect 1912 5652 1918 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2777 5655 2835 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3844 5664 4537 5692
rect 3844 5652 3850 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 5350 5692 5356 5704
rect 4755 5664 5356 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 10229 5695 10287 5701
rect 10229 5692 10241 5695
rect 8904 5664 10241 5692
rect 8904 5652 8910 5664
rect 10229 5661 10241 5664
rect 10275 5661 10287 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 10229 5655 10287 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 14292 5701 14320 5732
rect 14918 5720 14924 5732
rect 14976 5760 14982 5772
rect 18690 5769 18696 5772
rect 15545 5763 15603 5769
rect 15545 5760 15557 5763
rect 14976 5732 15557 5760
rect 14976 5720 14982 5732
rect 15545 5729 15557 5732
rect 15591 5729 15603 5763
rect 18684 5760 18696 5769
rect 18651 5732 18696 5760
rect 15545 5723 15603 5729
rect 18684 5723 18696 5732
rect 18690 5720 18696 5723
rect 18748 5720 18754 5772
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 14277 5655 14335 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18196 5664 18429 5692
rect 18196 5652 18202 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 5534 5624 5540 5636
rect 4120 5596 5540 5624
rect 4120 5584 4126 5596
rect 5534 5584 5540 5596
rect 5592 5584 5598 5636
rect 8021 5627 8079 5633
rect 8021 5593 8033 5627
rect 8067 5624 8079 5627
rect 8067 5596 10272 5624
rect 8067 5593 8079 5596
rect 8021 5587 8079 5593
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 4246 5556 4252 5568
rect 2363 5528 4252 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 7098 5556 7104 5568
rect 7055 5528 7104 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 7098 5516 7104 5528
rect 7156 5556 7162 5568
rect 8938 5556 8944 5568
rect 7156 5528 8944 5556
rect 7156 5516 7162 5528
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 10244 5556 10272 5596
rect 12526 5556 12532 5568
rect 10244 5528 12532 5556
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16540 5528 16681 5556
rect 16540 5516 16546 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19797 5559 19855 5565
rect 19797 5556 19809 5559
rect 19392 5528 19809 5556
rect 19392 5516 19398 5528
rect 19797 5525 19809 5528
rect 19843 5525 19855 5559
rect 19797 5519 19855 5525
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1765 5355 1823 5361
rect 1765 5321 1777 5355
rect 1811 5352 1823 5355
rect 2682 5352 2688 5364
rect 1811 5324 2688 5352
rect 1811 5321 1823 5324
rect 1765 5315 1823 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 6914 5352 6920 5364
rect 6871 5324 6920 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 8478 5352 8484 5364
rect 8435 5324 8484 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 12621 5355 12679 5361
rect 12621 5321 12633 5355
rect 12667 5352 12679 5355
rect 14642 5352 14648 5364
rect 12667 5324 14648 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 14918 5352 14924 5364
rect 14879 5324 14924 5352
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 4617 5287 4675 5293
rect 4617 5253 4629 5287
rect 4663 5284 4675 5287
rect 6638 5284 6644 5296
rect 4663 5256 6644 5284
rect 4663 5253 4675 5256
rect 4617 5247 4675 5253
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 13354 5284 13360 5296
rect 10827 5256 13360 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 13354 5244 13360 5256
rect 13412 5244 13418 5296
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2866 5216 2872 5228
rect 2455 5188 2872 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 3326 5216 3332 5228
rect 3287 5188 3332 5216
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4948 5188 5181 5216
rect 4948 5176 4954 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 5592 5188 7297 5216
rect 5592 5176 5598 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 8570 5216 8576 5228
rect 7515 5188 8576 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8938 5216 8944 5228
rect 8899 5188 8944 5216
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11296 5188 11345 5216
rect 11296 5176 11302 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 12894 5216 12900 5228
rect 11333 5179 11391 5185
rect 11440 5188 12900 5216
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 3936 5120 4997 5148
rect 3936 5108 3942 5120
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 8846 5148 8852 5160
rect 4985 5111 5043 5117
rect 8772 5120 8852 5148
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 4062 5080 4068 5092
rect 2179 5052 4068 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 7193 5083 7251 5089
rect 7193 5049 7205 5083
rect 7239 5080 7251 5083
rect 8386 5080 8392 5092
rect 7239 5052 8392 5080
rect 7239 5049 7251 5052
rect 7193 5043 7251 5049
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 8772 5089 8800 5120
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 11440 5148 11468 5188
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 9600 5120 11468 5148
rect 12437 5151 12495 5157
rect 8757 5083 8815 5089
rect 8757 5080 8769 5083
rect 8720 5052 8769 5080
rect 8720 5040 8726 5052
rect 8757 5049 8769 5052
rect 8803 5049 8815 5083
rect 9600 5080 9628 5120
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5148 13599 5151
rect 13587 5120 14504 5148
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 8757 5043 8815 5049
rect 8864 5052 9628 5080
rect 8864 5024 8892 5052
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 11112 5052 11253 5080
rect 11112 5040 11118 5052
rect 11241 5049 11253 5052
rect 11287 5049 11299 5083
rect 11241 5043 11299 5049
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3878 5012 3884 5024
rect 3476 4984 3884 5012
rect 3476 4972 3482 4984
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 5074 5012 5080 5024
rect 5035 4984 5080 5012
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 12452 5012 12480 5111
rect 14476 5092 14504 5120
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15344 5120 15761 5148
rect 15344 5108 15350 5120
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 15838 5148 15844 5160
rect 15795 5120 15844 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16016 5151 16074 5157
rect 16016 5117 16028 5151
rect 16062 5148 16074 5151
rect 16482 5148 16488 5160
rect 16062 5120 16488 5148
rect 16062 5117 16074 5120
rect 16016 5111 16074 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18138 5148 18144 5160
rect 18095 5120 18144 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 20254 5148 20260 5160
rect 20215 5120 20260 5148
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 13808 5083 13866 5089
rect 13808 5049 13820 5083
rect 13854 5080 13866 5083
rect 13906 5080 13912 5092
rect 13854 5052 13912 5080
rect 13854 5049 13866 5052
rect 13808 5043 13866 5049
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14458 5040 14464 5092
rect 14516 5040 14522 5092
rect 17770 5040 17776 5092
rect 17828 5080 17834 5092
rect 18294 5083 18352 5089
rect 18294 5080 18306 5083
rect 17828 5052 18306 5080
rect 17828 5040 17834 5052
rect 18294 5049 18306 5052
rect 18340 5049 18352 5083
rect 18294 5043 18352 5049
rect 18874 5040 18880 5092
rect 18932 5080 18938 5092
rect 18932 5052 20484 5080
rect 18932 5040 18938 5052
rect 14550 5012 14556 5024
rect 12452 4984 14556 5012
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 17126 5012 17132 5024
rect 17087 4984 17132 5012
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 18690 4972 18696 5024
rect 18748 5012 18754 5024
rect 20456 5021 20484 5052
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 18748 4984 19441 5012
rect 18748 4972 18754 4984
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 19429 4975 19487 4981
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 3016 4780 3157 4808
rect 3016 4768 3022 4780
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 4062 4808 4068 4820
rect 4023 4780 4068 4808
rect 3145 4771 3203 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 6822 4808 6828 4820
rect 6783 4780 6828 4808
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8846 4808 8852 4820
rect 8260 4780 8852 4808
rect 8260 4768 8266 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 13630 4808 13636 4820
rect 12492 4780 13636 4808
rect 12492 4768 12498 4780
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 19058 4808 19064 4820
rect 19019 4780 19064 4808
rect 19058 4768 19064 4780
rect 19116 4768 19122 4820
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 8662 4740 8668 4752
rect 2740 4712 8668 4740
rect 2740 4700 2746 4712
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 12710 4700 12716 4752
rect 12768 4749 12774 4752
rect 12768 4743 12832 4749
rect 12768 4709 12786 4743
rect 12820 4709 12832 4743
rect 12768 4703 12832 4709
rect 16660 4743 16718 4749
rect 16660 4709 16672 4743
rect 16706 4740 16718 4743
rect 17126 4740 17132 4752
rect 16706 4712 17132 4740
rect 16706 4709 16718 4712
rect 16660 4703 16718 4709
rect 12768 4700 12774 4703
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1452 4644 1777 4672
rect 1452 4632 1458 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 1765 4635 1823 4641
rect 2032 4675 2090 4681
rect 2032 4641 2044 4675
rect 2078 4672 2090 4675
rect 2866 4672 2872 4684
rect 2078 4644 2872 4672
rect 2078 4641 2090 4644
rect 2032 4635 2090 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5040 4644 5457 4672
rect 5040 4632 5046 4644
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5712 4675 5770 4681
rect 5712 4641 5724 4675
rect 5758 4672 5770 4675
rect 5994 4672 6000 4684
rect 5758 4644 6000 4672
rect 5758 4641 5770 4644
rect 5712 4635 5770 4641
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7616 4644 8033 4672
rect 7616 4632 7622 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10410 4672 10416 4684
rect 10091 4644 10416 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11471 4644 13676 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 10134 4604 10140 4616
rect 8260 4576 8305 4604
rect 10095 4576 10140 4604
rect 8260 4564 8266 4576
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10318 4604 10324 4616
rect 10279 4576 10324 4604
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12400 4576 12541 4604
rect 12400 4564 12406 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 13648 4604 13676 4644
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 13780 4644 15301 4672
rect 13780 4632 13786 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 15896 4644 16405 4672
rect 15896 4632 15902 4644
rect 16393 4641 16405 4644
rect 16439 4672 16451 4675
rect 18138 4672 18144 4684
rect 16439 4644 18144 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 15562 4604 15568 4616
rect 13648 4576 15568 4604
rect 12529 4567 12587 4573
rect 8220 4536 8248 4564
rect 6380 4508 8248 4536
rect 9677 4539 9735 4545
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 6380 4468 6408 4508
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 12158 4536 12164 4548
rect 9723 4508 12164 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 4948 4440 6408 4468
rect 4948 4428 4954 4440
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 6914 4468 6920 4480
rect 6696 4440 6920 4468
rect 6696 4428 6702 4440
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7650 4468 7656 4480
rect 7611 4440 7656 4468
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12434 4468 12440 4480
rect 11655 4440 12440 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 12544 4468 12572 4567
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 19150 4604 19156 4616
rect 19111 4576 19156 4604
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19334 4604 19340 4616
rect 19295 4576 19340 4604
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 14458 4536 14464 4548
rect 13464 4508 14464 4536
rect 13464 4468 13492 4508
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 13906 4468 13912 4480
rect 12544 4440 13492 4468
rect 13867 4440 13912 4468
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 15470 4468 15476 4480
rect 15431 4440 15476 4468
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 17770 4468 17776 4480
rect 17731 4440 17776 4468
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18693 4471 18751 4477
rect 18693 4437 18705 4471
rect 18739 4468 18751 4471
rect 19334 4468 19340 4480
rect 18739 4440 19340 4468
rect 18739 4437 18751 4440
rect 18693 4431 18751 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 4982 4264 4988 4276
rect 3436 4236 4988 4264
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2866 4128 2872 4140
rect 2547 4100 2872 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3436 4137 3464 4236
rect 4632 4208 4660 4236
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 9309 4267 9367 4273
rect 6871 4236 6960 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 4614 4156 4620 4208
rect 4672 4156 4678 4208
rect 4801 4199 4859 4205
rect 4801 4165 4813 4199
rect 4847 4196 4859 4199
rect 4890 4196 4896 4208
rect 4847 4168 4896 4196
rect 4847 4165 4859 4168
rect 4801 4159 4859 4165
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 6932 4196 6960 4236
rect 9309 4233 9321 4267
rect 9355 4264 9367 4267
rect 10134 4264 10140 4276
rect 9355 4236 10140 4264
rect 9355 4233 9367 4236
rect 9309 4227 9367 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 10928 4236 13124 4264
rect 10928 4224 10934 4236
rect 7098 4196 7104 4208
rect 6932 4168 7104 4196
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 11425 4199 11483 4205
rect 11425 4165 11437 4199
rect 11471 4196 11483 4199
rect 12526 4196 12532 4208
rect 11471 4168 12532 4196
rect 11471 4165 11483 4168
rect 11425 4159 11483 4165
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 12768 4168 13032 4196
rect 12768 4156 12774 4168
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6972 4100 7297 4128
rect 6972 4088 6978 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7285 4091 7343 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 9950 4128 9956 4140
rect 8168 4100 9812 4128
rect 9911 4100 9956 4128
rect 8168 4088 8174 4100
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3677 4063 3735 4069
rect 3677 4060 3689 4063
rect 3016 4032 3689 4060
rect 3016 4020 3022 4032
rect 3677 4029 3689 4032
rect 3723 4029 3735 4063
rect 3677 4023 3735 4029
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4120 4032 7328 4060
rect 4120 4020 4126 4032
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3992 5779 3995
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 5767 3964 7205 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7300 3992 7328 4032
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 7300 3964 9689 3992
rect 7193 3955 7251 3961
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 9784 3992 9812 4100
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 13004 4137 13032 4168
rect 12989 4131 13047 4137
rect 10100 4100 11284 4128
rect 10100 4088 10106 4100
rect 11256 4069 11284 4100
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 13096 4128 13124 4236
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 13688 4236 14780 4264
rect 13688 4224 13694 4236
rect 13832 4168 14688 4196
rect 13832 4128 13860 4168
rect 13096 4100 13860 4128
rect 12989 4091 13047 4097
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 13964 4100 14565 4128
rect 13964 4088 13970 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4029 11299 4063
rect 12710 4060 12716 4072
rect 11241 4023 11299 4029
rect 11348 4032 12716 4060
rect 11348 3992 11376 4032
rect 12710 4020 12716 4032
rect 12768 4060 12774 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12768 4032 12909 4060
rect 12768 4020 12774 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14240 4032 14381 4060
rect 14240 4020 14246 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 9784 3964 11376 3992
rect 12452 3964 14473 3992
rect 9677 3955 9735 3961
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2222 3924 2228 3936
rect 2183 3896 2228 3924
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 2406 3924 2412 3936
rect 2363 3896 2412 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 5074 3924 5080 3936
rect 3384 3896 5080 3924
rect 3384 3884 3390 3896
rect 5074 3884 5080 3896
rect 5132 3924 5138 3936
rect 9582 3924 9588 3936
rect 5132 3896 9588 3924
rect 5132 3884 5138 3896
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9640 3896 9781 3924
rect 9640 3884 9646 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 12342 3924 12348 3936
rect 11020 3896 12348 3924
rect 11020 3884 11026 3896
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12452 3933 12480 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14660 3992 14688 4168
rect 14752 4128 14780 4236
rect 17126 4196 17132 4208
rect 16500 4168 17132 4196
rect 16390 4128 16396 4140
rect 14752 4100 16396 4128
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16500 4137 16528 4168
rect 17126 4156 17132 4168
rect 17184 4156 17190 4208
rect 18046 4156 18052 4208
rect 18104 4156 18110 4208
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4097 16543 4131
rect 16485 4091 16543 4097
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 18064 4069 18092 4156
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 18782 4128 18788 4140
rect 18371 4100 18788 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 15252 4032 16313 4060
rect 15252 4020 15258 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 19702 4069 19708 4072
rect 19429 4063 19487 4069
rect 19429 4060 19441 4063
rect 18196 4032 19441 4060
rect 18196 4020 18202 4032
rect 19429 4029 19441 4032
rect 19475 4029 19487 4063
rect 19696 4060 19708 4069
rect 19663 4032 19708 4060
rect 19429 4023 19487 4029
rect 19696 4023 19708 4032
rect 19702 4020 19708 4023
rect 19760 4020 19766 4072
rect 17678 3992 17684 4004
rect 14660 3964 17684 3992
rect 14461 3955 14519 3961
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 19610 3992 19616 4004
rect 18012 3964 19616 3992
rect 18012 3952 18018 3964
rect 19610 3952 19616 3964
rect 19668 3992 19674 4004
rect 21818 3992 21824 4004
rect 19668 3964 21824 3992
rect 19668 3952 19674 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12805 3927 12863 3933
rect 12805 3893 12817 3927
rect 12851 3924 12863 3927
rect 12894 3924 12900 3936
rect 12851 3896 12900 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 15654 3924 15660 3936
rect 14047 3896 15660 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16206 3924 16212 3936
rect 16167 3896 16212 3924
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 18874 3924 18880 3936
rect 17368 3896 18880 3924
rect 17368 3884 17374 3896
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 20806 3924 20812 3936
rect 20767 3896 20812 3924
rect 20806 3884 20812 3896
rect 20864 3884 20870 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 2406 3720 2412 3732
rect 2367 3692 2412 3720
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 7156 3692 7205 3720
rect 7156 3680 7162 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 7193 3683 7251 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10134 3720 10140 3732
rect 9824 3692 10140 3720
rect 9824 3680 9830 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10962 3720 10968 3732
rect 10376 3692 10968 3720
rect 10376 3680 10382 3692
rect 10962 3680 10968 3692
rect 11020 3720 11026 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 11020 3692 11069 3720
rect 11020 3680 11026 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11057 3683 11115 3689
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 15470 3720 15476 3732
rect 14148 3692 15476 3720
rect 14148 3680 14154 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 15896 3692 16957 3720
rect 15896 3680 15902 3692
rect 16945 3689 16957 3692
rect 16991 3689 17003 3723
rect 16945 3683 17003 3689
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 19150 3720 19156 3732
rect 18095 3692 19156 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 198 3612 204 3664
rect 256 3652 262 3664
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 256 3624 2881 3652
rect 256 3612 262 3624
rect 2869 3621 2881 3624
rect 2915 3652 2927 3655
rect 3142 3652 3148 3664
rect 2915 3624 3148 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 11974 3652 11980 3664
rect 4120 3624 5672 3652
rect 4120 3612 4126 3624
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 2682 3448 2688 3460
rect 1084 3420 2688 3448
rect 1084 3408 1090 3420
rect 2682 3408 2688 3420
rect 2740 3448 2746 3460
rect 2792 3448 2820 3547
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4614 3584 4620 3596
rect 4028 3556 4620 3584
rect 4028 3544 4034 3556
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4890 3593 4896 3596
rect 4884 3584 4896 3593
rect 4851 3556 4896 3584
rect 4884 3547 4896 3556
rect 4890 3544 4896 3547
rect 4948 3544 4954 3596
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 5644 3516 5672 3624
rect 5828 3624 11980 3652
rect 5828 3516 5856 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12250 3652 12256 3664
rect 12211 3624 12256 3652
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 13872 3624 19748 3652
rect 13872 3612 13878 3624
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6788 3556 7420 3584
rect 6788 3544 6794 3556
rect 5644 3488 5856 3516
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7392 3525 7420 3556
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 8110 3584 8116 3596
rect 7524 3556 8116 3584
rect 7524 3544 7530 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 9766 3544 9772 3596
rect 9824 3544 9830 3596
rect 9950 3593 9956 3596
rect 9944 3584 9956 3593
rect 9911 3556 9956 3584
rect 9944 3547 9956 3556
rect 9950 3544 9956 3547
rect 10008 3544 10014 3596
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 11940 3556 12357 3584
rect 11940 3544 11946 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 12676 3556 13461 3584
rect 12676 3544 12682 3556
rect 13449 3553 13461 3556
rect 13495 3553 13507 3587
rect 13449 3547 13507 3553
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 13780 3556 13825 3584
rect 13780 3544 13786 3556
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 16850 3584 16856 3596
rect 15344 3556 15389 3584
rect 16811 3556 16856 3584
rect 15344 3544 15350 3556
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 18414 3584 18420 3596
rect 18375 3556 18420 3584
rect 18414 3544 18420 3556
rect 18472 3584 18478 3596
rect 19720 3593 19748 3624
rect 18877 3587 18935 3593
rect 18877 3584 18889 3587
rect 18472 3556 18889 3584
rect 18472 3544 18478 3556
rect 18877 3553 18889 3556
rect 18923 3553 18935 3587
rect 18877 3547 18935 3553
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 6972 3488 7297 3516
rect 6972 3476 6978 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 2740 3420 2820 3448
rect 2740 3408 2746 3420
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 4062 3448 4068 3460
rect 3292 3420 4068 3448
rect 3292 3408 3298 3420
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 5994 3448 6000 3460
rect 5907 3420 6000 3448
rect 5994 3408 6000 3420
rect 6052 3448 6058 3460
rect 7484 3448 7512 3544
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 9784 3516 9812 3544
rect 7616 3488 9812 3516
rect 12529 3519 12587 3525
rect 7616 3476 7622 3488
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12986 3516 12992 3528
rect 12575 3488 12992 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 17129 3519 17187 3525
rect 13872 3488 16344 3516
rect 13872 3476 13878 3488
rect 6052 3420 7512 3448
rect 16316 3448 16344 3488
rect 17129 3485 17141 3519
rect 17175 3516 17187 3519
rect 17770 3516 17776 3528
rect 17175 3488 17776 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3485 18567 3519
rect 18690 3516 18696 3528
rect 18651 3488 18696 3516
rect 18509 3479 18567 3485
rect 17957 3451 18015 3457
rect 17957 3448 17969 3451
rect 16316 3420 17969 3448
rect 6052 3408 6058 3420
rect 17957 3417 17969 3420
rect 18003 3448 18015 3451
rect 18524 3448 18552 3479
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 18003 3420 18552 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 6546 3380 6552 3392
rect 624 3352 6552 3380
rect 624 3340 630 3352
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6822 3380 6828 3392
rect 6783 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 10042 3380 10048 3392
rect 7524 3352 10048 3380
rect 7524 3340 7530 3352
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 10594 3380 10600 3392
rect 10376 3352 10600 3380
rect 10376 3340 10382 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 11885 3383 11943 3389
rect 11885 3380 11897 3383
rect 11848 3352 11897 3380
rect 11848 3340 11854 3352
rect 11885 3349 11897 3352
rect 11931 3349 11943 3383
rect 11885 3343 11943 3349
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 15473 3383 15531 3389
rect 15473 3380 15485 3383
rect 13320 3352 15485 3380
rect 13320 3340 13326 3352
rect 15473 3349 15485 3352
rect 15519 3349 15531 3383
rect 16482 3380 16488 3392
rect 16443 3352 16488 3380
rect 15473 3343 15531 3349
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 19889 3383 19947 3389
rect 19889 3349 19901 3383
rect 19935 3380 19947 3383
rect 21358 3380 21364 3392
rect 19935 3352 21364 3380
rect 19935 3349 19947 3352
rect 19889 3343 19947 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 3108 3148 5549 3176
rect 3108 3136 3114 3148
rect 5537 3145 5549 3148
rect 5583 3145 5595 3179
rect 5537 3139 5595 3145
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 7374 3176 7380 3188
rect 6236 3148 7380 3176
rect 6236 3136 6242 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 9858 3176 9864 3188
rect 7760 3148 9864 3176
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 1452 3012 1501 3040
rect 1452 3000 1458 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 7558 3040 7564 3052
rect 2556 3012 4292 3040
rect 2556 3000 2562 3012
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 4028 2944 4169 2972
rect 4028 2932 4034 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 4264 2972 4292 3012
rect 6472 3012 7564 3040
rect 6472 2972 6500 3012
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 7760 3049 7788 3148
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10502 3176 10508 3188
rect 10192 3148 10508 3176
rect 10192 3136 10198 3148
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 12250 3176 12256 3188
rect 10612 3148 12256 3176
rect 10612 3108 10640 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13170 3176 13176 3188
rect 12492 3148 12537 3176
rect 12820 3148 13176 3176
rect 12492 3136 12498 3148
rect 10060 3080 10640 3108
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8202 3040 8208 3052
rect 7975 3012 8208 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8846 3040 8852 3052
rect 8807 3012 8852 3040
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 4264 2944 6500 2972
rect 4157 2935 4215 2941
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 6604 2944 7665 2972
rect 6604 2932 6610 2944
rect 7653 2941 7665 2944
rect 7699 2972 7711 2975
rect 10060 2972 10088 3080
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 12820 3108 12848 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 16022 3176 16028 3188
rect 14700 3148 16028 3176
rect 14700 3136 14706 3148
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 20622 3136 20628 3188
rect 20680 3176 20686 3188
rect 20990 3176 20996 3188
rect 20680 3148 20996 3176
rect 20680 3136 20686 3148
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 10744 3080 12848 3108
rect 10744 3068 10750 3080
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 20806 3108 20812 3120
rect 14976 3080 20812 3108
rect 14976 3068 14982 3080
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 12802 3000 12808 3052
rect 12860 3040 12866 3052
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12860 3012 12909 3040
rect 12860 3000 12866 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13044 3012 13089 3040
rect 13044 3000 13050 3012
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 14550 3040 14556 3052
rect 13412 3012 14412 3040
rect 14511 3012 14556 3040
rect 13412 3000 13418 3012
rect 7699 2944 10088 2972
rect 11057 2975 11115 2981
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 11057 2941 11069 2975
rect 11103 2972 11115 2975
rect 12618 2972 12624 2984
rect 11103 2944 12624 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 14384 2981 14412 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 15620 3012 15853 3040
rect 15620 3000 15626 3012
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 16908 3012 16957 3040
rect 16908 3000 16914 3012
rect 16945 3009 16957 3012
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18966 3040 18972 3052
rect 18288 3012 18972 3040
rect 18288 3000 18294 3012
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19518 3040 19524 3052
rect 19479 3012 19524 3040
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 14379 2975 14437 2981
rect 14379 2941 14391 2975
rect 14425 2941 14437 2975
rect 15654 2972 15660 2984
rect 15615 2944 15660 2972
rect 14379 2935 14437 2941
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 16540 2944 18061 2972
rect 16540 2932 16546 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 19334 2972 19340 2984
rect 19295 2944 19340 2972
rect 18049 2935 18107 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 20809 2975 20867 2981
rect 20809 2941 20821 2975
rect 20855 2972 20867 2975
rect 22738 2972 22744 2984
rect 20855 2944 22744 2972
rect 20855 2941 20867 2944
rect 20809 2935 20867 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 1756 2907 1814 2913
rect 1756 2873 1768 2907
rect 1802 2904 1814 2907
rect 3050 2904 3056 2916
rect 1802 2876 3056 2904
rect 1802 2873 1814 2876
rect 1756 2867 1814 2873
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 4424 2907 4482 2913
rect 3160 2876 4108 2904
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3160 2836 3188 2876
rect 2832 2808 3188 2836
rect 2832 2796 2838 2808
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3970 2836 3976 2848
rect 3568 2808 3976 2836
rect 3568 2796 3574 2808
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4080 2836 4108 2876
rect 4424 2873 4436 2907
rect 4470 2904 4482 2907
rect 9116 2907 9174 2913
rect 4470 2876 9076 2904
rect 4470 2873 4482 2876
rect 4424 2867 4482 2873
rect 7006 2836 7012 2848
rect 4080 2808 7012 2836
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7282 2836 7288 2848
rect 7243 2808 7288 2836
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 9048 2836 9076 2876
rect 9116 2873 9128 2907
rect 9162 2904 9174 2907
rect 9674 2904 9680 2916
rect 9162 2876 9680 2904
rect 9162 2873 9174 2876
rect 9116 2867 9174 2873
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 11333 2907 11391 2913
rect 9824 2876 10364 2904
rect 9824 2864 9830 2876
rect 10042 2836 10048 2848
rect 9048 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2836 10106 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10100 2808 10241 2836
rect 10100 2796 10106 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 10336 2836 10364 2876
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 13722 2904 13728 2916
rect 11379 2876 13728 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 15194 2904 15200 2916
rect 13823 2876 15200 2904
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 10336 2808 12817 2836
rect 10229 2799 10287 2805
rect 12805 2805 12817 2808
rect 12851 2836 12863 2839
rect 13823 2836 13851 2876
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 17218 2904 17224 2916
rect 16040 2876 17224 2904
rect 12851 2808 13851 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 16040 2836 16068 2876
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 20254 2904 20260 2916
rect 18371 2876 20260 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 14608 2808 16068 2836
rect 14608 2796 14614 2808
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 18138 2836 18144 2848
rect 16172 2808 18144 2836
rect 16172 2796 16178 2808
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2280 2604 2421 2632
rect 2280 2592 2286 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 2409 2595 2467 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7340 2604 7389 2632
rect 7340 2592 7346 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 10410 2632 10416 2644
rect 8711 2604 10416 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 12434 2632 12440 2644
rect 11195 2604 12440 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 17218 2632 17224 2644
rect 14792 2604 17080 2632
rect 17179 2604 17224 2632
rect 14792 2592 14798 2604
rect 1946 2524 1952 2576
rect 2004 2564 2010 2576
rect 2869 2567 2927 2573
rect 2869 2564 2881 2567
rect 2004 2536 2881 2564
rect 2004 2524 2010 2536
rect 2869 2533 2881 2536
rect 2915 2564 2927 2567
rect 3970 2564 3976 2576
rect 2915 2536 3976 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 11241 2567 11299 2573
rect 4571 2536 8432 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 4246 2496 4252 2508
rect 2832 2468 2877 2496
rect 4207 2468 4252 2496
rect 2832 2456 2838 2468
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 6822 2496 6828 2508
rect 5583 2468 6828 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7650 2496 7656 2508
rect 7331 2468 7656 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8202 2428 8208 2440
rect 7607 2400 8208 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 5828 2360 5856 2391
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8404 2428 8432 2536
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11790 2564 11796 2576
rect 11287 2536 11796 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 12158 2524 12164 2576
rect 12216 2564 12222 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12216 2536 13001 2564
rect 12216 2524 12222 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 15286 2564 15292 2576
rect 12989 2527 13047 2533
rect 13096 2536 15292 2564
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 11146 2496 11152 2508
rect 9815 2468 11152 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 13096 2496 13124 2536
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 16025 2567 16083 2573
rect 16025 2533 16037 2567
rect 16071 2564 16083 2567
rect 16758 2564 16764 2576
rect 16071 2536 16764 2564
rect 16071 2533 16083 2536
rect 16025 2527 16083 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 11256 2468 13124 2496
rect 11256 2428 11284 2468
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13780 2468 14197 2496
rect 13780 2456 13786 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15746 2496 15752 2508
rect 15707 2468 15752 2496
rect 14185 2459 14243 2465
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 17052 2505 17080 2604
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 18196 2604 19625 2632
rect 18196 2592 18202 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 19613 2595 19671 2601
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 20162 2496 20168 2508
rect 19475 2468 20168 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 8404 2400 11284 2428
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 10781 2363 10839 2369
rect 5828 2332 7512 2360
rect 7484 2304 7512 2332
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11238 2360 11244 2372
rect 10827 2332 11244 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 7466 2252 7472 2304
rect 7524 2252 7530 2304
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 10962 2292 10968 2304
rect 9732 2264 10968 2292
rect 9732 2252 9738 2264
rect 10962 2252 10968 2264
rect 11020 2292 11026 2304
rect 11348 2292 11376 2391
rect 11514 2320 11520 2372
rect 11572 2360 11578 2372
rect 13096 2360 13124 2391
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13228 2400 13273 2428
rect 13228 2388 13234 2400
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 18340 2428 18368 2459
rect 20162 2456 20168 2468
rect 20220 2456 20226 2508
rect 14424 2400 18368 2428
rect 14424 2388 14430 2400
rect 11572 2332 13124 2360
rect 11572 2320 11578 2332
rect 11020 2264 11376 2292
rect 11020 2252 11026 2264
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 12860 2264 14381 2292
rect 12860 2252 12866 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 15068 2264 18521 2292
rect 15068 2252 15074 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3970 1572 3976 1624
rect 4028 1612 4034 1624
rect 10318 1612 10324 1624
rect 4028 1584 10324 1612
rect 4028 1572 4034 1584
rect 10318 1572 10324 1584
rect 10376 1572 10382 1624
rect 15470 1436 15476 1488
rect 15528 1476 15534 1488
rect 16114 1476 16120 1488
rect 15528 1448 16120 1476
rect 15528 1436 15534 1448
rect 16114 1436 16120 1448
rect 16172 1436 16178 1488
rect 12526 960 12532 1012
rect 12584 1000 12590 1012
rect 13722 1000 13728 1012
rect 12584 972 13728 1000
rect 12584 960 12590 972
rect 13722 960 13728 972
rect 13780 960 13786 1012
rect 19518 552 19524 604
rect 19576 592 19582 604
rect 19886 592 19892 604
rect 19576 564 19892 592
rect 19576 552 19582 564
rect 19886 552 19892 564
rect 19944 552 19950 604
<< via1 >>
rect 4068 20952 4120 21004
rect 12808 20952 12860 21004
rect 3976 20884 4028 20936
rect 12532 20884 12584 20936
rect 3792 20816 3844 20868
rect 13912 20816 13964 20868
rect 3884 20748 3936 20800
rect 13636 20748 13688 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 3976 20544 4028 20596
rect 12808 20587 12860 20596
rect 12808 20553 12817 20587
rect 12817 20553 12851 20587
rect 12851 20553 12860 20587
rect 12808 20544 12860 20553
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 4068 20476 4120 20528
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 5172 20340 5224 20392
rect 7104 20408 7156 20460
rect 7012 20340 7064 20392
rect 9772 20383 9824 20392
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 10876 20383 10928 20392
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 13728 20383 13780 20392
rect 13728 20349 13737 20383
rect 13737 20349 13771 20383
rect 13771 20349 13780 20383
rect 13728 20340 13780 20349
rect 11244 20272 11296 20324
rect 3516 20204 3568 20256
rect 7012 20204 7064 20256
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 10876 20000 10928 20052
rect 12532 20000 12584 20052
rect 2136 19907 2188 19916
rect 2136 19873 2145 19907
rect 2145 19873 2179 19907
rect 2179 19873 2188 19907
rect 2136 19864 2188 19873
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 4160 19864 4212 19916
rect 8208 19932 8260 19984
rect 9772 19932 9824 19984
rect 13728 19932 13780 19984
rect 5356 19907 5408 19916
rect 5356 19873 5365 19907
rect 5365 19873 5399 19907
rect 5399 19873 5408 19907
rect 5356 19864 5408 19873
rect 6644 19907 6696 19916
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 6644 19873 6653 19907
rect 6653 19873 6687 19907
rect 6687 19873 6696 19907
rect 6644 19864 6696 19873
rect 8300 19907 8352 19916
rect 8300 19873 8309 19907
rect 8309 19873 8343 19907
rect 8343 19873 8352 19907
rect 8300 19864 8352 19873
rect 8760 19864 8812 19916
rect 10508 19864 10560 19916
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 8668 19796 8720 19848
rect 10968 19796 11020 19848
rect 8760 19728 8812 19780
rect 10048 19728 10100 19780
rect 11244 19864 11296 19916
rect 17224 19907 17276 19916
rect 12440 19728 12492 19780
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 3884 19660 3936 19712
rect 8576 19660 8628 19712
rect 13636 19728 13688 19780
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 2228 19456 2280 19508
rect 7656 19456 7708 19508
rect 8300 19456 8352 19508
rect 12440 19499 12492 19508
rect 12440 19465 12449 19499
rect 12449 19465 12483 19499
rect 12483 19465 12492 19499
rect 12440 19456 12492 19465
rect 5632 19388 5684 19440
rect 12624 19388 12676 19440
rect 5172 19320 5224 19372
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 11428 19320 11480 19372
rect 14004 19320 14056 19372
rect 6736 19184 6788 19236
rect 2412 19116 2464 19168
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 4896 19116 4948 19168
rect 8484 19252 8536 19304
rect 12992 19184 13044 19236
rect 20904 19184 20956 19236
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 9496 19159 9548 19168
rect 7288 19116 7340 19125
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 9680 19116 9732 19168
rect 9772 19116 9824 19168
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 20720 19159 20772 19168
rect 12900 19116 12952 19125
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 4620 18912 4672 18964
rect 5172 18844 5224 18896
rect 2412 18819 2464 18828
rect 2412 18785 2421 18819
rect 2421 18785 2455 18819
rect 2455 18785 2464 18819
rect 2412 18776 2464 18785
rect 3792 18708 3844 18760
rect 7472 18912 7524 18964
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 12808 18912 12860 18964
rect 7564 18844 7616 18896
rect 11428 18844 11480 18896
rect 8944 18776 8996 18828
rect 10600 18776 10652 18828
rect 12624 18776 12676 18828
rect 7104 18708 7156 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 11060 18708 11112 18760
rect 4068 18572 4120 18624
rect 9772 18572 9824 18624
rect 11980 18572 12032 18624
rect 12716 18572 12768 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 5172 18368 5224 18420
rect 5724 18368 5776 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 20720 18368 20772 18420
rect 12624 18275 12676 18284
rect 3424 18164 3476 18216
rect 3792 18164 3844 18216
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 6644 18164 6696 18216
rect 7104 18164 7156 18216
rect 9772 18164 9824 18216
rect 12716 18164 12768 18216
rect 5448 18096 5500 18148
rect 7472 18096 7524 18148
rect 4068 18028 4120 18080
rect 8300 18096 8352 18148
rect 11060 18096 11112 18148
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 14004 18071 14056 18080
rect 14004 18037 14013 18071
rect 14013 18037 14047 18071
rect 14047 18037 14056 18071
rect 14004 18028 14056 18037
rect 19248 18028 19300 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 4896 17867 4948 17876
rect 4896 17833 4905 17867
rect 4905 17833 4939 17867
rect 4939 17833 4948 17867
rect 4896 17824 4948 17833
rect 7288 17824 7340 17876
rect 4344 17688 4396 17740
rect 2412 17620 2464 17672
rect 6184 17688 6236 17740
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 9496 17824 9548 17876
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 12992 17867 13044 17876
rect 8300 17756 8352 17808
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 8944 17688 8996 17740
rect 9772 17688 9824 17740
rect 10692 17688 10744 17740
rect 11152 17688 11204 17740
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 7564 17663 7616 17672
rect 5448 17620 5500 17629
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 8484 17552 8536 17604
rect 4068 17484 4120 17536
rect 7012 17484 7064 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 4068 17280 4120 17332
rect 5448 17280 5500 17332
rect 5540 17280 5592 17332
rect 9772 17280 9824 17332
rect 10692 17280 10744 17332
rect 12900 17280 12952 17332
rect 3792 17119 3844 17128
rect 3792 17085 3801 17119
rect 3801 17085 3835 17119
rect 3835 17085 3844 17119
rect 3792 17076 3844 17085
rect 9772 17144 9824 17196
rect 10324 17144 10376 17196
rect 12716 17144 12768 17196
rect 5172 17076 5224 17128
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 6920 17076 6972 17128
rect 3700 17008 3752 17060
rect 4988 17008 5040 17060
rect 5356 17008 5408 17060
rect 4160 16940 4212 16992
rect 9772 17008 9824 17060
rect 11704 17008 11756 17060
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 8300 16940 8352 16949
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 10416 16940 10468 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2136 16736 2188 16788
rect 3700 16736 3752 16788
rect 9680 16736 9732 16788
rect 10692 16736 10744 16788
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 4252 16600 4304 16652
rect 5540 16600 5592 16652
rect 6920 16668 6972 16720
rect 8300 16668 8352 16720
rect 8392 16600 8444 16652
rect 4988 16532 5040 16584
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 8208 16532 8260 16584
rect 10416 16600 10468 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 11152 16600 11204 16652
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 3608 16192 3660 16244
rect 4344 16192 4396 16244
rect 4988 16192 5040 16244
rect 9772 16192 9824 16244
rect 11152 16167 11204 16176
rect 11152 16133 11161 16167
rect 11161 16133 11195 16167
rect 11195 16133 11204 16167
rect 11152 16124 11204 16133
rect 2320 15988 2372 16040
rect 3976 15988 4028 16040
rect 6828 15988 6880 16040
rect 6920 15988 6972 16040
rect 9588 15988 9640 16040
rect 9864 15988 9916 16040
rect 11704 15988 11756 16040
rect 5448 15920 5500 15972
rect 8300 15920 8352 15972
rect 10140 15920 10192 15972
rect 4068 15852 4120 15904
rect 8484 15852 8536 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 8852 15852 8904 15904
rect 13176 15852 13228 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 4436 15648 4488 15700
rect 5264 15648 5316 15700
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 5540 15648 5592 15700
rect 4804 15580 4856 15632
rect 7748 15648 7800 15700
rect 9956 15648 10008 15700
rect 10140 15648 10192 15700
rect 2228 15555 2280 15564
rect 2228 15521 2237 15555
rect 2237 15521 2271 15555
rect 2271 15521 2280 15555
rect 2228 15512 2280 15521
rect 3976 15512 4028 15564
rect 2872 15444 2924 15496
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 10692 15580 10744 15632
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 5448 15444 5500 15496
rect 5264 15376 5316 15428
rect 9220 15512 9272 15564
rect 11888 15555 11940 15564
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 11888 15521 11922 15555
rect 11922 15521 11940 15555
rect 11888 15512 11940 15521
rect 8392 15444 8444 15453
rect 5540 15308 5592 15360
rect 8852 15308 8904 15360
rect 9772 15308 9824 15360
rect 10600 15376 10652 15428
rect 11244 15376 11296 15428
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 4068 15104 4120 15156
rect 10048 15104 10100 15156
rect 11244 15104 11296 15156
rect 3976 15036 4028 15088
rect 4344 15036 4396 15088
rect 4896 15036 4948 15088
rect 5172 15079 5224 15088
rect 5172 15045 5181 15079
rect 5181 15045 5215 15079
rect 5215 15045 5224 15079
rect 5172 15036 5224 15045
rect 11888 15104 11940 15156
rect 4712 14968 4764 15020
rect 7012 14968 7064 15020
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2596 14900 2648 14952
rect 3424 14832 3476 14884
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 3792 14832 3844 14841
rect 5540 14900 5592 14952
rect 7380 14900 7432 14952
rect 12440 15036 12492 15088
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 11796 14943 11848 14952
rect 11796 14909 11805 14943
rect 11805 14909 11839 14943
rect 11839 14909 11848 14943
rect 11796 14900 11848 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 12348 14832 12400 14884
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 4436 14764 4488 14816
rect 4896 14764 4948 14816
rect 7288 14764 7340 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3976 14560 4028 14612
rect 4252 14492 4304 14544
rect 4436 14535 4488 14544
rect 4436 14501 4445 14535
rect 4445 14501 4479 14535
rect 4479 14501 4488 14535
rect 4436 14492 4488 14501
rect 1492 14424 1544 14476
rect 2872 14399 2924 14408
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 4712 14560 4764 14612
rect 7748 14560 7800 14612
rect 8208 14560 8260 14612
rect 8484 14560 8536 14612
rect 12348 14560 12400 14612
rect 5816 14492 5868 14544
rect 11244 14492 11296 14544
rect 7564 14424 7616 14476
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 11704 14424 11756 14476
rect 1768 14288 1820 14340
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 2872 14220 2924 14272
rect 7748 14356 7800 14408
rect 6736 14288 6788 14340
rect 7196 14288 7248 14340
rect 5264 14220 5316 14272
rect 5540 14220 5592 14272
rect 8484 14288 8536 14340
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 3884 14016 3936 14068
rect 7748 14016 7800 14068
rect 10416 14016 10468 14068
rect 2504 13948 2556 14000
rect 1768 13880 1820 13932
rect 3332 13880 3384 13932
rect 3976 13880 4028 13932
rect 3056 13812 3108 13864
rect 7380 13948 7432 14000
rect 5540 13880 5592 13932
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 11704 13880 11756 13932
rect 5724 13812 5776 13864
rect 10600 13812 10652 13864
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 3240 13676 3292 13728
rect 4344 13676 4396 13728
rect 7288 13744 7340 13796
rect 5632 13676 5684 13728
rect 8392 13676 8444 13728
rect 8760 13744 8812 13796
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 10600 13676 10652 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2228 13472 2280 13524
rect 3148 13472 3200 13524
rect 4160 13472 4212 13524
rect 5816 13472 5868 13524
rect 7380 13472 7432 13524
rect 8208 13472 8260 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 10324 13515 10376 13524
rect 8484 13472 8536 13481
rect 10324 13481 10333 13515
rect 10333 13481 10367 13515
rect 10367 13481 10376 13515
rect 10324 13472 10376 13481
rect 11704 13472 11756 13524
rect 2872 13447 2924 13456
rect 2872 13413 2881 13447
rect 2881 13413 2915 13447
rect 2915 13413 2924 13447
rect 2872 13404 2924 13413
rect 3424 13404 3476 13456
rect 3792 13336 3844 13388
rect 3976 13268 4028 13320
rect 2964 13200 3016 13252
rect 5632 13404 5684 13456
rect 10416 13404 10468 13456
rect 4344 13336 4396 13388
rect 7012 13336 7064 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 11152 13336 11204 13388
rect 8760 13268 8812 13320
rect 11244 13268 11296 13320
rect 3516 13132 3568 13184
rect 6276 13132 6328 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1584 12928 1636 12980
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 11796 12928 11848 12980
rect 4804 12792 4856 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 2044 12724 2096 12776
rect 4436 12724 4488 12776
rect 7564 12724 7616 12776
rect 3332 12656 3384 12708
rect 6552 12656 6604 12708
rect 7840 12724 7892 12776
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 8208 12656 8260 12708
rect 9588 12656 9640 12708
rect 9680 12656 9732 12708
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 9128 12631 9180 12640
rect 5632 12588 5684 12597
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 3240 12384 3292 12436
rect 7012 12384 7064 12436
rect 7380 12384 7432 12436
rect 4436 12316 4488 12368
rect 11244 12316 11296 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 4160 12248 4212 12300
rect 4252 12248 4304 12300
rect 6920 12248 6972 12300
rect 9496 12248 9548 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 8300 12223 8352 12232
rect 2596 12112 2648 12164
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 11704 12248 11756 12300
rect 5540 12112 5592 12164
rect 9680 12112 9732 12164
rect 3424 12044 3476 12096
rect 11152 12044 11204 12096
rect 20628 12044 20680 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 6276 11840 6328 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 10968 11840 11020 11892
rect 12072 11840 12124 11892
rect 12900 11840 12952 11892
rect 8208 11704 8260 11756
rect 9404 11704 9456 11756
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 2044 11636 2096 11688
rect 4344 11636 4396 11688
rect 4804 11679 4856 11688
rect 4804 11645 4838 11679
rect 4838 11645 4856 11679
rect 4804 11636 4856 11645
rect 5540 11636 5592 11688
rect 5816 11636 5868 11688
rect 7104 11636 7156 11688
rect 8576 11679 8628 11688
rect 8576 11645 8610 11679
rect 8610 11645 8628 11679
rect 8576 11636 8628 11645
rect 9128 11636 9180 11688
rect 11060 11679 11112 11688
rect 2596 11568 2648 11620
rect 2780 11568 2832 11620
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11152 11636 11204 11688
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6552 11500 6604 11552
rect 8392 11500 8444 11552
rect 8760 11500 8812 11552
rect 10048 11500 10100 11552
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 10600 11500 10652 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 13268 11543 13320 11552
rect 11152 11500 11204 11509
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 20444 11500 20496 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2320 11296 2372 11348
rect 6828 11296 6880 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 8300 11296 8352 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 9496 11296 9548 11348
rect 5908 11228 5960 11280
rect 6000 11228 6052 11280
rect 3424 11160 3476 11212
rect 4436 11160 4488 11212
rect 3516 11092 3568 11144
rect 4988 11092 5040 11144
rect 5172 11024 5224 11076
rect 7380 11024 7432 11076
rect 7656 11024 7708 11076
rect 9220 11160 9272 11212
rect 10876 11160 10928 11212
rect 11704 11160 11756 11212
rect 12348 11160 12400 11212
rect 12808 11203 12860 11212
rect 12808 11169 12842 11203
rect 12842 11169 12860 11203
rect 12808 11160 12860 11169
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 15844 11135 15896 11144
rect 8576 11092 8628 11101
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 11704 11067 11756 11076
rect 11704 11033 11713 11067
rect 11713 11033 11747 11067
rect 11747 11033 11756 11067
rect 11704 11024 11756 11033
rect 3700 10956 3752 11008
rect 13912 10999 13964 11008
rect 13912 10965 13921 10999
rect 13921 10965 13955 10999
rect 13955 10965 13964 10999
rect 13912 10956 13964 10965
rect 19984 11024 20036 11076
rect 17408 10956 17460 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1676 10752 1728 10804
rect 3976 10752 4028 10804
rect 4804 10752 4856 10804
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 3516 10616 3568 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 3884 10591 3936 10600
rect 3884 10557 3918 10591
rect 3918 10557 3936 10591
rect 3884 10548 3936 10557
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9864 10548 9916 10600
rect 10232 10752 10284 10804
rect 12256 10752 12308 10804
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 13820 10684 13872 10693
rect 16028 10684 16080 10736
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11704 10548 11756 10600
rect 12348 10548 12400 10600
rect 14740 10616 14792 10668
rect 9680 10480 9732 10532
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 10508 10412 10560 10421
rect 11060 10412 11112 10464
rect 11980 10412 12032 10464
rect 13544 10480 13596 10532
rect 13728 10412 13780 10464
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 19432 10412 19484 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2596 10208 2648 10260
rect 4068 10208 4120 10260
rect 6828 10208 6880 10260
rect 8576 10208 8628 10260
rect 11060 10208 11112 10260
rect 12348 10208 12400 10260
rect 9956 10140 10008 10192
rect 10784 10140 10836 10192
rect 1676 10115 1728 10124
rect 1676 10081 1710 10115
rect 1710 10081 1728 10115
rect 1676 10072 1728 10081
rect 4252 10072 4304 10124
rect 6276 10072 6328 10124
rect 9680 10072 9732 10124
rect 12440 10072 12492 10124
rect 16120 10072 16172 10124
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 5080 10004 5132 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 8576 10004 8628 10056
rect 9404 10004 9456 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 3792 9936 3844 9988
rect 10416 9936 10468 9988
rect 12808 9936 12860 9988
rect 15200 10004 15252 10056
rect 18052 10004 18104 10056
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 9404 9868 9456 9920
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 1676 9664 1728 9716
rect 5724 9664 5776 9716
rect 4160 9596 4212 9648
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 1400 9460 1452 9512
rect 3516 9460 3568 9512
rect 5448 9460 5500 9512
rect 16120 9664 16172 9716
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 11888 9596 11940 9648
rect 12072 9596 12124 9648
rect 12164 9596 12216 9648
rect 19432 9596 19484 9648
rect 19892 9596 19944 9648
rect 6368 9460 6420 9512
rect 2504 9392 2556 9444
rect 2596 9392 2648 9444
rect 2872 9392 2924 9444
rect 4896 9392 4948 9444
rect 7380 9460 7432 9512
rect 10784 9528 10836 9580
rect 12348 9528 12400 9580
rect 12900 9528 12952 9580
rect 13912 9528 13964 9580
rect 8576 9460 8628 9512
rect 10968 9460 11020 9512
rect 14924 9460 14976 9512
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 6460 9367 6512 9376
rect 5172 9324 5224 9333
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 7380 9324 7432 9376
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 14740 9324 14792 9376
rect 16304 9392 16356 9444
rect 19616 9392 19668 9444
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1492 9120 1544 9172
rect 4896 9120 4948 9172
rect 5356 9052 5408 9104
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 6000 9052 6052 9104
rect 4344 8984 4396 9036
rect 5540 8984 5592 9036
rect 11060 9120 11112 9172
rect 11704 9120 11756 9172
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 14648 9052 14700 9104
rect 16212 9120 16264 9172
rect 16304 9120 16356 9172
rect 11060 9027 11112 9036
rect 11060 8993 11094 9027
rect 11094 8993 11112 9027
rect 11060 8984 11112 8993
rect 12256 8984 12308 9036
rect 17500 9052 17552 9104
rect 16028 9027 16080 9036
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 18880 8984 18932 9036
rect 4903 8959 4955 8968
rect 4903 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4955 8959
rect 4903 8916 4955 8925
rect 3884 8780 3936 8832
rect 4068 8780 4120 8832
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 16488 8916 16540 8968
rect 19340 8916 19392 8968
rect 7380 8780 7432 8832
rect 8484 8780 8536 8832
rect 9404 8780 9456 8832
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 15200 8780 15252 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1952 8576 2004 8628
rect 3056 8576 3108 8628
rect 5172 8576 5224 8628
rect 5356 8576 5408 8628
rect 9312 8576 9364 8628
rect 9956 8619 10008 8628
rect 3608 8508 3660 8560
rect 3792 8508 3844 8560
rect 6552 8508 6604 8560
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 10140 8576 10192 8628
rect 10416 8576 10468 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 4068 8483 4120 8492
rect 2504 8440 2556 8449
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 6000 8440 6052 8492
rect 9404 8440 9456 8492
rect 2964 8372 3016 8424
rect 3884 8372 3936 8424
rect 7380 8372 7432 8424
rect 8852 8372 8904 8424
rect 8944 8372 8996 8424
rect 10784 8440 10836 8492
rect 13084 8440 13136 8492
rect 14464 8576 14516 8628
rect 17868 8576 17920 8628
rect 18604 8508 18656 8560
rect 20168 8440 20220 8492
rect 11796 8372 11848 8424
rect 15292 8372 15344 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 19524 8372 19576 8424
rect 2780 8304 2832 8356
rect 3056 8304 3108 8356
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4804 8304 4856 8356
rect 6828 8304 6880 8356
rect 9496 8304 9548 8356
rect 13452 8347 13504 8356
rect 13452 8313 13486 8347
rect 13486 8313 13504 8347
rect 13452 8304 13504 8313
rect 19064 8304 19116 8356
rect 4068 8236 4120 8288
rect 9036 8236 9088 8288
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 3424 8032 3476 8084
rect 4896 8032 4948 8084
rect 6000 8032 6052 8084
rect 6736 8032 6788 8084
rect 11244 8032 11296 8084
rect 18880 8075 18932 8084
rect 2228 7896 2280 7948
rect 6460 7964 6512 8016
rect 5540 7939 5592 7948
rect 5540 7905 5574 7939
rect 5574 7905 5592 7939
rect 5540 7896 5592 7905
rect 6736 7896 6788 7948
rect 9588 7964 9640 8016
rect 12164 7964 12216 8016
rect 14556 7964 14608 8016
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 19800 7964 19852 8016
rect 7748 7896 7800 7948
rect 10232 7896 10284 7948
rect 11704 7896 11756 7948
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 4252 7828 4304 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 14188 7871 14240 7880
rect 8300 7760 8352 7812
rect 9128 7760 9180 7812
rect 7380 7692 7432 7744
rect 8392 7692 8444 7744
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 15200 7828 15252 7880
rect 16488 7896 16540 7948
rect 17776 7939 17828 7948
rect 17776 7905 17810 7939
rect 17810 7905 17828 7939
rect 17776 7896 17828 7905
rect 18788 7896 18840 7948
rect 10048 7692 10100 7744
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 11888 7692 11940 7744
rect 13452 7692 13504 7744
rect 16028 7692 16080 7744
rect 18972 7692 19024 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 7748 7488 7800 7540
rect 6828 7420 6880 7472
rect 10416 7420 10468 7472
rect 20904 7488 20956 7540
rect 22284 7488 22336 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 7104 7352 7156 7404
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 12164 7352 12216 7404
rect 18880 7352 18932 7404
rect 3700 7284 3752 7336
rect 6920 7284 6972 7336
rect 7564 7284 7616 7336
rect 8208 7284 8260 7336
rect 9036 7284 9088 7336
rect 12716 7284 12768 7336
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 13728 7284 13780 7336
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 14464 7284 14516 7336
rect 16028 7284 16080 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 1676 7259 1728 7268
rect 1676 7225 1710 7259
rect 1710 7225 1728 7259
rect 1676 7216 1728 7225
rect 4068 7216 4120 7268
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 4252 7148 4304 7200
rect 7012 7148 7064 7200
rect 8668 7216 8720 7268
rect 13912 7216 13964 7268
rect 14372 7216 14424 7268
rect 10232 7148 10284 7200
rect 10600 7148 10652 7200
rect 11980 7148 12032 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 12624 7148 12676 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 19156 7148 19208 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2228 6987 2280 6996
rect 2228 6953 2237 6987
rect 2237 6953 2271 6987
rect 2271 6953 2280 6987
rect 2228 6944 2280 6953
rect 4160 6944 4212 6996
rect 13268 6987 13320 6996
rect 3332 6876 3384 6928
rect 3976 6876 4028 6928
rect 3700 6808 3752 6860
rect 4252 6876 4304 6928
rect 8852 6876 8904 6928
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 7472 6808 7524 6860
rect 8576 6808 8628 6860
rect 13268 6953 13277 6987
rect 13277 6953 13311 6987
rect 13311 6953 13320 6987
rect 13268 6944 13320 6953
rect 15844 6944 15896 6996
rect 18512 6944 18564 6996
rect 19800 6944 19852 6996
rect 9680 6876 9732 6928
rect 12440 6876 12492 6928
rect 19340 6876 19392 6928
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 17408 6808 17460 6860
rect 19616 6808 19668 6860
rect 2596 6740 2648 6792
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 9864 6740 9916 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 1676 6672 1728 6724
rect 3884 6672 3936 6724
rect 4068 6604 4120 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 8668 6604 8720 6656
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 12624 6740 12676 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 13820 6740 13872 6792
rect 16028 6740 16080 6792
rect 17776 6740 17828 6792
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 14004 6672 14056 6724
rect 14464 6715 14516 6724
rect 14464 6681 14473 6715
rect 14473 6681 14507 6715
rect 14507 6681 14516 6715
rect 14464 6672 14516 6681
rect 15292 6715 15344 6724
rect 15292 6681 15301 6715
rect 15301 6681 15335 6715
rect 15335 6681 15344 6715
rect 15292 6672 15344 6681
rect 18420 6672 18472 6724
rect 12532 6604 12584 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2504 6400 2556 6452
rect 5080 6400 5132 6452
rect 3424 6332 3476 6384
rect 8576 6400 8628 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 19800 6400 19852 6452
rect 2780 6264 2832 6316
rect 2964 6264 3016 6316
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 5356 6264 5408 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 9496 6332 9548 6384
rect 12256 6332 12308 6384
rect 5540 6264 5592 6316
rect 9680 6264 9732 6316
rect 10048 6264 10100 6316
rect 13360 6264 13412 6316
rect 14556 6264 14608 6316
rect 16488 6264 16540 6316
rect 6000 6196 6052 6248
rect 7472 6196 7524 6248
rect 10416 6239 10468 6248
rect 10416 6205 10439 6239
rect 10439 6205 10468 6239
rect 10416 6196 10468 6205
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 13912 6196 13964 6248
rect 18144 6196 18196 6248
rect 3516 6128 3568 6180
rect 6920 6128 6972 6180
rect 7104 6171 7156 6180
rect 7104 6137 7138 6171
rect 7138 6137 7156 6171
rect 7104 6128 7156 6137
rect 14740 6128 14792 6180
rect 19340 6171 19392 6180
rect 19340 6137 19374 6171
rect 19374 6137 19392 6171
rect 19340 6128 19392 6137
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 3976 6060 4028 6112
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 11336 6060 11388 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 11704 6060 11756 6112
rect 12348 6060 12400 6112
rect 15752 6060 15804 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2136 5856 2188 5908
rect 5540 5856 5592 5908
rect 2320 5788 2372 5840
rect 3792 5788 3844 5840
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 6000 5788 6052 5840
rect 8392 5856 8444 5908
rect 9404 5856 9456 5908
rect 11060 5856 11112 5908
rect 11336 5856 11388 5908
rect 8852 5788 8904 5840
rect 11244 5788 11296 5840
rect 11520 5788 11572 5840
rect 16120 5856 16172 5908
rect 6828 5720 6880 5772
rect 6920 5720 6972 5772
rect 9680 5720 9732 5772
rect 10048 5720 10100 5772
rect 12348 5720 12400 5772
rect 13084 5720 13136 5772
rect 1860 5652 1912 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3792 5652 3844 5704
rect 5356 5652 5408 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 8852 5652 8904 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 14924 5720 14976 5772
rect 18696 5763 18748 5772
rect 18696 5729 18730 5763
rect 18730 5729 18748 5763
rect 18696 5720 18748 5729
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 18144 5652 18196 5704
rect 4068 5584 4120 5636
rect 5540 5584 5592 5636
rect 4252 5516 4304 5568
rect 7104 5516 7156 5568
rect 8944 5516 8996 5568
rect 12532 5516 12584 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 16488 5516 16540 5568
rect 19340 5516 19392 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 2688 5312 2740 5364
rect 6920 5312 6972 5364
rect 8484 5312 8536 5364
rect 14648 5312 14700 5364
rect 14924 5355 14976 5364
rect 14924 5321 14933 5355
rect 14933 5321 14967 5355
rect 14967 5321 14976 5355
rect 14924 5312 14976 5321
rect 6644 5244 6696 5296
rect 13360 5244 13412 5296
rect 2872 5176 2924 5228
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4896 5176 4948 5228
rect 5540 5176 5592 5228
rect 8576 5176 8628 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 11244 5176 11296 5228
rect 3884 5108 3936 5160
rect 4068 5040 4120 5092
rect 8392 5040 8444 5092
rect 8668 5040 8720 5092
rect 8852 5108 8904 5160
rect 12900 5176 12952 5228
rect 11060 5040 11112 5092
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 3424 4972 3476 5024
rect 3884 4972 3936 5024
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 5080 4972 5132 4981
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 15292 5108 15344 5160
rect 15844 5108 15896 5160
rect 16488 5108 16540 5160
rect 18144 5108 18196 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 13912 5040 13964 5092
rect 14464 5040 14516 5092
rect 17776 5040 17828 5092
rect 18880 5040 18932 5092
rect 14556 4972 14608 5024
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 18696 4972 18748 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2964 4768 3016 4820
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 6828 4811 6880 4820
rect 6828 4777 6837 4811
rect 6837 4777 6871 4811
rect 6871 4777 6880 4811
rect 6828 4768 6880 4777
rect 8208 4768 8260 4820
rect 8852 4768 8904 4820
rect 12440 4768 12492 4820
rect 13636 4768 13688 4820
rect 19064 4811 19116 4820
rect 19064 4777 19073 4811
rect 19073 4777 19107 4811
rect 19107 4777 19116 4811
rect 19064 4768 19116 4777
rect 2688 4700 2740 4752
rect 8668 4700 8720 4752
rect 12716 4700 12768 4752
rect 17132 4700 17184 4752
rect 1400 4632 1452 4684
rect 2872 4632 2924 4684
rect 4988 4632 5040 4684
rect 6000 4632 6052 4684
rect 7564 4632 7616 4684
rect 10416 4632 10468 4684
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 10140 4607 10192 4616
rect 8208 4564 8260 4573
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 12348 4564 12400 4616
rect 13728 4632 13780 4684
rect 15844 4632 15896 4684
rect 18144 4632 18196 4684
rect 4896 4428 4948 4480
rect 12164 4496 12216 4548
rect 6644 4428 6696 4480
rect 6920 4428 6972 4480
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 12440 4428 12492 4480
rect 15568 4564 15620 4616
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 14464 4496 14516 4548
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 13912 4428 13964 4437
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 17776 4471 17828 4480
rect 17776 4437 17785 4471
rect 17785 4437 17819 4471
rect 17819 4437 17828 4471
rect 17776 4428 17828 4437
rect 19340 4428 19392 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2872 4088 2924 4140
rect 4988 4224 5040 4276
rect 4620 4156 4672 4208
rect 4896 4156 4948 4208
rect 10140 4224 10192 4276
rect 10876 4224 10928 4276
rect 7104 4156 7156 4208
rect 12532 4156 12584 4208
rect 12716 4156 12768 4208
rect 6920 4088 6972 4140
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 8116 4088 8168 4140
rect 9956 4131 10008 4140
rect 2964 4020 3016 4072
rect 4068 4020 4120 4072
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10048 4088 10100 4140
rect 13636 4224 13688 4276
rect 13912 4088 13964 4140
rect 12716 4020 12768 4072
rect 14188 4020 14240 4072
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2412 3884 2464 3936
rect 3332 3884 3384 3936
rect 5080 3884 5132 3936
rect 9588 3884 9640 3936
rect 10968 3884 11020 3936
rect 12348 3884 12400 3936
rect 16396 4088 16448 4140
rect 17132 4156 17184 4208
rect 18052 4156 18104 4208
rect 15200 4020 15252 4072
rect 18788 4088 18840 4140
rect 18144 4020 18196 4072
rect 19708 4063 19760 4072
rect 19708 4029 19742 4063
rect 19742 4029 19760 4063
rect 19708 4020 19760 4029
rect 17684 3952 17736 4004
rect 17960 3952 18012 4004
rect 19616 3952 19668 4004
rect 21824 3952 21876 4004
rect 12900 3884 12952 3936
rect 15660 3884 15712 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16212 3927 16264 3936
rect 16212 3893 16221 3927
rect 16221 3893 16255 3927
rect 16255 3893 16264 3927
rect 16212 3884 16264 3893
rect 17316 3884 17368 3936
rect 18880 3884 18932 3936
rect 20812 3927 20864 3936
rect 20812 3893 20821 3927
rect 20821 3893 20855 3927
rect 20855 3893 20864 3927
rect 20812 3884 20864 3893
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 7104 3680 7156 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 9772 3680 9824 3732
rect 10140 3680 10192 3732
rect 10324 3680 10376 3732
rect 10968 3680 11020 3732
rect 14096 3680 14148 3732
rect 15476 3680 15528 3732
rect 15844 3680 15896 3732
rect 19156 3680 19208 3732
rect 204 3612 256 3664
rect 3148 3612 3200 3664
rect 4068 3612 4120 3664
rect 1032 3408 1084 3460
rect 2688 3408 2740 3460
rect 3976 3544 4028 3596
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 4896 3587 4948 3596
rect 4896 3553 4930 3587
rect 4930 3553 4948 3587
rect 4896 3544 4948 3553
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 11980 3612 12032 3664
rect 12256 3655 12308 3664
rect 12256 3621 12265 3655
rect 12265 3621 12299 3655
rect 12299 3621 12308 3655
rect 12256 3612 12308 3621
rect 13820 3612 13872 3664
rect 6736 3544 6788 3596
rect 6920 3476 6972 3528
rect 7472 3544 7524 3596
rect 8116 3544 8168 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 9772 3544 9824 3596
rect 9956 3587 10008 3596
rect 9956 3553 9990 3587
rect 9990 3553 10008 3587
rect 9956 3544 10008 3553
rect 11888 3544 11940 3596
rect 12624 3544 12676 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 16856 3587 16908 3596
rect 15292 3544 15344 3553
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 3240 3408 3292 3460
rect 4068 3408 4120 3460
rect 6000 3451 6052 3460
rect 6000 3417 6009 3451
rect 6009 3417 6043 3451
rect 6043 3417 6052 3451
rect 7564 3476 7616 3528
rect 12992 3476 13044 3528
rect 13820 3476 13872 3528
rect 17776 3476 17828 3528
rect 18696 3519 18748 3528
rect 6000 3408 6052 3417
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 572 3340 624 3392
rect 6552 3340 6604 3392
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 7472 3340 7524 3392
rect 10048 3340 10100 3392
rect 10324 3340 10376 3392
rect 10600 3340 10652 3392
rect 11796 3340 11848 3392
rect 13268 3340 13320 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 21364 3340 21416 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 3056 3136 3108 3188
rect 6184 3136 6236 3188
rect 7380 3136 7432 3188
rect 1400 3000 1452 3052
rect 2504 3000 2556 3052
rect 3976 2932 4028 2984
rect 7564 3000 7616 3052
rect 9864 3136 9916 3188
rect 10140 3136 10192 3188
rect 10508 3136 10560 3188
rect 12256 3136 12308 3188
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 8208 3000 8260 3052
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 6552 2932 6604 2984
rect 10692 3068 10744 3120
rect 13176 3136 13228 3188
rect 14648 3136 14700 3188
rect 16028 3136 16080 3188
rect 20628 3136 20680 3188
rect 20996 3136 21048 3188
rect 14924 3068 14976 3120
rect 20812 3068 20864 3120
rect 12808 3000 12860 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13360 3000 13412 3052
rect 14556 3043 14608 3052
rect 12624 2932 12676 2984
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 15568 3000 15620 3052
rect 16856 3000 16908 3052
rect 18236 3000 18288 3052
rect 18972 3000 19024 3052
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 16488 2932 16540 2984
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 22744 2932 22796 2984
rect 3056 2864 3108 2916
rect 2780 2796 2832 2848
rect 3516 2796 3568 2848
rect 3976 2796 4028 2848
rect 7012 2796 7064 2848
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 9680 2864 9732 2916
rect 9772 2864 9824 2916
rect 10048 2796 10100 2848
rect 13728 2864 13780 2916
rect 15200 2864 15252 2916
rect 14556 2796 14608 2848
rect 17224 2864 17276 2916
rect 20260 2864 20312 2916
rect 16120 2796 16172 2848
rect 18144 2796 18196 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2228 2592 2280 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7288 2592 7340 2644
rect 10416 2592 10468 2644
rect 12440 2592 12492 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 14740 2592 14792 2644
rect 17224 2635 17276 2644
rect 1952 2524 2004 2576
rect 3976 2524 4028 2576
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 4252 2499 4304 2508
rect 2780 2456 2832 2465
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 6828 2456 6880 2508
rect 7656 2456 7708 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 8208 2388 8260 2440
rect 11796 2524 11848 2576
rect 12164 2524 12216 2576
rect 11152 2456 11204 2508
rect 15292 2524 15344 2576
rect 16764 2524 16816 2576
rect 13728 2456 13780 2508
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 17224 2601 17233 2635
rect 17233 2601 17267 2635
rect 17267 2601 17276 2635
rect 17224 2592 17276 2601
rect 18144 2592 18196 2644
rect 11244 2320 11296 2372
rect 7472 2252 7524 2304
rect 9680 2252 9732 2304
rect 10968 2252 11020 2304
rect 11520 2320 11572 2372
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 14372 2388 14424 2440
rect 20168 2456 20220 2508
rect 12808 2252 12860 2304
rect 15016 2252 15068 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3976 1572 4028 1624
rect 10324 1572 10376 1624
rect 15476 1436 15528 1488
rect 16120 1436 16172 1488
rect 12532 960 12584 1012
rect 13728 960 13780 1012
rect 19524 552 19576 604
rect 19892 552 19944 604
<< metal2 >>
rect 4802 22672 4858 22681
rect 4802 22607 4858 22616
rect 3790 22264 3846 22273
rect 3790 22199 3846 22208
rect 3804 20874 3832 22199
rect 3882 21720 3938 21729
rect 3882 21655 3938 21664
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3896 20806 3924 21655
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 21010 4108 21247
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3884 20800 3936 20806
rect 3988 20777 4016 20878
rect 3884 20742 3936 20748
rect 3974 20768 4030 20777
rect 3974 20703 4030 20712
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 16794 2176 19858
rect 2240 19514 2268 20334
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 2410 19952 2466 19961
rect 2410 19887 2412 19896
rect 2464 19887 2466 19896
rect 2412 19858 2464 19864
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 3528 19417 3556 20198
rect 3988 19825 4016 20538
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4080 20369 4108 20470
rect 4066 20360 4122 20369
rect 4066 20295 4122 20304
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 18834 2452 19110
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3804 18222 3832 18702
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 7410 1440 9454
rect 1504 9178 1532 14418
rect 1582 14240 1638 14249
rect 1582 14175 1638 14184
rect 1596 12986 1624 14175
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1688 10810 1716 14894
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1780 13938 1808 14282
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 10690 1808 13874
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1688 10662 1808 10690
rect 1688 10130 1716 10662
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9722 1716 10066
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1964 8634 1992 13670
rect 2240 13530 2268 15506
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 11694 2084 12718
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2332 11354 2360 15982
rect 2424 14793 2452 17614
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 15745 2912 16526
rect 2870 15736 2926 15745
rect 2870 15671 2926 15680
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2410 14784 2466 14793
rect 2410 14719 2466 14728
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2424 10606 2452 14214
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 2516 10606 2544 13942
rect 2608 12170 2636 14894
rect 2884 14414 2912 15438
rect 3436 15162 3464 18158
rect 3804 17134 3832 18158
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3712 16794 3740 17002
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 2872 14408 2924 14414
rect 2792 14368 2872 14396
rect 2792 13274 2820 14368
rect 2872 14350 2924 14356
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13462 2912 14214
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2792 13246 2912 13274
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2792 11626 2820 12242
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2608 10674 2636 11562
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2608 10266 2636 10610
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2516 8498 2544 9386
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 4690 1440 7346
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 6730 1716 7210
rect 2240 7002 2268 7890
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 2516 6458 2544 7822
rect 2608 6798 2636 9386
rect 2792 8362 2820 11562
rect 2884 9738 2912 13246
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2875 9710 2912 9738
rect 2875 9450 2903 9710
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2976 8430 3004 13194
rect 3068 8634 3096 13806
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3160 13530 3188 13670
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3252 12442 3280 13670
rect 3344 12714 3372 13874
rect 3436 13462 3464 14826
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3514 13288 3570 13297
rect 3514 13223 3570 13232
rect 3528 13190 3556 13223
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3422 12880 3478 12889
rect 3422 12815 3478 12824
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 11898 3372 12650
rect 3436 12102 3464 12815
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3238 9072 3294 9081
rect 3238 9007 3294 9016
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6798 2820 7142
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5914 2176 6054
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 204 3664 256 3670
rect 204 3606 256 3612
rect 216 480 244 3606
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 584 480 612 3334
rect 1044 480 1072 3402
rect 1412 3058 1440 4626
rect 1490 4584 1546 4593
rect 1490 4519 1546 4528
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1504 480 1532 4519
rect 1872 3942 1900 5646
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4865 2268 4966
rect 2226 4856 2282 4865
rect 2226 4791 2282 4800
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 2650 2268 3878
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 1964 480 1992 2518
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2332 241 2360 5782
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3738 2452 3878
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2516 1578 2544 2994
rect 2608 2961 2636 6734
rect 2792 6322 2820 6734
rect 2976 6322 3004 8366
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5370 2728 5714
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2700 3466 2728 4694
rect 2884 4690 2912 5170
rect 2976 4826 3004 5646
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 4146 2912 4626
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2884 3194 2912 4082
rect 2976 4078 3004 4762
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3068 3924 3096 8298
rect 3146 4720 3202 4729
rect 3146 4655 3202 4664
rect 2976 3896 3096 3924
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2594 2952 2650 2961
rect 2594 2887 2650 2896
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2514 2820 2790
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2424 1550 2544 1578
rect 2424 480 2452 1550
rect 2792 626 2820 2450
rect 2976 649 3004 3896
rect 3160 3670 3188 4655
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 3194 3096 3470
rect 3252 3466 3280 9007
rect 3436 8090 3464 11154
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 10674 3556 11086
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3528 9518 3556 10610
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3620 8566 3648 16186
rect 3804 16028 3832 17070
rect 3896 16561 3924 19654
rect 4172 18986 4200 19858
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 3988 18958 4200 18986
rect 4632 18970 4660 19110
rect 4620 18964 4672 18970
rect 3988 18057 4016 18958
rect 4620 18906 4672 18912
rect 4066 18864 4122 18873
rect 4066 18799 4122 18808
rect 4080 18630 4108 18799
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4066 18456 4122 18465
rect 4421 18448 4717 18468
rect 4066 18391 4122 18400
rect 4080 18086 4108 18391
rect 4068 18080 4120 18086
rect 3974 18048 4030 18057
rect 4068 18022 4120 18028
rect 3974 17983 4030 17992
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4068 17536 4120 17542
rect 4066 17504 4068 17513
rect 4120 17504 4122 17513
rect 4066 17439 4122 17448
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 17105 4108 17274
rect 4066 17096 4122 17105
rect 4066 17031 4122 17040
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3882 16552 3938 16561
rect 3882 16487 3938 16496
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 3976 16040 4028 16046
rect 3804 16000 3976 16028
rect 3976 15982 4028 15988
rect 3988 15570 4016 15982
rect 4080 15910 4108 16079
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4066 15600 4122 15609
rect 3976 15564 4028 15570
rect 4172 15586 4200 16934
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4122 15558 4200 15586
rect 4066 15535 4122 15544
rect 3976 15506 4028 15512
rect 3988 15094 4016 15506
rect 4066 15192 4122 15201
rect 4066 15127 4068 15136
rect 4120 15127 4122 15136
rect 4068 15098 4120 15104
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3804 13394 3832 14826
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 14074 3924 14758
rect 4066 14648 4122 14657
rect 3976 14612 4028 14618
rect 4122 14606 4200 14634
rect 4066 14583 4122 14592
rect 3976 14554 4028 14560
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3988 13938 4016 14554
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4066 13832 4122 13841
rect 4066 13767 4122 13776
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12986 4016 13262
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3988 12730 4016 12922
rect 3896 12702 4016 12730
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3790 10976 3846 10985
rect 3712 10033 3740 10950
rect 3790 10911 3846 10920
rect 3698 10024 3754 10033
rect 3804 9994 3832 10911
rect 3896 10606 3924 12702
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3988 10810 4016 11319
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 4080 10266 4108 13767
rect 4172 13530 4200 14606
rect 4264 14550 4292 16594
rect 4356 16250 4384 17682
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4356 16130 4384 16186
rect 4356 16102 4476 16130
rect 4448 15706 4476 16102
rect 4816 15858 4844 22607
rect 5722 22520 5778 23000
rect 17222 22520 17278 23000
rect 5172 20392 5224 20398
rect 5224 20352 5580 20380
rect 5172 20334 5224 20340
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 17882 4936 19110
rect 5184 18902 5212 19314
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5184 18426 5212 18838
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16590 5028 17002
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 16250 5028 16526
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4816 15830 4936 15858
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4356 13734 4384 15030
rect 4712 15020 4764 15026
rect 4816 15008 4844 15574
rect 4908 15094 4936 15830
rect 5184 15094 5212 17070
rect 5368 17066 5396 19858
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5460 17678 5488 18090
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5460 17338 5488 17614
rect 5552 17338 5580 20352
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5644 19446 5672 19790
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 5736 18426 5764 22520
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7012 20392 7064 20398
rect 6932 20352 7012 20380
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 6656 18222 6684 19858
rect 6932 19258 6960 20352
rect 7012 20334 7064 20340
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6748 19242 6960 19258
rect 6736 19236 6960 19242
rect 6788 19230 6960 19236
rect 6736 19178 6788 19184
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 15706 5488 15914
rect 5552 15706 5580 16594
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5276 15434 5304 15642
rect 5460 15502 5488 15642
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 4764 14980 4844 15008
rect 4712 14962 4764 14968
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14550 4476 14758
rect 4724 14618 4752 14962
rect 4908 14822 4936 15030
rect 5552 14958 5580 15302
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4356 13394 4384 13670
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4252 12300 4304 12306
rect 4356 12288 4384 13330
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4448 12374 4476 12718
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4304 12260 4384 12288
rect 4252 12242 4304 12248
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3698 9959 3754 9968
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 4172 9654 4200 12242
rect 4356 11694 4384 12260
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4816 11694 4844 12786
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4264 11218 4476 11234
rect 4264 11212 4488 11218
rect 4264 11206 4436 11212
rect 4264 10130 4292 11206
rect 4436 11154 4488 11160
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4816 10810 4844 11630
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4908 9450 4936 14758
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 9178 4936 9386
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3344 5234 3372 6870
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3330 5128 3386 5137
rect 3330 5063 3386 5072
rect 3344 4842 3372 5063
rect 3436 5030 3464 6326
rect 3620 6254 3648 8502
rect 3804 8294 3832 8502
rect 3896 8430 3924 8774
rect 4080 8498 4108 8774
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3712 6866 3740 7278
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3344 4814 3464 4842
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3068 2922 3096 3130
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 3068 2446 3096 2858
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2962 640 3018 649
rect 2792 598 2912 626
rect 2884 480 2912 598
rect 2962 575 3018 584
rect 3344 480 3372 3878
rect 3436 3505 3464 4814
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3528 2854 3556 6122
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3620 2009 3648 6190
rect 3606 2000 3662 2009
rect 3606 1935 3662 1944
rect 3712 1057 3740 6258
rect 3804 5846 3832 8230
rect 4080 8129 4108 8230
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 3974 7712 4030 7721
rect 3974 7647 4030 7656
rect 3988 6934 4016 7647
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 7177 4108 7210
rect 4264 7206 4292 7822
rect 4252 7200 4304 7206
rect 4066 7168 4122 7177
rect 4252 7142 4304 7148
rect 4066 7103 4122 7112
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4066 6760 4122 6769
rect 3884 6724 3936 6730
rect 4066 6695 4122 6704
rect 3884 6666 3936 6672
rect 3896 6322 3924 6666
rect 4080 6662 4108 6695
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 4066 6216 4122 6225
rect 4172 6202 4200 6938
rect 4264 6934 4292 7142
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4122 6174 4200 6202
rect 4066 6151 4122 6160
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3698 1048 3754 1057
rect 3698 983 3754 992
rect 3804 480 3832 5646
rect 3988 5522 4016 6054
rect 4356 5930 4384 8978
rect 4903 8968 4955 8974
rect 5000 8956 5028 11086
rect 5184 11082 5212 12582
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4955 8928 5028 8956
rect 4903 8910 4955 8916
rect 4908 8894 4943 8910
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4172 5902 4384 5930
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5642 4108 5743
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3988 5494 4108 5522
rect 4080 5273 4108 5494
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3896 5166 3924 5199
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 2553 3924 4966
rect 4080 4826 4108 5034
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 4080 4078 4108 4383
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 4080 3670 4108 3839
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3988 2990 4016 3538
rect 4066 3496 4122 3505
rect 4066 3431 4068 3440
rect 4120 3431 4122 3440
rect 4068 3402 4120 3408
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3988 2582 4016 2790
rect 3976 2576 4028 2582
rect 3882 2544 3938 2553
rect 3976 2518 4028 2524
rect 3882 2479 3938 2488
rect 3976 1624 4028 1630
rect 3974 1592 3976 1601
rect 4028 1592 4030 1601
rect 3974 1527 4030 1536
rect 4172 1034 4200 5902
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 2514 4292 5510
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4632 3602 4660 4150
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1306 4844 8298
rect 4908 8090 4936 8894
rect 4896 8084 4948 8090
rect 4948 8044 5028 8072
rect 4896 8026 4948 8032
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4486 4936 5170
rect 5000 4690 5028 8044
rect 5092 6458 5120 9998
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5184 8634 5212 9318
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4214 4936 4422
rect 5000 4282 5028 4626
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4908 3602 4936 4150
rect 5092 3942 5120 4966
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5276 3754 5304 14214
rect 5552 13938 5580 14214
rect 5828 13938 5856 14486
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13462 5672 13670
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5552 11694 5580 12106
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 9110 5396 9522
rect 5460 9518 5488 9862
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 6322 5396 8570
rect 5552 7954 5580 8978
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 6656 5500 6662
rect 5552 6644 5580 7890
rect 5500 6616 5580 6644
rect 5448 6598 5500 6604
rect 5552 6322 5580 6616
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5368 5710 5396 6258
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5914 5580 6054
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5552 5234 5580 5578
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5644 4808 5672 12582
rect 5736 9722 5764 13806
rect 5828 13530 5856 13874
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5998 11792 6054 11801
rect 5998 11727 6054 11736
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5092 3726 5304 3754
rect 5552 4780 5672 4808
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4724 1278 4844 1306
rect 4172 1006 4292 1034
rect 4264 480 4292 1006
rect 4724 480 4752 1278
rect 5092 480 5120 3726
rect 5552 480 5580 4780
rect 5828 3210 5856 11630
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11286 5948 11494
rect 6012 11286 6040 11727
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9110 6040 9998
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6012 8498 6040 9046
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 8090 6040 8434
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6012 5846 6040 6190
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 3466 6040 4626
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5828 3182 6040 3210
rect 6196 3194 6224 17682
rect 7024 17542 7052 20198
rect 7116 18766 7144 20402
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 19990 8248 20198
rect 9784 19990 9812 20334
rect 10888 20058 10916 20334
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 8208 19984 8260 19990
rect 9772 19984 9824 19990
rect 8208 19926 8260 19932
rect 8666 19952 8722 19961
rect 8300 19916 8352 19922
rect 9772 19926 9824 19932
rect 11256 19922 11284 20266
rect 12544 20058 12572 20878
rect 12820 20602 12848 20946
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 8666 19887 8722 19896
rect 8760 19916 8812 19922
rect 8300 19858 8352 19864
rect 8312 19514 8340 19858
rect 8680 19854 8708 19887
rect 8760 19858 8812 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8588 19718 8616 19790
rect 8772 19786 8800 19858
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7104 18216 7156 18222
rect 7208 18204 7236 18702
rect 7156 18176 7236 18204
rect 7104 18158 7156 18164
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6840 16046 6868 17070
rect 6932 16726 6960 17070
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6920 16584 6972 16590
rect 7116 16572 7144 18158
rect 7300 17882 7328 19110
rect 7484 18970 7512 19314
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7484 18154 7512 18906
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 6972 16544 7144 16572
rect 6920 16526 6972 16532
rect 6932 16046 6960 16526
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6748 14346 6776 15506
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 7024 13394 7052 14962
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 11898 6316 13126
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6564 11558 6592 12650
rect 7024 12442 7052 13330
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 6866 6316 10066
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6380 4842 6408 9454
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8022 6500 9318
rect 6564 8566 6592 11494
rect 6932 11354 6960 12242
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6840 10266 6868 11290
rect 7116 10674 7144 11630
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6748 7954 6776 8026
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6840 7478 6868 8298
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6186 6960 7278
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6380 4814 6500 4842
rect 6012 480 6040 3182
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6472 480 6500 4814
rect 6656 4486 6684 5238
rect 6840 4826 6868 5714
rect 6932 5370 6960 5714
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6840 4026 6868 4762
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4146 6960 4422
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6748 3998 6868 4026
rect 6748 3602 6776 3998
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6564 2990 6592 3334
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6840 2514 6868 3334
rect 6932 2650 6960 3470
rect 7024 2961 7052 7142
rect 7116 6186 7144 7346
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7116 5574 7144 6122
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7116 3738 7144 4150
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7010 2952 7066 2961
rect 7010 2887 7066 2896
rect 7024 2854 7052 2887
rect 7012 2848 7064 2854
rect 7208 2802 7236 14282
rect 7300 13802 7328 14758
rect 7392 14006 7420 14894
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7392 13530 7420 13942
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7378 13424 7434 13433
rect 7378 13359 7434 13368
rect 7392 12442 7420 13359
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7392 9518 7420 11018
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8838 7420 9318
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8430 7420 8774
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7750 7420 8366
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7392 7324 7420 7686
rect 7484 7426 7512 17682
rect 7576 17678 7604 18838
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 14482 7604 14758
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 12782 7604 14418
rect 7668 13569 7696 19450
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8312 17814 8340 18090
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8312 16726 8340 16934
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8404 16658 8432 18022
rect 8496 17610 8524 19246
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8956 17746 8984 18770
rect 9508 17882 9536 19110
rect 9692 18970 9720 19110
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9784 18630 9812 19110
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9784 17746 9812 18158
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7746 15736 7802 15745
rect 7886 15728 8182 15748
rect 7746 15671 7748 15680
rect 7800 15671 7802 15680
rect 7748 15642 7800 15648
rect 8220 15570 8248 16526
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 15978 8340 16390
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8404 15502 8432 16594
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8208 14816 8260 14822
rect 7746 14784 7802 14793
rect 8208 14758 8260 14764
rect 7746 14719 7802 14728
rect 7760 14618 7788 14719
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8220 14618 8248 14758
rect 8496 14618 8524 15846
rect 8772 15026 8800 15846
rect 8864 15366 8892 15846
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 14074 7788 14350
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7654 13560 7710 13569
rect 7654 13495 7710 13504
rect 7760 13410 7788 14010
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13530 8248 14418
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13530 8432 13670
rect 8496 13530 8524 14282
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 7656 13388 7708 13394
rect 7760 13382 7880 13410
rect 7656 13330 7708 13336
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7668 11082 7696 13330
rect 7852 12782 7880 13382
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 11762 8248 12650
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8312 11354 8340 12174
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11354 8432 11494
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8496 8838 8524 13466
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11150 8616 11630
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 10266 8616 10406
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9518 8616 9998
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7546 7788 7890
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7484 7398 7788 7426
rect 7564 7336 7616 7342
rect 7392 7296 7564 7324
rect 7564 7278 7616 7284
rect 7472 6860 7524 6866
rect 7576 6848 7604 7278
rect 7524 6820 7604 6848
rect 7472 6802 7524 6808
rect 7484 6254 7512 6802
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3602 7512 4082
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7576 3534 7604 4626
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7012 2790 7064 2796
rect 7107 2774 7236 2802
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7107 2666 7135 2774
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7024 2638 7135 2666
rect 7300 2650 7328 2790
rect 7288 2644 7340 2650
rect 7024 2530 7052 2638
rect 7288 2586 7340 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6932 2502 7052 2530
rect 6932 480 6960 2502
rect 7392 480 7420 3130
rect 7484 2310 7512 3334
rect 7576 3058 7604 3470
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7668 2514 7696 4422
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7760 1306 7788 7398
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8220 4826 8248 7278
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4616 8168 4622
rect 8114 4584 8116 4593
rect 8208 4616 8260 4622
rect 8168 4584 8170 4593
rect 8208 4558 8260 4564
rect 8114 4519 8170 4528
rect 8128 4146 8156 4519
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 2938 8156 3538
rect 8220 3058 8248 4558
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8128 2910 8248 2938
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 2446 8248 2910
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7760 1278 7880 1306
rect 7852 480 7880 1278
rect 8312 480 8340 7754
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 5914 8432 7686
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8496 5370 8524 7822
rect 8588 6866 8616 7822
rect 8680 7392 8708 14758
rect 8772 13802 8800 14962
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8772 13326 8800 13738
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8758 12336 8814 12345
rect 8758 12271 8814 12280
rect 8772 11558 8800 12271
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 9382 8892 10610
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8864 8430 8892 9318
rect 8956 8430 8984 17682
rect 9784 17626 9812 17682
rect 9784 17598 9904 17626
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9784 17202 9812 17274
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 11694 9168 12582
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9232 11336 9260 15506
rect 9600 12714 9628 15982
rect 9692 14482 9720 16730
rect 9784 16250 9812 17002
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9876 16046 9904 17598
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9968 15706 9996 16934
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 12306 9720 12650
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9140 11308 9260 11336
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8680 7364 8800 7392
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6458 8616 6802
rect 8680 6662 8708 7210
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8588 5234 8616 6394
rect 8680 5710 8708 6598
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8404 3738 8432 5034
rect 8680 4758 8708 5034
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8772 480 8800 7364
rect 9048 7342 9076 8230
rect 9140 7818 9168 11308
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8864 5846 8892 6870
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5166 8892 5646
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5234 8984 5510
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8852 5024 8904 5030
rect 8904 4984 8984 5012
rect 8852 4966 8904 4972
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8864 3058 8892 4762
rect 8956 4729 8984 4984
rect 8942 4720 8998 4729
rect 8942 4655 8998 4664
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9232 480 9260 11154
rect 9416 10062 9444 11698
rect 9508 11354 9536 12242
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11898 9720 12106
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9586 10432 9642 10441
rect 9692 10418 9720 10474
rect 9642 10390 9720 10418
rect 9586 10367 9642 10376
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9926 9444 9998
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9692 9178 9720 10066
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9324 8537 9352 8570
rect 9310 8528 9366 8537
rect 9416 8498 9444 8774
rect 9310 8463 9366 8472
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 5914 9444 8434
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 6390 9536 8298
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9600 3942 9628 7958
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9692 6322 9720 6870
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9692 3602 9720 5714
rect 9784 3738 9812 15302
rect 10060 15162 10088 19722
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10336 16674 10364 17138
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10152 16646 10364 16674
rect 10428 16658 10456 16934
rect 10416 16652 10468 16658
rect 10152 15978 10180 16646
rect 10416 16594 10468 16600
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15706 10180 15914
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10336 13530 10364 14758
rect 10428 14074 10456 14758
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10428 13462 10456 13670
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10520 12986 10548 19858
rect 10968 19848 11020 19854
rect 11020 19808 11192 19836
rect 10968 19790 11020 19796
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10612 16658 10640 18770
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18154 11100 18702
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 17882 11100 18090
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11164 17746 11192 19808
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 12452 19514 12480 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12636 19446 12664 20334
rect 13648 19786 13676 20742
rect 13924 20602 13952 20810
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13740 19990 13768 20334
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 17236 19922 17264 22520
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 11440 18902 11468 19314
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12820 18970 12848 19110
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11440 18612 11468 18838
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 11256 18584 11468 18612
rect 11980 18624 12032 18630
rect 11256 18426 11284 18584
rect 11980 18566 12032 18572
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10704 17338 10732 17682
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10704 16794 10732 17274
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 10612 15434 10640 16594
rect 11164 16182 11192 16594
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11716 16046 11744 17002
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13734 10640 13806
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10612 12866 10640 13670
rect 10428 12838 10640 12866
rect 10428 12356 10456 12838
rect 10704 12356 10732 15574
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 15162 11284 15370
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11900 15162 11928 15506
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11256 14550 11284 15098
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11164 12850 11192 13330
rect 11256 13326 11284 14486
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11716 13938 11744 14418
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13530 11744 13874
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11808 12986 11836 14894
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10336 12328 10456 12356
rect 10520 12328 10732 12356
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9876 10606 9904 11834
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 10060 11558 10088 11591
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 10810 10272 11494
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 8634 9996 10134
rect 10336 9874 10364 12328
rect 10520 10470 10548 12328
rect 10980 11898 11008 12582
rect 11164 12102 11192 12786
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11256 11762 11284 12310
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11060 11688 11112 11694
rect 11152 11688 11204 11694
rect 11060 11630 11112 11636
rect 11150 11656 11152 11665
rect 11204 11656 11206 11665
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10414 10024 10470 10033
rect 10414 9959 10416 9968
rect 10468 9959 10470 9968
rect 10416 9930 10468 9936
rect 10336 9846 10456 9874
rect 10428 8634 10456 9846
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 4049 9904 6734
rect 10060 6322 10088 7686
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5778 10088 6258
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10152 4808 10180 8570
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7206 10272 7890
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 6798 10272 7142
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10428 6254 10456 7414
rect 10520 7188 10548 10406
rect 10612 9654 10640 11494
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10782 10704 10838 10713
rect 10782 10639 10784 10648
rect 10836 10639 10838 10648
rect 10784 10610 10836 10616
rect 10796 10198 10824 10610
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10796 9586 10824 10134
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10796 8498 10824 9522
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10600 7200 10652 7206
rect 10520 7160 10600 7188
rect 10600 7142 10652 7148
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5710 10456 6190
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10152 4780 10272 4808
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10152 4282 10180 4558
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9862 4040 9918 4049
rect 9862 3975 9918 3984
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 2922 9812 3538
rect 9876 3194 9904 3975
rect 9968 3602 9996 4082
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9968 3097 9996 3538
rect 10060 3398 10088 4082
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10152 3194 10180 3674
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9954 3088 10010 3097
rect 9954 3023 10010 3032
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9586 2680 9642 2689
rect 9586 2615 9642 2624
rect 9600 480 9628 2615
rect 9692 2310 9720 2858
rect 10048 2848 10100 2854
rect 10046 2816 10048 2825
rect 10100 2816 10102 2825
rect 10046 2751 10102 2760
rect 10244 2666 10272 4780
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 3738 10364 4558
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10060 2638 10272 2666
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10060 480 10088 2638
rect 10336 1630 10364 3334
rect 10428 2650 10456 4626
rect 10612 3398 10640 7142
rect 10888 4282 10916 11154
rect 11072 10470 11100 11630
rect 11150 11591 11206 11600
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10980 3942 11008 9454
rect 11072 9178 11100 10202
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 7750 11100 8978
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11072 5098 11100 5850
rect 11164 5114 11192 11494
rect 11716 11218 11744 12242
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11716 10606 11744 11018
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11716 8634 11744 9114
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11256 7410 11284 8026
rect 11716 7954 11744 8570
rect 11808 8430 11836 12922
rect 11992 12458 12020 18566
rect 12636 18290 12664 18770
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12728 18222 12756 18566
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12728 17202 12756 18158
rect 12912 17338 12940 19110
rect 13004 17882 13032 19178
rect 14016 18086 14044 19314
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20720 19168 20772 19174
rect 19246 19136 19302 19145
rect 14817 19068 15113 19088
rect 20720 19110 20772 19116
rect 19246 19071 19302 19080
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 19260 18086 19288 19071
rect 20732 18426 20760 19110
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14958 12480 15030
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 14618 12388 14826
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 11891 12430 12020 12458
rect 11891 12356 11919 12430
rect 11891 12328 11928 12356
rect 11900 9654 11928 12328
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11900 6798 11928 7686
rect 11992 7206 12020 10406
rect 12084 9654 12112 11834
rect 12268 10810 12296 12718
rect 12912 11898 12940 16934
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12176 8922 12204 9590
rect 12268 9042 12296 10746
rect 12360 10606 12388 11154
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 10266 12388 10542
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 10033 12480 10066
rect 12438 10024 12494 10033
rect 12820 9994 12848 11154
rect 12438 9959 12494 9968
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9586 12940 9862
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12176 8894 12296 8922
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8022 12204 8774
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12176 7410 12204 7958
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 12268 6474 12296 8894
rect 12176 6446 12296 6474
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11348 5914 11376 6054
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11532 5846 11560 6054
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11256 5234 11284 5782
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11060 5092 11112 5098
rect 11164 5086 11284 5114
rect 11060 5034 11112 5040
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10324 1624 10376 1630
rect 10324 1566 10376 1572
rect 10520 480 10548 3130
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10704 1306 10732 3062
rect 10980 2310 11008 3674
rect 11164 2514 11192 4966
rect 11256 2689 11284 5086
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11242 2680 11298 2689
rect 11242 2615 11298 2624
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11256 2378 11560 2394
rect 11244 2372 11572 2378
rect 11296 2366 11520 2372
rect 11244 2314 11296 2320
rect 11520 2314 11572 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 1986 11744 6054
rect 12176 4672 12204 6446
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12084 4644 12204 4672
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11900 3602 11928 3975
rect 11978 3768 12034 3777
rect 11978 3703 12034 3712
rect 11992 3670 12020 3703
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12084 3482 12112 4644
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11900 3454 12112 3482
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 2582 11836 3334
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11440 1958 11744 1986
rect 10704 1278 11008 1306
rect 10980 480 11008 1278
rect 11440 480 11468 1958
rect 11900 480 11928 3454
rect 12176 2582 12204 4490
rect 12268 3670 12296 6326
rect 12360 6118 12388 9522
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12452 6934 12480 7142
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12636 6798 12664 7142
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12728 6746 12756 7278
rect 12728 6718 12848 6746
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6254 12572 6598
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 4622 12388 5714
rect 12532 5568 12584 5574
rect 12716 5568 12768 5574
rect 12584 5516 12664 5522
rect 12532 5510 12664 5516
rect 12716 5510 12768 5516
rect 12544 5494 12664 5510
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12452 4486 12480 4762
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12268 3194 12296 3606
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12360 480 12388 3878
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12452 2650 12480 3130
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12544 1018 12572 4150
rect 12636 3602 12664 5494
rect 12728 4758 12756 5510
rect 12820 5114 12848 6718
rect 12912 5234 12940 7278
rect 13096 5778 13124 8434
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12820 5086 12940 5114
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12728 4214 12756 4694
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12716 4072 12768 4078
rect 12768 4020 12848 4026
rect 12716 4014 12848 4020
rect 12728 3998 12848 4014
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12820 3058 12848 3998
rect 12912 3942 12940 5086
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3097 13032 3470
rect 13188 3194 13216 15846
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 13268 11552 13320 11558
rect 20444 11552 20496 11558
rect 13268 11494 13320 11500
rect 19706 11520 19762 11529
rect 13280 7002 13308 11494
rect 14817 11452 15113 11472
rect 20444 11494 20496 11500
rect 19706 11455 19762 11464
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 10736 13872 10742
rect 13818 10704 13820 10713
rect 13872 10704 13874 10713
rect 13818 10639 13874 10648
rect 13924 10554 13952 10950
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 13556 10538 13952 10554
rect 13544 10532 13952 10538
rect 13596 10526 13952 10532
rect 13544 10474 13596 10480
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 6322 13400 9998
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9178 13492 9318
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13464 7750 13492 8298
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 6798 13492 7686
rect 13740 7342 13768 10406
rect 13924 9586 13952 10526
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14752 9382 14780 10610
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 14924 9512 14976 9518
rect 15212 9466 15240 9998
rect 14976 9460 15240 9466
rect 14924 9454 15240 9460
rect 14936 9438 15240 9454
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13832 6458 13860 6734
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13924 6254 13952 7210
rect 14016 6730 14044 7278
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12990 3088 13046 3097
rect 12808 3052 12860 3058
rect 12990 3023 12992 3032
rect 12808 2994 12860 3000
rect 13044 3023 13046 3032
rect 12992 2994 13044 3000
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12636 2650 12664 2926
rect 13174 2816 13230 2825
rect 13174 2751 13230 2760
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13188 2446 13216 2751
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12532 1012 12584 1018
rect 12532 954 12584 960
rect 12820 480 12848 2246
rect 13280 480 13308 3334
rect 13372 3058 13400 5238
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13648 4282 13676 4762
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 3602 13768 4626
rect 13924 4486 13952 5034
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 4146 13952 4422
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14200 4078 14228 7822
rect 14476 7342 14504 8570
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 8022 14596 8230
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 13818 3768 13874 3777
rect 13818 3703 13874 3712
rect 14096 3732 14148 3738
rect 13832 3670 13860 3703
rect 14096 3674 14148 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13832 2961 13860 3470
rect 13818 2952 13874 2961
rect 13728 2916 13780 2922
rect 13818 2887 13874 2896
rect 13728 2858 13780 2864
rect 13740 2514 13768 2858
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13728 1012 13780 1018
rect 13728 954 13780 960
rect 13740 480 13768 954
rect 14108 480 14136 3674
rect 14384 2446 14412 7210
rect 14476 6730 14504 7278
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14476 5098 14504 6666
rect 14568 6322 14596 7958
rect 14660 6866 14688 9046
rect 15212 8838 15240 9438
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15212 7886 15240 8774
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15212 6610 15240 7822
rect 15304 6730 15332 8366
rect 15856 7002 15884 11086
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 16040 9042 16068 10678
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16132 9722 16160 10066
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16132 8974 16160 9658
rect 16224 9178 16252 10406
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16316 9178 16344 9386
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 7954 16528 8910
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 7342 16068 7686
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 16040 6798 16068 7278
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15212 6582 15332 6610
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14476 4554 14504 5034
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14568 3058 14596 4966
rect 14660 3194 14688 5306
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14568 480 14596 2790
rect 14752 2650 14780 6122
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14936 5370 14964 5714
rect 15304 5710 15332 6582
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15304 5166 15332 5646
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14924 3120 14976 3126
rect 14922 3088 14924 3097
rect 14976 3088 14978 3097
rect 14922 3023 14978 3032
rect 15212 2922 15240 4014
rect 15488 3738 15516 4422
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 15304 2582 15332 3538
rect 15580 3058 15608 4558
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15672 2990 15700 3878
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15764 2514 15792 6054
rect 16132 5914 16160 6054
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16500 5574 16528 6258
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16500 5166 16528 5510
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 15856 4690 15884 5102
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 15856 3738 15884 3878
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 16224 3369 16252 3878
rect 16210 3360 16266 3369
rect 16210 3295 16266 3304
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16040 2530 16068 3130
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15948 2502 16068 2530
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 480 15056 2246
rect 15476 1488 15528 1494
rect 15476 1430 15528 1436
rect 15488 480 15516 1430
rect 15948 480 15976 2502
rect 16132 1494 16160 2790
rect 16120 1488 16172 1494
rect 16120 1430 16172 1436
rect 16408 480 16436 4082
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16500 2990 16528 3334
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16776 2582 16804 8366
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3058 16896 3538
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16960 2938 16988 8230
rect 17420 6866 17448 10950
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9110 17540 10066
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17788 6798 17816 7890
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4758 17172 4966
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17144 4214 17172 4694
rect 17788 4486 17816 5034
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17316 3936 17368 3942
rect 17696 3913 17724 3946
rect 17316 3878 17368 3884
rect 17682 3904 17738 3913
rect 16868 2910 16988 2938
rect 17224 2916 17276 2922
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16868 480 16896 2910
rect 17224 2858 17276 2864
rect 17236 2650 17264 2858
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17328 480 17356 3878
rect 17682 3839 17738 3848
rect 17788 3534 17816 4422
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17880 3380 17908 8570
rect 18064 8430 18092 9998
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 19444 9654 19472 10406
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18064 4214 18092 7142
rect 18432 6730 18460 7142
rect 18524 7002 18552 7142
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5710 18184 6190
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18156 5166 18184 5646
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4690 18184 5102
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18156 4078 18184 4626
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 4072 18196 4078
rect 17958 4040 18014 4049
rect 18144 4014 18196 4020
rect 17958 3975 17960 3984
rect 18012 3975 18014 3984
rect 17960 3946 18012 3952
rect 18418 3632 18474 3641
rect 18418 3567 18420 3576
rect 18472 3567 18474 3576
rect 18420 3538 18472 3544
rect 17788 3352 17908 3380
rect 17788 480 17816 3352
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18156 2650 18184 2790
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18248 2394 18276 2994
rect 18156 2366 18276 2394
rect 18156 1986 18184 2366
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1958 18276 1986
rect 18248 480 18276 1958
rect 18616 480 18644 8502
rect 18892 8090 18920 8978
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18708 5030 18736 5714
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18708 3534 18736 4966
rect 18800 4146 18828 7890
rect 18892 7410 18920 8026
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18892 3942 18920 5034
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18984 3058 19012 7686
rect 19076 4826 19104 8298
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19168 4706 19196 7142
rect 19352 6934 19380 8910
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19352 5574 19380 6122
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19076 4678 19196 4706
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19076 480 19104 4678
rect 19352 4622 19380 5510
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19168 3738 19196 4558
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19352 2990 19380 4422
rect 19536 3058 19564 8366
rect 19628 7342 19656 9386
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19628 4010 19656 6802
rect 19720 4078 19748 11455
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19812 7002 19840 7958
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19812 6458 19840 6734
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19904 610 19932 9590
rect 19524 604 19576 610
rect 19524 546 19576 552
rect 19892 604 19944 610
rect 19892 546 19944 552
rect 19536 480 19564 546
rect 19996 480 20024 11018
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20180 2514 20208 8434
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20272 2922 20300 5102
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20456 480 20484 11494
rect 20640 3194 20668 12038
rect 20916 7546 20944 19178
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20824 3126 20852 3878
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 21008 2666 21036 3130
rect 20916 2638 21036 2666
rect 20916 480 20944 2638
rect 21376 480 21404 3334
rect 21836 480 21864 3946
rect 22296 480 22324 7482
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22756 480 22784 2926
rect 2318 232 2374 241
rect 2318 167 2374 176
rect 2410 0 2466 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4250 0 4306 480
rect 4710 0 4766 480
rect 5078 0 5134 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8298 0 8354 480
rect 8758 0 8814 480
rect 9218 0 9274 480
rect 9586 0 9642 480
rect 10046 0 10102 480
rect 10506 0 10562 480
rect 10966 0 11022 480
rect 11426 0 11482 480
rect 11886 0 11942 480
rect 12346 0 12402 480
rect 12806 0 12862 480
rect 13266 0 13322 480
rect 13726 0 13782 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16394 0 16450 480
rect 16854 0 16910 480
rect 17314 0 17370 480
rect 17774 0 17830 480
rect 18234 0 18290 480
rect 18602 0 18658 480
rect 19062 0 19118 480
rect 19522 0 19578 480
rect 19982 0 20038 480
rect 20442 0 20498 480
rect 20902 0 20958 480
rect 21362 0 21418 480
rect 21822 0 21878 480
rect 22282 0 22338 480
rect 22742 0 22798 480
<< via2 >>
rect 4802 22616 4858 22672
rect 3790 22208 3846 22264
rect 3882 21664 3938 21720
rect 4066 21256 4122 21312
rect 3974 20712 4030 20768
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 2410 19916 2466 19952
rect 2410 19896 2412 19916
rect 2412 19896 2464 19916
rect 2464 19896 2466 19916
rect 4066 20304 4122 20360
rect 3974 19760 4030 19816
rect 3514 19352 3570 19408
rect 1582 14184 1638 14240
rect 2870 15680 2926 15736
rect 2410 14728 2466 14784
rect 3514 13232 3570 13288
rect 3422 12824 3478 12880
rect 3238 9016 3294 9072
rect 1490 4528 1546 4584
rect 2226 4800 2282 4856
rect 3146 4664 3202 4720
rect 2594 2896 2650 2952
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4066 18808 4122 18864
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4066 18400 4122 18456
rect 3974 17992 4030 18048
rect 4066 17484 4068 17504
rect 4068 17484 4120 17504
rect 4120 17484 4122 17504
rect 4066 17448 4122 17484
rect 4066 17040 4122 17096
rect 3882 16496 3938 16552
rect 4066 16088 4122 16144
rect 4066 15544 4122 15600
rect 4066 15156 4122 15192
rect 4066 15136 4068 15156
rect 4068 15136 4120 15156
rect 4120 15136 4122 15156
rect 4066 14592 4122 14648
rect 4066 13776 4122 13832
rect 3790 10920 3846 10976
rect 3698 9968 3754 10024
rect 3974 11328 4030 11384
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 3330 5072 3386 5128
rect 2962 584 3018 640
rect 3422 3440 3478 3496
rect 3606 1944 3662 2000
rect 4066 8064 4122 8120
rect 3974 7656 4030 7712
rect 4066 7112 4122 7168
rect 4066 6704 4122 6760
rect 4066 6160 4122 6216
rect 3698 992 3754 1048
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4066 5752 4122 5808
rect 3882 5208 3938 5264
rect 4066 5208 4122 5264
rect 4066 4392 4122 4448
rect 4066 3848 4122 3904
rect 4066 3460 4122 3496
rect 4066 3440 4068 3460
rect 4068 3440 4120 3460
rect 4120 3440 4122 3460
rect 3882 2488 3938 2544
rect 3974 1572 3976 1592
rect 3976 1572 4028 1592
rect 4028 1572 4030 1592
rect 3974 1536 4030 1572
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5998 11736 6054 11792
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8666 19896 8722 19952
rect 7010 2896 7066 2952
rect 7378 13368 7434 13424
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7746 15700 7802 15736
rect 7746 15680 7748 15700
rect 7748 15680 7800 15700
rect 7800 15680 7802 15700
rect 7746 14728 7802 14784
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7654 13504 7710 13560
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8114 4564 8116 4584
rect 8116 4564 8168 4584
rect 8168 4564 8170 4584
rect 8114 4528 8170 4564
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8758 12280 8814 12336
rect 8942 4664 8998 4720
rect 9586 10376 9642 10432
rect 9310 8472 9366 8528
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10046 11600 10102 11656
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11150 11636 11152 11656
rect 11152 11636 11204 11656
rect 11204 11636 11206 11656
rect 10414 9988 10470 10024
rect 10414 9968 10416 9988
rect 10416 9968 10468 9988
rect 10468 9968 10470 9988
rect 10782 10668 10838 10704
rect 10782 10648 10784 10668
rect 10784 10648 10836 10668
rect 10836 10648 10838 10668
rect 9862 3984 9918 4040
rect 9954 3032 10010 3088
rect 9586 2624 9642 2680
rect 10046 2796 10048 2816
rect 10048 2796 10100 2816
rect 10100 2796 10102 2816
rect 10046 2760 10102 2796
rect 11150 11600 11206 11636
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 19246 19080 19302 19136
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 12438 9968 12494 10024
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11242 2624 11298 2680
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11886 3984 11942 4040
rect 11978 3712 12034 3768
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 19706 11464 19762 11520
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 13818 10684 13820 10704
rect 13820 10684 13872 10704
rect 13872 10684 13874 10704
rect 13818 10648 13874 10684
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 12990 3052 13046 3088
rect 12990 3032 12992 3052
rect 12992 3032 13044 3052
rect 13044 3032 13046 3052
rect 13174 2760 13230 2816
rect 13818 3712 13874 3768
rect 13818 2896 13874 2952
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14922 3068 14924 3088
rect 14924 3068 14976 3088
rect 14976 3068 14978 3088
rect 14922 3032 14978 3068
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16210 3304 16266 3360
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 17682 3848 17738 3904
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 17958 4004 18014 4040
rect 17958 3984 17960 4004
rect 17960 3984 18012 4004
rect 18012 3984 18014 4004
rect 18418 3596 18474 3632
rect 18418 3576 18420 3596
rect 18420 3576 18472 3596
rect 18472 3576 18474 3596
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 2318 176 2374 232
<< metal3 >>
rect 0 22674 480 22704
rect 4797 22674 4863 22677
rect 0 22672 4863 22674
rect 0 22616 4802 22672
rect 4858 22616 4863 22672
rect 0 22614 4863 22616
rect 0 22584 480 22614
rect 4797 22611 4863 22614
rect 0 22266 480 22296
rect 3785 22266 3851 22269
rect 0 22264 3851 22266
rect 0 22208 3790 22264
rect 3846 22208 3851 22264
rect 0 22206 3851 22208
rect 0 22176 480 22206
rect 3785 22203 3851 22206
rect 0 21722 480 21752
rect 3877 21722 3943 21725
rect 0 21720 3943 21722
rect 0 21664 3882 21720
rect 3938 21664 3943 21720
rect 0 21662 3943 21664
rect 0 21632 480 21662
rect 3877 21659 3943 21662
rect 0 21314 480 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 480 21254
rect 4061 21251 4127 21254
rect 0 20770 480 20800
rect 3969 20770 4035 20773
rect 0 20768 4035 20770
rect 0 20712 3974 20768
rect 4030 20712 4035 20768
rect 0 20710 4035 20712
rect 0 20680 480 20710
rect 3969 20707 4035 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20362 480 20392
rect 4061 20362 4127 20365
rect 0 20360 4127 20362
rect 0 20304 4066 20360
rect 4122 20304 4127 20360
rect 0 20302 4127 20304
rect 0 20272 480 20302
rect 4061 20299 4127 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 2405 19954 2471 19957
rect 8661 19954 8727 19957
rect 2405 19952 8727 19954
rect 2405 19896 2410 19952
rect 2466 19896 8666 19952
rect 8722 19896 8727 19952
rect 2405 19894 8727 19896
rect 2405 19891 2471 19894
rect 8661 19891 8727 19894
rect 0 19818 480 19848
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19728 480 19758
rect 3969 19755 4035 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 480 19440
rect 3509 19410 3575 19413
rect 0 19408 3575 19410
rect 0 19352 3514 19408
rect 3570 19352 3575 19408
rect 0 19350 3575 19352
rect 0 19320 480 19350
rect 3509 19347 3575 19350
rect 19241 19138 19307 19141
rect 22520 19138 23000 19168
rect 19241 19136 23000 19138
rect 19241 19080 19246 19136
rect 19302 19080 23000 19136
rect 19241 19078 23000 19080
rect 19241 19075 19307 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 22520 19048 23000 19078
rect 14805 19007 15125 19008
rect 0 18866 480 18896
rect 4061 18866 4127 18869
rect 0 18864 4127 18866
rect 0 18808 4066 18864
rect 4122 18808 4127 18864
rect 0 18806 4127 18808
rect 0 18776 480 18806
rect 4061 18803 4127 18806
rect 4409 18528 4729 18529
rect 0 18458 480 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 480 18398
rect 4061 18395 4127 18398
rect 0 18050 480 18080
rect 3969 18050 4035 18053
rect 0 18048 4035 18050
rect 0 17992 3974 18048
rect 4030 17992 4035 18048
rect 0 17990 4035 17992
rect 0 17960 480 17990
rect 3969 17987 4035 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 0 17506 480 17536
rect 4061 17506 4127 17509
rect 0 17504 4127 17506
rect 0 17448 4066 17504
rect 4122 17448 4127 17504
rect 0 17446 4127 17448
rect 0 17416 480 17446
rect 4061 17443 4127 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17098 480 17128
rect 4061 17098 4127 17101
rect 0 17096 4127 17098
rect 0 17040 4066 17096
rect 4122 17040 4127 17096
rect 0 17038 4127 17040
rect 0 17008 480 17038
rect 4061 17035 4127 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 480 16584
rect 3877 16554 3943 16557
rect 0 16552 3943 16554
rect 0 16496 3882 16552
rect 3938 16496 3943 16552
rect 0 16494 3943 16496
rect 0 16464 480 16494
rect 3877 16491 3943 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 480 16176
rect 4061 16146 4127 16149
rect 0 16144 4127 16146
rect 0 16088 4066 16144
rect 4122 16088 4127 16144
rect 0 16086 4127 16088
rect 0 16056 480 16086
rect 4061 16083 4127 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 2865 15738 2931 15741
rect 7741 15738 7807 15741
rect 2865 15736 7807 15738
rect 2865 15680 2870 15736
rect 2926 15680 7746 15736
rect 7802 15680 7807 15736
rect 2865 15678 7807 15680
rect 2865 15675 2931 15678
rect 7741 15675 7807 15678
rect 0 15602 480 15632
rect 4061 15602 4127 15605
rect 0 15600 4127 15602
rect 0 15544 4066 15600
rect 4122 15544 4127 15600
rect 0 15542 4127 15544
rect 0 15512 480 15542
rect 4061 15539 4127 15542
rect 4409 15264 4729 15265
rect 0 15194 480 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 4061 15194 4127 15197
rect 0 15192 4127 15194
rect 0 15136 4066 15192
rect 4122 15136 4127 15192
rect 0 15134 4127 15136
rect 0 15104 480 15134
rect 4061 15131 4127 15134
rect 2405 14786 2471 14789
rect 7741 14786 7807 14789
rect 2405 14784 7807 14786
rect 2405 14728 2410 14784
rect 2466 14728 7746 14784
rect 7802 14728 7807 14784
rect 2405 14726 7807 14728
rect 2405 14723 2471 14726
rect 7741 14723 7807 14726
rect 7874 14720 8194 14721
rect 0 14650 480 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 4061 14650 4127 14653
rect 0 14648 4127 14650
rect 0 14592 4066 14648
rect 4122 14592 4127 14648
rect 0 14590 4127 14592
rect 0 14560 480 14590
rect 4061 14587 4127 14590
rect 0 14242 480 14272
rect 1577 14242 1643 14245
rect 0 14240 1643 14242
rect 0 14184 1582 14240
rect 1638 14184 1643 14240
rect 0 14182 1643 14184
rect 0 14152 480 14182
rect 1577 14179 1643 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 0 13834 480 13864
rect 4061 13834 4127 13837
rect 0 13832 4127 13834
rect 0 13776 4066 13832
rect 4122 13776 4127 13832
rect 0 13774 4127 13776
rect 0 13744 480 13774
rect 4061 13771 4127 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 7649 13562 7715 13565
rect 7606 13560 7715 13562
rect 7606 13504 7654 13560
rect 7710 13504 7715 13560
rect 7606 13499 7715 13504
rect 7373 13426 7439 13429
rect 7606 13426 7666 13499
rect 7373 13424 7666 13426
rect 7373 13368 7378 13424
rect 7434 13368 7666 13424
rect 7373 13366 7666 13368
rect 7373 13363 7439 13366
rect 0 13290 480 13320
rect 3509 13290 3575 13293
rect 0 13288 3575 13290
rect 0 13232 3514 13288
rect 3570 13232 3575 13288
rect 0 13230 3575 13232
rect 0 13200 480 13230
rect 3509 13227 3575 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 480 12912
rect 3417 12882 3483 12885
rect 0 12880 3483 12882
rect 0 12824 3422 12880
rect 3478 12824 3483 12880
rect 0 12822 3483 12824
rect 0 12792 480 12822
rect 3417 12819 3483 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12338 480 12368
rect 8753 12338 8819 12341
rect 0 12336 8819 12338
rect 0 12280 8758 12336
rect 8814 12280 8819 12336
rect 0 12278 8819 12280
rect 0 12248 480 12278
rect 8753 12275 8819 12278
rect 4409 12000 4729 12001
rect 0 11930 480 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 0 11870 4170 11930
rect 0 11840 480 11870
rect 4110 11794 4170 11870
rect 5993 11794 6059 11797
rect 4110 11792 6059 11794
rect 4110 11736 5998 11792
rect 6054 11736 6059 11792
rect 4110 11734 6059 11736
rect 5993 11731 6059 11734
rect 10041 11658 10107 11661
rect 11145 11658 11211 11661
rect 10041 11656 11211 11658
rect 10041 11600 10046 11656
rect 10102 11600 11150 11656
rect 11206 11600 11211 11656
rect 10041 11598 11211 11600
rect 10041 11595 10107 11598
rect 11145 11595 11211 11598
rect 19701 11522 19767 11525
rect 22520 11522 23000 11552
rect 19701 11520 23000 11522
rect 19701 11464 19706 11520
rect 19762 11464 23000 11520
rect 19701 11462 23000 11464
rect 19701 11459 19767 11462
rect 7874 11456 8194 11457
rect 0 11386 480 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 22520 11432 23000 11462
rect 14805 11391 15125 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 480 11326
rect 3969 11323 4035 11326
rect 0 10978 480 11008
rect 3785 10978 3851 10981
rect 0 10976 3851 10978
rect 0 10920 3790 10976
rect 3846 10920 3851 10976
rect 0 10918 3851 10920
rect 0 10888 480 10918
rect 3785 10915 3851 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 10777 10706 10843 10709
rect 13813 10706 13879 10709
rect 10777 10704 13879 10706
rect 10777 10648 10782 10704
rect 10838 10648 13818 10704
rect 13874 10648 13879 10704
rect 10777 10646 13879 10648
rect 10777 10643 10843 10646
rect 13813 10643 13879 10646
rect 4846 10510 8402 10570
rect 0 10434 480 10464
rect 4846 10434 4906 10510
rect 0 10374 4906 10434
rect 8342 10434 8402 10510
rect 9581 10434 9647 10437
rect 8342 10432 9647 10434
rect 8342 10376 9586 10432
rect 9642 10376 9647 10432
rect 8342 10374 9647 10376
rect 0 10344 480 10374
rect 9581 10371 9647 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 0 10026 480 10056
rect 3693 10026 3759 10029
rect 0 10024 3759 10026
rect 0 9968 3698 10024
rect 3754 9968 3759 10024
rect 0 9966 3759 9968
rect 0 9936 480 9966
rect 3693 9963 3759 9966
rect 10409 10026 10475 10029
rect 12433 10026 12499 10029
rect 10409 10024 12499 10026
rect 10409 9968 10414 10024
rect 10470 9968 12438 10024
rect 12494 9968 12499 10024
rect 10409 9966 12499 9968
rect 10409 9963 10475 9966
rect 12433 9963 12499 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 0 9482 480 9512
rect 9438 9482 9444 9484
rect 0 9422 9444 9482
rect 0 9392 480 9422
rect 9438 9420 9444 9422
rect 9508 9420 9514 9484
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 480 9104
rect 3233 9074 3299 9077
rect 0 9072 3299 9074
rect 0 9016 3238 9072
rect 3294 9016 3299 9072
rect 0 9014 3299 9016
rect 0 8984 480 9014
rect 3233 9011 3299 9014
rect 4409 8736 4729 8737
rect 0 8666 480 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 0 8606 4170 8666
rect 0 8576 480 8606
rect 4110 8530 4170 8606
rect 9305 8530 9371 8533
rect 4110 8528 9371 8530
rect 4110 8472 9310 8528
rect 9366 8472 9371 8528
rect 4110 8470 9371 8472
rect 9305 8467 9371 8470
rect 7874 8192 8194 8193
rect 0 8122 480 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 0 7714 480 7744
rect 3969 7714 4035 7717
rect 0 7712 4035 7714
rect 0 7656 3974 7712
rect 4030 7656 4035 7712
rect 0 7654 4035 7656
rect 0 7624 480 7654
rect 3969 7651 4035 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 480 5296
rect 3877 5266 3943 5269
rect 0 5264 3943 5266
rect 0 5208 3882 5264
rect 3938 5208 3943 5264
rect 0 5206 3943 5208
rect 0 5176 480 5206
rect 3877 5203 3943 5206
rect 4061 5266 4127 5269
rect 4061 5264 4170 5266
rect 4061 5208 4066 5264
rect 4122 5208 4170 5264
rect 4061 5203 4170 5208
rect 3325 5130 3391 5133
rect 4110 5130 4170 5203
rect 3325 5128 4170 5130
rect 3325 5072 3330 5128
rect 3386 5072 4170 5128
rect 3325 5070 4170 5072
rect 3325 5067 3391 5070
rect 7874 4928 8194 4929
rect 0 4858 480 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 2221 4858 2287 4861
rect 0 4856 2287 4858
rect 0 4800 2226 4856
rect 2282 4800 2287 4856
rect 0 4798 2287 4800
rect 0 4768 480 4798
rect 2221 4795 2287 4798
rect 3141 4722 3207 4725
rect 8937 4722 9003 4725
rect 3141 4720 9003 4722
rect 3141 4664 3146 4720
rect 3202 4664 8942 4720
rect 8998 4664 9003 4720
rect 3141 4662 9003 4664
rect 3141 4659 3207 4662
rect 8937 4659 9003 4662
rect 1485 4586 1551 4589
rect 8109 4586 8175 4589
rect 1485 4584 8175 4586
rect 1485 4528 1490 4584
rect 1546 4528 8114 4584
rect 8170 4528 8175 4584
rect 1485 4526 8175 4528
rect 1485 4523 1551 4526
rect 8109 4523 8175 4526
rect 0 4450 480 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 480 4390
rect 4061 4387 4127 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 9857 4042 9923 4045
rect 11881 4042 11947 4045
rect 17953 4042 18019 4045
rect 9857 4040 18019 4042
rect 9857 3984 9862 4040
rect 9918 3984 11886 4040
rect 11942 3984 17958 4040
rect 18014 3984 18019 4040
rect 9857 3982 18019 3984
rect 9857 3979 9923 3982
rect 11881 3979 11947 3982
rect 17953 3979 18019 3982
rect 0 3906 480 3936
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 480 3846
rect 4061 3843 4127 3846
rect 17677 3906 17743 3909
rect 22520 3906 23000 3936
rect 17677 3904 23000 3906
rect 17677 3848 17682 3904
rect 17738 3848 23000 3904
rect 17677 3846 23000 3848
rect 17677 3843 17743 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22520 3816 23000 3846
rect 14805 3775 15125 3776
rect 11973 3770 12039 3773
rect 13813 3770 13879 3773
rect 11973 3768 13879 3770
rect 11973 3712 11978 3768
rect 12034 3712 13818 3768
rect 13874 3712 13879 3768
rect 11973 3710 13879 3712
rect 11973 3707 12039 3710
rect 13813 3707 13879 3710
rect 9438 3572 9444 3636
rect 9508 3634 9514 3636
rect 18413 3634 18479 3637
rect 9508 3632 18479 3634
rect 9508 3576 18418 3632
rect 18474 3576 18479 3632
rect 9508 3574 18479 3576
rect 9508 3572 9514 3574
rect 18413 3571 18479 3574
rect 0 3498 480 3528
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3408 480 3438
rect 3417 3435 3483 3438
rect 4061 3498 4127 3501
rect 4061 3496 12266 3498
rect 4061 3440 4066 3496
rect 4122 3440 12266 3496
rect 4061 3438 12266 3440
rect 4061 3435 4127 3438
rect 12206 3362 12266 3438
rect 16205 3362 16271 3365
rect 12206 3360 16271 3362
rect 12206 3304 16210 3360
rect 16266 3304 16271 3360
rect 12206 3302 16271 3304
rect 16205 3299 16271 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 9949 3090 10015 3093
rect 12985 3090 13051 3093
rect 14917 3090 14983 3093
rect 9949 3088 14983 3090
rect 9949 3032 9954 3088
rect 10010 3032 12990 3088
rect 13046 3032 14922 3088
rect 14978 3032 14983 3088
rect 9949 3030 14983 3032
rect 9949 3027 10015 3030
rect 12985 3027 13051 3030
rect 14917 3027 14983 3030
rect 0 2954 480 2984
rect 2589 2954 2655 2957
rect 0 2952 2655 2954
rect 0 2896 2594 2952
rect 2650 2896 2655 2952
rect 0 2894 2655 2896
rect 0 2864 480 2894
rect 2589 2891 2655 2894
rect 7005 2954 7071 2957
rect 13813 2954 13879 2957
rect 7005 2952 13879 2954
rect 7005 2896 7010 2952
rect 7066 2896 13818 2952
rect 13874 2896 13879 2952
rect 7005 2894 13879 2896
rect 7005 2891 7071 2894
rect 13813 2891 13879 2894
rect 10041 2818 10107 2821
rect 13169 2818 13235 2821
rect 10041 2816 13235 2818
rect 10041 2760 10046 2816
rect 10102 2760 13174 2816
rect 13230 2760 13235 2816
rect 10041 2758 13235 2760
rect 10041 2755 10107 2758
rect 13169 2755 13235 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 9581 2682 9647 2685
rect 11237 2682 11303 2685
rect 9581 2680 11303 2682
rect 9581 2624 9586 2680
rect 9642 2624 11242 2680
rect 11298 2624 11303 2680
rect 9581 2622 11303 2624
rect 9581 2619 9647 2622
rect 11237 2619 11303 2622
rect 0 2546 480 2576
rect 3877 2546 3943 2549
rect 0 2544 3943 2546
rect 0 2488 3882 2544
rect 3938 2488 3943 2544
rect 0 2486 3943 2488
rect 0 2456 480 2486
rect 3877 2483 3943 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 480 2032
rect 3601 2002 3667 2005
rect 0 2000 3667 2002
rect 0 1944 3606 2000
rect 3662 1944 3667 2000
rect 0 1942 3667 1944
rect 0 1912 480 1942
rect 3601 1939 3667 1942
rect 0 1594 480 1624
rect 3969 1594 4035 1597
rect 0 1592 4035 1594
rect 0 1536 3974 1592
rect 4030 1536 4035 1592
rect 0 1534 4035 1536
rect 0 1504 480 1534
rect 3969 1531 4035 1534
rect 0 1050 480 1080
rect 3693 1050 3759 1053
rect 0 1048 3759 1050
rect 0 992 3698 1048
rect 3754 992 3759 1048
rect 0 990 3759 992
rect 0 960 480 990
rect 3693 987 3759 990
rect 0 642 480 672
rect 2957 642 3023 645
rect 0 640 3023 642
rect 0 584 2962 640
rect 3018 584 3023 640
rect 0 582 3023 584
rect 0 552 480 582
rect 2957 579 3023 582
rect 0 234 480 264
rect 2313 234 2379 237
rect 0 232 2379 234
rect 0 176 2318 232
rect 2374 176 2379 232
rect 0 174 2379 176
rect 0 144 480 174
rect 2313 171 2379 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 9444 9420 9508 9484
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 9444 3572 9508 3636
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 9443 9484 9509 9485
rect 9443 9420 9444 9484
rect 9508 9420 9509 9484
rect 9443 9419 9509 9420
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 9446 3637 9506 9419
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 9443 3636 9509 3637
rect 9443 3572 9444 3636
rect 9508 3572 9509 3636
rect 9443 3571 9509 3572
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_20 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1604681595
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_76
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8832 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1604681595
transform 1 0 10028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _112_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15732 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1604681595
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_164
timestamp 1604681595
transform 1 0 16192 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1604681595
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_191
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204
timestamp 1604681595
transform 1 0 19872 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _071_
timestamp 1604681595
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_54
timestamp 1604681595
transform 1 0 6072 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_82
timestamp 1604681595
transform 1 0 8648 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_126
timestamp 1604681595
transform 1 0 12696 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_140
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_176
timestamp 1604681595
transform 1 0 17296 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_195
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1604681595
transform 1 0 19596 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_17
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_41
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_49
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_83
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_190
timestamp 1604681595
transform 1 0 18584 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_198
timestamp 1604681595
transform 1 0 19320 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_35
timestamp 1604681595
transform 1 0 4324 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_63
timestamp 1604681595
transform 1 0 6900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12512 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_116
timestamp 1604681595
transform 1 0 11776 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_140
timestamp 1604681595
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_182
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_200
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_16
timestamp 1604681595
transform 1 0 2576 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_47
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_88
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1604681595
transform 1 0 10304 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_151
timestamp 1604681595
transform 1 0 14996 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_200
timestamp 1604681595
transform 1 0 19504 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_212
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1656 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_22
timestamp 1604681595
transform 1 0 3128 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1604681595
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_103
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_127
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_130
timestamp 1604681595
transform 1 0 13064 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_170
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_167
timestamp 1604681595
transform 1 0 16468 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_48
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_119
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_137
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1604681595
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1604681595
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_175
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_189
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_55
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6900 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_72
timestamp 1604681595
transform 1 0 7728 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_96
timestamp 1604681595
transform 1 0 9936 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1604681595
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_146
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1604681595
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1604681595
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1604681595
transform 1 0 21068 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_19
timestamp 1604681595
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_61
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11960 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_109
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_134
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_194
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_17
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_34
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_42
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1604681595
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_88
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1604681595
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_162
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 16744 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_211
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_57
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_81
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1604681595
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_104
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17388 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_174
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_25
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7452 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_97
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_139
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_137
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_177
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_196
timestamp 1604681595
transform 1 0 19136 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_19
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6900 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_139
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 18492 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_38
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5520 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_140
timestamp 1604681595
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_199
timestamp 1604681595
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_94
timestamp 1604681595
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_200
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1604681595
transform 1 0 19964 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_6
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_38
timestamp 1604681595
transform 1 0 4600 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_72
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_133
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 1472 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_8
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_70
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_72
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 10304 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_88
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_100
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_99
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 1604681595
transform 1 0 10580 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_111
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_126
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_138
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_150
timestamp 1604681595
transform 1 0 14904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1604681595
transform 1 0 17112 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_14
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 4508 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_31
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_65
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_89
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_126
timestamp 1604681595
transform 1 0 12696 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_138
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_150
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1604681595
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_43
timestamp 1604681595
transform 1 0 5060 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_82
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_136
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1604681595
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_12
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_24
timestamp 1604681595
transform 1 0 3312 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_94
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1604681595
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1604681595
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1604681595
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_18
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1604681595
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_48
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11592 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_18
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4324 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_84
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_134
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_155
timestamp 1604681595
transform 1 0 15364 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_167
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_6
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_17
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_55
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_45
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6900 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_79
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_83
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_100
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_112
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_130
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_142
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_134
timestamp 1604681595
transform 1 0 13432 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1604681595
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1604681595
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1604681595
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_38
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_50
timestamp 1604681595
transform 1 0 5704 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 1604681595
transform 1 0 12236 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1604681595
transform 1 0 2760 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_48
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6992 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_92
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_165
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_6
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1604681595
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_104
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 13432 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_126
timestamp 1604681595
transform 1 0 12696 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_31
timestamp 1604681595
transform 1 0 3956 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1604681595
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_55
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1604681595
transform 1 0 8740 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 10672 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_96
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_108
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_144
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_168
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_17
timestamp 1604681595
transform 1 0 2668 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_38
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 6624 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5336 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_52
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1604681595
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_99
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_107
timestamp 1604681595
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_115
timestamp 1604681595
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 13524 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_127
timestamp 1604681595
transform 1 0 12788 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_139
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _070_
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_176
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_188
timestamp 1604681595
transform 1 0 18400 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_18
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_30
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_38
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 5336 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_50
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_79
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 10856 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1604681595
transform 1 0 14076 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1604681595
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_199
timestamp 1604681595
transform 1 0 19412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 22282 0 22338 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 5722 22520 5778 23000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 22742 0 22798 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 17222 22520 17278 23000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 21822 0 21878 480 6 bottom_right_grid_pin_1_
port 12 nsew default input
rlabel metal3 s 22520 11432 23000 11552 6 ccff_head
port 13 nsew default input
rlabel metal3 s 22520 19048 23000 19168 6 ccff_tail
port 14 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[10]
port 16 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 17 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 18 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 19 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 20 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[15]
port 21 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 22 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[17]
port 23 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 24 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[19]
port 25 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 26 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 27 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 28 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 29 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 30 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 31 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 32 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[8]
port 33 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 34 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 35 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[10]
port 36 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[11]
port 37 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 38 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[13]
port 39 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 40 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[15]
port 41 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[16]
port 42 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[17]
port 43 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[18]
port 44 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[19]
port 45 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[1]
port 46 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_left_out[2]
port 47 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 48 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[4]
port 49 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 50 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[6]
port 51 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 52 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[8]
port 53 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[9]
port 54 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_in[0]
port 55 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[10]
port 56 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[11]
port 57 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[12]
port 58 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[13]
port 59 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[14]
port 60 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[15]
port 61 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[16]
port 62 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[17]
port 63 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[18]
port 64 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[19]
port 65 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[1]
port 66 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[2]
port 67 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[3]
port 68 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[4]
port 69 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[5]
port 70 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[6]
port 71 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[7]
port 72 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[8]
port 73 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[9]
port 74 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_out[0]
port 75 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[10]
port 76 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[11]
port 77 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[12]
port 78 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[13]
port 79 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[14]
port 80 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[15]
port 81 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 chany_bottom_out[16]
port 82 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[17]
port 83 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[18]
port 84 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[19]
port 85 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[1]
port 86 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[2]
port 87 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[3]
port 88 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[4]
port 89 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[5]
port 90 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[6]
port 91 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[7]
port 92 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[8]
port 93 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[9]
port 94 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 95 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 96 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 97 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 98 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 99 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 100 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 101 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 102 nsew default input
rlabel metal3 s 0 22584 480 22704 6 left_top_grid_pin_1_
port 103 nsew default input
rlabel metal3 s 22520 3816 23000 3936 6 prog_clk
port 104 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 105 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 106 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
