magic
tech sky130A
magscale 1 2
timestamp 1606236529
<< viali >>
rect 5587 9129 5621 9163
rect 5403 8993 5437 9027
rect 4759 7973 4793 8007
rect 4667 7837 4701 7871
rect 5311 7837 5345 7871
rect 3195 6341 3229 6375
rect 3563 6205 3597 6239
rect 3931 6137 3965 6171
rect 5162 5729 5196 5763
rect 5265 5525 5299 5559
rect 4759 4709 4793 4743
rect 4667 4573 4701 4607
rect 5219 4573 5253 4607
rect 1631 4029 1665 4063
rect 1898 3961 1932 3995
rect 3011 3893 3045 3927
<< metal1 >>
rect 38 14714 6754 14736
rect 38 14662 2180 14714
rect 2232 14662 2244 14714
rect 2296 14662 2308 14714
rect 2360 14662 2372 14714
rect 2424 14662 4444 14714
rect 4496 14662 4508 14714
rect 4560 14662 4572 14714
rect 4624 14662 4636 14714
rect 4688 14662 6754 14714
rect 38 14640 6754 14662
rect 38 14170 6754 14192
rect 38 14118 1048 14170
rect 1100 14118 1112 14170
rect 1164 14118 1176 14170
rect 1228 14118 1240 14170
rect 1292 14118 3312 14170
rect 3364 14118 3376 14170
rect 3428 14118 3440 14170
rect 3492 14118 3504 14170
rect 3556 14118 5576 14170
rect 5628 14118 5640 14170
rect 5692 14118 5704 14170
rect 5756 14118 5768 14170
rect 5820 14118 6754 14170
rect 38 14096 6754 14118
rect 38 13626 6754 13648
rect 38 13574 2180 13626
rect 2232 13574 2244 13626
rect 2296 13574 2308 13626
rect 2360 13574 2372 13626
rect 2424 13574 4444 13626
rect 4496 13574 4508 13626
rect 4560 13574 4572 13626
rect 4624 13574 4636 13626
rect 4688 13574 6754 13626
rect 38 13552 6754 13574
rect 38 13082 6754 13104
rect 38 13030 1048 13082
rect 1100 13030 1112 13082
rect 1164 13030 1176 13082
rect 1228 13030 1240 13082
rect 1292 13030 3312 13082
rect 3364 13030 3376 13082
rect 3428 13030 3440 13082
rect 3492 13030 3504 13082
rect 3556 13030 5576 13082
rect 5628 13030 5640 13082
rect 5692 13030 5704 13082
rect 5756 13030 5768 13082
rect 5820 13030 6754 13082
rect 38 13008 6754 13030
rect 1340 12588 1346 12640
rect 1398 12628 1404 12640
rect 3180 12628 3186 12640
rect 1398 12600 3186 12628
rect 1398 12588 1404 12600
rect 3180 12588 3186 12600
rect 3238 12588 3244 12640
rect 38 12538 6754 12560
rect 38 12486 2180 12538
rect 2232 12486 2244 12538
rect 2296 12486 2308 12538
rect 2360 12486 2372 12538
rect 2424 12486 4444 12538
rect 4496 12486 4508 12538
rect 4560 12486 4572 12538
rect 4624 12486 4636 12538
rect 4688 12486 6754 12538
rect 38 12464 6754 12486
rect 38 11994 6754 12016
rect 38 11942 1048 11994
rect 1100 11942 1112 11994
rect 1164 11942 1176 11994
rect 1228 11942 1240 11994
rect 1292 11942 3312 11994
rect 3364 11942 3376 11994
rect 3428 11942 3440 11994
rect 3492 11942 3504 11994
rect 3556 11942 5576 11994
rect 5628 11942 5640 11994
rect 5692 11942 5704 11994
rect 5756 11942 5768 11994
rect 5820 11942 6754 11994
rect 38 11920 6754 11942
rect 38 11450 6754 11472
rect 38 11398 2180 11450
rect 2232 11398 2244 11450
rect 2296 11398 2308 11450
rect 2360 11398 2372 11450
rect 2424 11398 4444 11450
rect 4496 11398 4508 11450
rect 4560 11398 4572 11450
rect 4624 11398 4636 11450
rect 4688 11398 6754 11450
rect 38 11376 6754 11398
rect 38 10906 6754 10928
rect 38 10854 1048 10906
rect 1100 10854 1112 10906
rect 1164 10854 1176 10906
rect 1228 10854 1240 10906
rect 1292 10854 3312 10906
rect 3364 10854 3376 10906
rect 3428 10854 3440 10906
rect 3492 10854 3504 10906
rect 3556 10854 5576 10906
rect 5628 10854 5640 10906
rect 5692 10854 5704 10906
rect 5756 10854 5768 10906
rect 5820 10854 6754 10906
rect 38 10832 6754 10854
rect 38 10362 6754 10384
rect 38 10310 2180 10362
rect 2232 10310 2244 10362
rect 2296 10310 2308 10362
rect 2360 10310 2372 10362
rect 2424 10310 4444 10362
rect 4496 10310 4508 10362
rect 4560 10310 4572 10362
rect 4624 10310 4636 10362
rect 4688 10310 6754 10362
rect 38 10288 6754 10310
rect 38 9818 6754 9840
rect 38 9766 1048 9818
rect 1100 9766 1112 9818
rect 1164 9766 1176 9818
rect 1228 9766 1240 9818
rect 1292 9766 3312 9818
rect 3364 9766 3376 9818
rect 3428 9766 3440 9818
rect 3492 9766 3504 9818
rect 3556 9766 5576 9818
rect 5628 9766 5640 9818
rect 5692 9766 5704 9818
rect 5756 9766 5768 9818
rect 5820 9766 6754 9818
rect 38 9744 6754 9766
rect 38 9274 6754 9296
rect 38 9222 2180 9274
rect 2232 9222 2244 9274
rect 2296 9222 2308 9274
rect 2360 9222 2372 9274
rect 2424 9222 4444 9274
rect 4496 9222 4508 9274
rect 4560 9222 4572 9274
rect 4624 9222 4636 9274
rect 4688 9222 6754 9274
rect 38 9200 6754 9222
rect 5388 9120 5394 9172
rect 5446 9160 5452 9172
rect 5575 9163 5633 9169
rect 5575 9160 5587 9163
rect 5446 9132 5587 9160
rect 5446 9120 5452 9132
rect 5575 9129 5587 9132
rect 5621 9129 5633 9163
rect 5575 9123 5633 9129
rect 5388 9024 5394 9036
rect 5349 8996 5394 9024
rect 5388 8984 5394 8996
rect 5446 8984 5452 9036
rect 38 8730 6754 8752
rect 38 8678 1048 8730
rect 1100 8678 1112 8730
rect 1164 8678 1176 8730
rect 1228 8678 1240 8730
rect 1292 8678 3312 8730
rect 3364 8678 3376 8730
rect 3428 8678 3440 8730
rect 3492 8678 3504 8730
rect 3556 8678 5576 8730
rect 5628 8678 5640 8730
rect 5692 8678 5704 8730
rect 5756 8678 5768 8730
rect 5820 8678 6754 8730
rect 38 8656 6754 8678
rect 38 8186 6754 8208
rect 38 8134 2180 8186
rect 2232 8134 2244 8186
rect 2296 8134 2308 8186
rect 2360 8134 2372 8186
rect 2424 8134 4444 8186
rect 4496 8134 4508 8186
rect 4560 8134 4572 8186
rect 4624 8134 4636 8186
rect 4688 8134 6754 8186
rect 38 8112 6754 8134
rect 4284 7964 4290 8016
rect 4342 8004 4348 8016
rect 4747 8007 4805 8013
rect 4747 8004 4759 8007
rect 4342 7976 4759 8004
rect 4342 7964 4348 7976
rect 4747 7973 4759 7976
rect 4793 7973 4805 8007
rect 4747 7967 4805 7973
rect 4655 7871 4713 7877
rect 4655 7837 4667 7871
rect 4701 7868 4713 7871
rect 4744 7868 4750 7880
rect 4701 7840 4750 7868
rect 4701 7837 4713 7840
rect 4655 7831 4713 7837
rect 4744 7828 4750 7840
rect 4802 7828 4808 7880
rect 5296 7868 5302 7880
rect 5257 7840 5302 7868
rect 5296 7828 5302 7840
rect 5354 7828 5360 7880
rect 38 7642 6754 7664
rect 38 7590 1048 7642
rect 1100 7590 1112 7642
rect 1164 7590 1176 7642
rect 1228 7590 1240 7642
rect 1292 7590 3312 7642
rect 3364 7590 3376 7642
rect 3428 7590 3440 7642
rect 3492 7590 3504 7642
rect 3556 7590 5576 7642
rect 5628 7590 5640 7642
rect 5692 7590 5704 7642
rect 5756 7590 5768 7642
rect 5820 7590 6754 7642
rect 38 7568 6754 7590
rect 38 7098 6754 7120
rect 38 7046 2180 7098
rect 2232 7046 2244 7098
rect 2296 7046 2308 7098
rect 2360 7046 2372 7098
rect 2424 7046 4444 7098
rect 4496 7046 4508 7098
rect 4560 7046 4572 7098
rect 4624 7046 4636 7098
rect 4688 7046 6754 7098
rect 38 7024 6754 7046
rect 38 6554 6754 6576
rect 38 6502 1048 6554
rect 1100 6502 1112 6554
rect 1164 6502 1176 6554
rect 1228 6502 1240 6554
rect 1292 6502 3312 6554
rect 3364 6502 3376 6554
rect 3428 6502 3440 6554
rect 3492 6502 3504 6554
rect 3556 6502 5576 6554
rect 5628 6502 5640 6554
rect 5692 6502 5704 6554
rect 5756 6502 5768 6554
rect 5820 6502 6754 6554
rect 38 6480 6754 6502
rect 3180 6372 3186 6384
rect 3141 6344 3186 6372
rect 3180 6332 3186 6344
rect 3238 6332 3244 6384
rect 3551 6239 3609 6245
rect 3551 6205 3563 6239
rect 3597 6236 3609 6239
rect 3640 6236 3646 6248
rect 3597 6208 3646 6236
rect 3597 6205 3609 6208
rect 3551 6199 3609 6205
rect 3640 6196 3646 6208
rect 3698 6196 3704 6248
rect 3916 6168 3922 6180
rect 3877 6140 3922 6168
rect 3916 6128 3922 6140
rect 3974 6168 3980 6180
rect 4284 6168 4290 6180
rect 3974 6140 4290 6168
rect 3974 6128 3980 6140
rect 4284 6128 4290 6140
rect 4342 6128 4348 6180
rect 38 6010 6754 6032
rect 38 5958 2180 6010
rect 2232 5958 2244 6010
rect 2296 5958 2308 6010
rect 2360 5958 2372 6010
rect 2424 5958 4444 6010
rect 4496 5958 4508 6010
rect 4560 5958 4572 6010
rect 4624 5958 4636 6010
rect 4688 5958 6754 6010
rect 38 5936 6754 5958
rect 3916 5720 3922 5772
rect 3974 5760 3980 5772
rect 5150 5763 5208 5769
rect 5150 5760 5162 5763
rect 3974 5732 5162 5760
rect 3974 5720 3980 5732
rect 5150 5729 5162 5732
rect 5196 5729 5208 5763
rect 5150 5723 5208 5729
rect 4744 5516 4750 5568
rect 4802 5556 4808 5568
rect 5253 5559 5311 5565
rect 5253 5556 5265 5559
rect 4802 5528 5265 5556
rect 4802 5516 4808 5528
rect 5253 5525 5265 5528
rect 5299 5525 5311 5559
rect 5253 5519 5311 5525
rect 38 5466 6754 5488
rect 38 5414 1048 5466
rect 1100 5414 1112 5466
rect 1164 5414 1176 5466
rect 1228 5414 1240 5466
rect 1292 5414 3312 5466
rect 3364 5414 3376 5466
rect 3428 5414 3440 5466
rect 3492 5414 3504 5466
rect 3556 5414 5576 5466
rect 5628 5414 5640 5466
rect 5692 5414 5704 5466
rect 5756 5414 5768 5466
rect 5820 5414 6754 5466
rect 38 5392 6754 5414
rect 38 4922 6754 4944
rect 38 4870 2180 4922
rect 2232 4870 2244 4922
rect 2296 4870 2308 4922
rect 2360 4870 2372 4922
rect 2424 4870 4444 4922
rect 4496 4870 4508 4922
rect 4560 4870 4572 4922
rect 4624 4870 4636 4922
rect 4688 4870 6754 4922
rect 38 4848 6754 4870
rect 4744 4740 4750 4752
rect 4705 4712 4750 4740
rect 4744 4700 4750 4712
rect 4802 4700 4808 4752
rect 4655 4607 4713 4613
rect 4655 4573 4667 4607
rect 4701 4573 4713 4607
rect 5204 4604 5210 4616
rect 5165 4576 5210 4604
rect 4655 4567 4713 4573
rect 4670 4536 4698 4567
rect 5204 4564 5210 4576
rect 5262 4564 5268 4616
rect 6768 4536 6774 4548
rect 4670 4508 6774 4536
rect 6768 4496 6774 4508
rect 6826 4496 6832 4548
rect 38 4378 6754 4400
rect 38 4326 1048 4378
rect 1100 4326 1112 4378
rect 1164 4326 1176 4378
rect 1228 4326 1240 4378
rect 1292 4326 3312 4378
rect 3364 4326 3376 4378
rect 3428 4326 3440 4378
rect 3492 4326 3504 4378
rect 3556 4326 5576 4378
rect 5628 4326 5640 4378
rect 5692 4326 5704 4378
rect 5756 4326 5768 4378
rect 5820 4326 6754 4378
rect 38 4304 6754 4326
rect 52 4020 58 4072
rect 110 4060 116 4072
rect 1619 4063 1677 4069
rect 1619 4060 1631 4063
rect 110 4032 1631 4060
rect 110 4020 116 4032
rect 1619 4029 1631 4032
rect 1665 4029 1677 4063
rect 1619 4023 1677 4029
rect 1886 3995 1944 4001
rect 1886 3961 1898 3995
rect 1932 3992 1944 3995
rect 2076 3992 2082 4004
rect 1932 3964 2082 3992
rect 1932 3961 1944 3964
rect 1886 3955 1944 3961
rect 2076 3952 2082 3964
rect 2134 3952 2140 4004
rect 2999 3927 3057 3933
rect 2999 3893 3011 3927
rect 3045 3924 3057 3927
rect 3640 3924 3646 3936
rect 3045 3896 3646 3924
rect 3045 3893 3057 3896
rect 2999 3887 3057 3893
rect 3640 3884 3646 3896
rect 3698 3924 3704 3936
rect 4744 3924 4750 3936
rect 3698 3896 4750 3924
rect 3698 3884 3704 3896
rect 4744 3884 4750 3896
rect 4802 3884 4808 3936
rect 38 3834 6754 3856
rect 38 3782 2180 3834
rect 2232 3782 2244 3834
rect 2296 3782 2308 3834
rect 2360 3782 2372 3834
rect 2424 3782 4444 3834
rect 4496 3782 4508 3834
rect 4560 3782 4572 3834
rect 4624 3782 4636 3834
rect 4688 3782 6754 3834
rect 38 3760 6754 3782
rect 38 3290 6754 3312
rect 38 3238 1048 3290
rect 1100 3238 1112 3290
rect 1164 3238 1176 3290
rect 1228 3238 1240 3290
rect 1292 3238 3312 3290
rect 3364 3238 3376 3290
rect 3428 3238 3440 3290
rect 3492 3238 3504 3290
rect 3556 3238 5576 3290
rect 5628 3238 5640 3290
rect 5692 3238 5704 3290
rect 5756 3238 5768 3290
rect 5820 3238 6754 3290
rect 38 3216 6754 3238
rect 38 2746 6754 2768
rect 38 2694 2180 2746
rect 2232 2694 2244 2746
rect 2296 2694 2308 2746
rect 2360 2694 2372 2746
rect 2424 2694 4444 2746
rect 4496 2694 4508 2746
rect 4560 2694 4572 2746
rect 4624 2694 4636 2746
rect 4688 2694 6754 2746
rect 38 2672 6754 2694
rect 38 2202 6754 2224
rect 38 2150 1048 2202
rect 1100 2150 1112 2202
rect 1164 2150 1176 2202
rect 1228 2150 1240 2202
rect 1292 2150 3312 2202
rect 3364 2150 3376 2202
rect 3428 2150 3440 2202
rect 3492 2150 3504 2202
rect 3556 2150 5576 2202
rect 5628 2150 5640 2202
rect 5692 2150 5704 2202
rect 5756 2150 5768 2202
rect 5820 2150 6754 2202
rect 38 2128 6754 2150
<< via1 >>
rect 2180 14662 2232 14714
rect 2244 14662 2296 14714
rect 2308 14662 2360 14714
rect 2372 14662 2424 14714
rect 4444 14662 4496 14714
rect 4508 14662 4560 14714
rect 4572 14662 4624 14714
rect 4636 14662 4688 14714
rect 1048 14118 1100 14170
rect 1112 14118 1164 14170
rect 1176 14118 1228 14170
rect 1240 14118 1292 14170
rect 3312 14118 3364 14170
rect 3376 14118 3428 14170
rect 3440 14118 3492 14170
rect 3504 14118 3556 14170
rect 5576 14118 5628 14170
rect 5640 14118 5692 14170
rect 5704 14118 5756 14170
rect 5768 14118 5820 14170
rect 2180 13574 2232 13626
rect 2244 13574 2296 13626
rect 2308 13574 2360 13626
rect 2372 13574 2424 13626
rect 4444 13574 4496 13626
rect 4508 13574 4560 13626
rect 4572 13574 4624 13626
rect 4636 13574 4688 13626
rect 1048 13030 1100 13082
rect 1112 13030 1164 13082
rect 1176 13030 1228 13082
rect 1240 13030 1292 13082
rect 3312 13030 3364 13082
rect 3376 13030 3428 13082
rect 3440 13030 3492 13082
rect 3504 13030 3556 13082
rect 5576 13030 5628 13082
rect 5640 13030 5692 13082
rect 5704 13030 5756 13082
rect 5768 13030 5820 13082
rect 1346 12588 1398 12640
rect 3186 12588 3238 12640
rect 2180 12486 2232 12538
rect 2244 12486 2296 12538
rect 2308 12486 2360 12538
rect 2372 12486 2424 12538
rect 4444 12486 4496 12538
rect 4508 12486 4560 12538
rect 4572 12486 4624 12538
rect 4636 12486 4688 12538
rect 1048 11942 1100 11994
rect 1112 11942 1164 11994
rect 1176 11942 1228 11994
rect 1240 11942 1292 11994
rect 3312 11942 3364 11994
rect 3376 11942 3428 11994
rect 3440 11942 3492 11994
rect 3504 11942 3556 11994
rect 5576 11942 5628 11994
rect 5640 11942 5692 11994
rect 5704 11942 5756 11994
rect 5768 11942 5820 11994
rect 2180 11398 2232 11450
rect 2244 11398 2296 11450
rect 2308 11398 2360 11450
rect 2372 11398 2424 11450
rect 4444 11398 4496 11450
rect 4508 11398 4560 11450
rect 4572 11398 4624 11450
rect 4636 11398 4688 11450
rect 1048 10854 1100 10906
rect 1112 10854 1164 10906
rect 1176 10854 1228 10906
rect 1240 10854 1292 10906
rect 3312 10854 3364 10906
rect 3376 10854 3428 10906
rect 3440 10854 3492 10906
rect 3504 10854 3556 10906
rect 5576 10854 5628 10906
rect 5640 10854 5692 10906
rect 5704 10854 5756 10906
rect 5768 10854 5820 10906
rect 2180 10310 2232 10362
rect 2244 10310 2296 10362
rect 2308 10310 2360 10362
rect 2372 10310 2424 10362
rect 4444 10310 4496 10362
rect 4508 10310 4560 10362
rect 4572 10310 4624 10362
rect 4636 10310 4688 10362
rect 1048 9766 1100 9818
rect 1112 9766 1164 9818
rect 1176 9766 1228 9818
rect 1240 9766 1292 9818
rect 3312 9766 3364 9818
rect 3376 9766 3428 9818
rect 3440 9766 3492 9818
rect 3504 9766 3556 9818
rect 5576 9766 5628 9818
rect 5640 9766 5692 9818
rect 5704 9766 5756 9818
rect 5768 9766 5820 9818
rect 2180 9222 2232 9274
rect 2244 9222 2296 9274
rect 2308 9222 2360 9274
rect 2372 9222 2424 9274
rect 4444 9222 4496 9274
rect 4508 9222 4560 9274
rect 4572 9222 4624 9274
rect 4636 9222 4688 9274
rect 5394 9120 5446 9172
rect 5394 9027 5446 9036
rect 5394 8993 5403 9027
rect 5403 8993 5437 9027
rect 5437 8993 5446 9027
rect 5394 8984 5446 8993
rect 1048 8678 1100 8730
rect 1112 8678 1164 8730
rect 1176 8678 1228 8730
rect 1240 8678 1292 8730
rect 3312 8678 3364 8730
rect 3376 8678 3428 8730
rect 3440 8678 3492 8730
rect 3504 8678 3556 8730
rect 5576 8678 5628 8730
rect 5640 8678 5692 8730
rect 5704 8678 5756 8730
rect 5768 8678 5820 8730
rect 2180 8134 2232 8186
rect 2244 8134 2296 8186
rect 2308 8134 2360 8186
rect 2372 8134 2424 8186
rect 4444 8134 4496 8186
rect 4508 8134 4560 8186
rect 4572 8134 4624 8186
rect 4636 8134 4688 8186
rect 4290 7964 4342 8016
rect 4750 7828 4802 7880
rect 5302 7871 5354 7880
rect 5302 7837 5311 7871
rect 5311 7837 5345 7871
rect 5345 7837 5354 7871
rect 5302 7828 5354 7837
rect 1048 7590 1100 7642
rect 1112 7590 1164 7642
rect 1176 7590 1228 7642
rect 1240 7590 1292 7642
rect 3312 7590 3364 7642
rect 3376 7590 3428 7642
rect 3440 7590 3492 7642
rect 3504 7590 3556 7642
rect 5576 7590 5628 7642
rect 5640 7590 5692 7642
rect 5704 7590 5756 7642
rect 5768 7590 5820 7642
rect 2180 7046 2232 7098
rect 2244 7046 2296 7098
rect 2308 7046 2360 7098
rect 2372 7046 2424 7098
rect 4444 7046 4496 7098
rect 4508 7046 4560 7098
rect 4572 7046 4624 7098
rect 4636 7046 4688 7098
rect 1048 6502 1100 6554
rect 1112 6502 1164 6554
rect 1176 6502 1228 6554
rect 1240 6502 1292 6554
rect 3312 6502 3364 6554
rect 3376 6502 3428 6554
rect 3440 6502 3492 6554
rect 3504 6502 3556 6554
rect 5576 6502 5628 6554
rect 5640 6502 5692 6554
rect 5704 6502 5756 6554
rect 5768 6502 5820 6554
rect 3186 6375 3238 6384
rect 3186 6341 3195 6375
rect 3195 6341 3229 6375
rect 3229 6341 3238 6375
rect 3186 6332 3238 6341
rect 3646 6196 3698 6248
rect 3922 6171 3974 6180
rect 3922 6137 3931 6171
rect 3931 6137 3965 6171
rect 3965 6137 3974 6171
rect 3922 6128 3974 6137
rect 4290 6128 4342 6180
rect 2180 5958 2232 6010
rect 2244 5958 2296 6010
rect 2308 5958 2360 6010
rect 2372 5958 2424 6010
rect 4444 5958 4496 6010
rect 4508 5958 4560 6010
rect 4572 5958 4624 6010
rect 4636 5958 4688 6010
rect 3922 5720 3974 5772
rect 4750 5516 4802 5568
rect 1048 5414 1100 5466
rect 1112 5414 1164 5466
rect 1176 5414 1228 5466
rect 1240 5414 1292 5466
rect 3312 5414 3364 5466
rect 3376 5414 3428 5466
rect 3440 5414 3492 5466
rect 3504 5414 3556 5466
rect 5576 5414 5628 5466
rect 5640 5414 5692 5466
rect 5704 5414 5756 5466
rect 5768 5414 5820 5466
rect 2180 4870 2232 4922
rect 2244 4870 2296 4922
rect 2308 4870 2360 4922
rect 2372 4870 2424 4922
rect 4444 4870 4496 4922
rect 4508 4870 4560 4922
rect 4572 4870 4624 4922
rect 4636 4870 4688 4922
rect 4750 4743 4802 4752
rect 4750 4709 4759 4743
rect 4759 4709 4793 4743
rect 4793 4709 4802 4743
rect 4750 4700 4802 4709
rect 5210 4607 5262 4616
rect 5210 4573 5219 4607
rect 5219 4573 5253 4607
rect 5253 4573 5262 4607
rect 5210 4564 5262 4573
rect 6774 4496 6826 4548
rect 1048 4326 1100 4378
rect 1112 4326 1164 4378
rect 1176 4326 1228 4378
rect 1240 4326 1292 4378
rect 3312 4326 3364 4378
rect 3376 4326 3428 4378
rect 3440 4326 3492 4378
rect 3504 4326 3556 4378
rect 5576 4326 5628 4378
rect 5640 4326 5692 4378
rect 5704 4326 5756 4378
rect 5768 4326 5820 4378
rect 58 4020 110 4072
rect 2082 3952 2134 4004
rect 3646 3884 3698 3936
rect 4750 3884 4802 3936
rect 2180 3782 2232 3834
rect 2244 3782 2296 3834
rect 2308 3782 2360 3834
rect 2372 3782 2424 3834
rect 4444 3782 4496 3834
rect 4508 3782 4560 3834
rect 4572 3782 4624 3834
rect 4636 3782 4688 3834
rect 1048 3238 1100 3290
rect 1112 3238 1164 3290
rect 1176 3238 1228 3290
rect 1240 3238 1292 3290
rect 3312 3238 3364 3290
rect 3376 3238 3428 3290
rect 3440 3238 3492 3290
rect 3504 3238 3556 3290
rect 5576 3238 5628 3290
rect 5640 3238 5692 3290
rect 5704 3238 5756 3290
rect 5768 3238 5820 3290
rect 2180 2694 2232 2746
rect 2244 2694 2296 2746
rect 2308 2694 2360 2746
rect 2372 2694 2424 2746
rect 4444 2694 4496 2746
rect 4508 2694 4560 2746
rect 4572 2694 4624 2746
rect 4636 2694 4688 2746
rect 1048 2150 1100 2202
rect 1112 2150 1164 2202
rect 1176 2150 1228 2202
rect 1240 2150 1292 2202
rect 3312 2150 3364 2202
rect 3376 2150 3428 2202
rect 3440 2150 3492 2202
rect 3504 2150 3556 2202
rect 5576 2150 5628 2202
rect 5640 2150 5692 2202
rect 5704 2150 5756 2202
rect 5768 2150 5820 2202
<< metal2 >>
rect 1160 16520 1216 17000
rect 5668 16520 5724 17000
rect 1174 14362 1202 16520
rect 2154 14716 2450 14736
rect 2210 14714 2234 14716
rect 2290 14714 2314 14716
rect 2370 14714 2394 14716
rect 2232 14662 2234 14714
rect 2296 14662 2308 14714
rect 2370 14662 2372 14714
rect 2210 14660 2234 14662
rect 2290 14660 2314 14662
rect 2370 14660 2394 14662
rect 2154 14640 2450 14660
rect 4418 14716 4714 14736
rect 4474 14714 4498 14716
rect 4554 14714 4578 14716
rect 4634 14714 4658 14716
rect 4496 14662 4498 14714
rect 4560 14662 4572 14714
rect 4634 14662 4636 14714
rect 4474 14660 4498 14662
rect 4554 14660 4578 14662
rect 4634 14660 4658 14662
rect 4418 14640 4714 14660
rect 4288 14376 4344 14385
rect 1174 14334 1386 14362
rect 1022 14172 1318 14192
rect 1078 14170 1102 14172
rect 1158 14170 1182 14172
rect 1238 14170 1262 14172
rect 1100 14118 1102 14170
rect 1164 14118 1176 14170
rect 1238 14118 1240 14170
rect 1078 14116 1102 14118
rect 1158 14116 1182 14118
rect 1238 14116 1262 14118
rect 1022 14096 1318 14116
rect 1022 13084 1318 13104
rect 1078 13082 1102 13084
rect 1158 13082 1182 13084
rect 1238 13082 1262 13084
rect 1100 13030 1102 13082
rect 1164 13030 1176 13082
rect 1238 13030 1240 13082
rect 1078 13028 1102 13030
rect 1158 13028 1182 13030
rect 1238 13028 1262 13030
rect 1022 13008 1318 13028
rect 1358 12646 1386 14334
rect 5682 14362 5710 16520
rect 4288 14311 4344 14320
rect 5314 14334 5710 14362
rect 3286 14172 3582 14192
rect 3342 14170 3366 14172
rect 3422 14170 3446 14172
rect 3502 14170 3526 14172
rect 3364 14118 3366 14170
rect 3428 14118 3440 14170
rect 3502 14118 3504 14170
rect 3342 14116 3366 14118
rect 3422 14116 3446 14118
rect 3502 14116 3526 14118
rect 3286 14096 3582 14116
rect 2154 13628 2450 13648
rect 2210 13626 2234 13628
rect 2290 13626 2314 13628
rect 2370 13626 2394 13628
rect 2232 13574 2234 13626
rect 2296 13574 2308 13626
rect 2370 13574 2372 13626
rect 2210 13572 2234 13574
rect 2290 13572 2314 13574
rect 2370 13572 2394 13574
rect 2154 13552 2450 13572
rect 3286 13084 3582 13104
rect 3342 13082 3366 13084
rect 3422 13082 3446 13084
rect 3502 13082 3526 13084
rect 3364 13030 3366 13082
rect 3428 13030 3440 13082
rect 3502 13030 3504 13082
rect 3342 13028 3366 13030
rect 3422 13028 3446 13030
rect 3502 13028 3526 13030
rect 3286 13008 3582 13028
rect 1346 12640 1398 12646
rect 1346 12582 1398 12588
rect 3186 12640 3238 12646
rect 3186 12582 3238 12588
rect 2154 12540 2450 12560
rect 2210 12538 2234 12540
rect 2290 12538 2314 12540
rect 2370 12538 2394 12540
rect 2232 12486 2234 12538
rect 2296 12486 2308 12538
rect 2370 12486 2372 12538
rect 2210 12484 2234 12486
rect 2290 12484 2314 12486
rect 2370 12484 2394 12486
rect 2154 12464 2450 12484
rect 1022 11996 1318 12016
rect 1078 11994 1102 11996
rect 1158 11994 1182 11996
rect 1238 11994 1262 11996
rect 1100 11942 1102 11994
rect 1164 11942 1176 11994
rect 1238 11942 1240 11994
rect 1078 11940 1102 11942
rect 1158 11940 1182 11942
rect 1238 11940 1262 11942
rect 1022 11920 1318 11940
rect 2154 11452 2450 11472
rect 2210 11450 2234 11452
rect 2290 11450 2314 11452
rect 2370 11450 2394 11452
rect 2232 11398 2234 11450
rect 2296 11398 2308 11450
rect 2370 11398 2372 11450
rect 2210 11396 2234 11398
rect 2290 11396 2314 11398
rect 2370 11396 2394 11398
rect 2154 11376 2450 11396
rect 1022 10908 1318 10928
rect 1078 10906 1102 10908
rect 1158 10906 1182 10908
rect 1238 10906 1262 10908
rect 1100 10854 1102 10906
rect 1164 10854 1176 10906
rect 1238 10854 1240 10906
rect 1078 10852 1102 10854
rect 1158 10852 1182 10854
rect 1238 10852 1262 10854
rect 1022 10832 1318 10852
rect 2154 10364 2450 10384
rect 2210 10362 2234 10364
rect 2290 10362 2314 10364
rect 2370 10362 2394 10364
rect 2232 10310 2234 10362
rect 2296 10310 2308 10362
rect 2370 10310 2372 10362
rect 2210 10308 2234 10310
rect 2290 10308 2314 10310
rect 2370 10308 2394 10310
rect 2154 10288 2450 10308
rect 1022 9820 1318 9840
rect 1078 9818 1102 9820
rect 1158 9818 1182 9820
rect 1238 9818 1262 9820
rect 1100 9766 1102 9818
rect 1164 9766 1176 9818
rect 1238 9766 1240 9818
rect 1078 9764 1102 9766
rect 1158 9764 1182 9766
rect 1238 9764 1262 9766
rect 1022 9744 1318 9764
rect 2154 9276 2450 9296
rect 2210 9274 2234 9276
rect 2290 9274 2314 9276
rect 2370 9274 2394 9276
rect 2232 9222 2234 9274
rect 2296 9222 2308 9274
rect 2370 9222 2372 9274
rect 2210 9220 2234 9222
rect 2290 9220 2314 9222
rect 2370 9220 2394 9222
rect 2154 9200 2450 9220
rect 1022 8732 1318 8752
rect 1078 8730 1102 8732
rect 1158 8730 1182 8732
rect 1238 8730 1262 8732
rect 1100 8678 1102 8730
rect 1164 8678 1176 8730
rect 1238 8678 1240 8730
rect 1078 8676 1102 8678
rect 1158 8676 1182 8678
rect 1238 8676 1262 8678
rect 1022 8656 1318 8676
rect 2154 8188 2450 8208
rect 2210 8186 2234 8188
rect 2290 8186 2314 8188
rect 2370 8186 2394 8188
rect 2232 8134 2234 8186
rect 2296 8134 2308 8186
rect 2370 8134 2372 8186
rect 2210 8132 2234 8134
rect 2290 8132 2314 8134
rect 2370 8132 2394 8134
rect 2154 8112 2450 8132
rect 1022 7644 1318 7664
rect 1078 7642 1102 7644
rect 1158 7642 1182 7644
rect 1238 7642 1262 7644
rect 1100 7590 1102 7642
rect 1164 7590 1176 7642
rect 1238 7590 1240 7642
rect 1078 7588 1102 7590
rect 1158 7588 1182 7590
rect 1238 7588 1262 7590
rect 1022 7568 1318 7588
rect 2154 7100 2450 7120
rect 2210 7098 2234 7100
rect 2290 7098 2314 7100
rect 2370 7098 2394 7100
rect 2232 7046 2234 7098
rect 2296 7046 2308 7098
rect 2370 7046 2372 7098
rect 2210 7044 2234 7046
rect 2290 7044 2314 7046
rect 2370 7044 2394 7046
rect 2154 7024 2450 7044
rect 1022 6556 1318 6576
rect 1078 6554 1102 6556
rect 1158 6554 1182 6556
rect 1238 6554 1262 6556
rect 1100 6502 1102 6554
rect 1164 6502 1176 6554
rect 1238 6502 1240 6554
rect 1078 6500 1102 6502
rect 1158 6500 1182 6502
rect 1238 6500 1262 6502
rect 1022 6480 1318 6500
rect 3198 6390 3226 12582
rect 3286 11996 3582 12016
rect 3342 11994 3366 11996
rect 3422 11994 3446 11996
rect 3502 11994 3526 11996
rect 3364 11942 3366 11994
rect 3428 11942 3440 11994
rect 3502 11942 3504 11994
rect 3342 11940 3366 11942
rect 3422 11940 3446 11942
rect 3502 11940 3526 11942
rect 3286 11920 3582 11940
rect 3286 10908 3582 10928
rect 3342 10906 3366 10908
rect 3422 10906 3446 10908
rect 3502 10906 3526 10908
rect 3364 10854 3366 10906
rect 3428 10854 3440 10906
rect 3502 10854 3504 10906
rect 3342 10852 3366 10854
rect 3422 10852 3446 10854
rect 3502 10852 3526 10854
rect 3286 10832 3582 10852
rect 3286 9820 3582 9840
rect 3342 9818 3366 9820
rect 3422 9818 3446 9820
rect 3502 9818 3526 9820
rect 3364 9766 3366 9818
rect 3428 9766 3440 9818
rect 3502 9766 3504 9818
rect 3342 9764 3366 9766
rect 3422 9764 3446 9766
rect 3502 9764 3526 9766
rect 3286 9744 3582 9764
rect 3286 8732 3582 8752
rect 3342 8730 3366 8732
rect 3422 8730 3446 8732
rect 3502 8730 3526 8732
rect 3364 8678 3366 8730
rect 3428 8678 3440 8730
rect 3502 8678 3504 8730
rect 3342 8676 3366 8678
rect 3422 8676 3446 8678
rect 3502 8676 3526 8678
rect 3286 8656 3582 8676
rect 4302 8022 4330 14311
rect 4418 13628 4714 13648
rect 4474 13626 4498 13628
rect 4554 13626 4578 13628
rect 4634 13626 4658 13628
rect 4496 13574 4498 13626
rect 4560 13574 4572 13626
rect 4634 13574 4636 13626
rect 4474 13572 4498 13574
rect 4554 13572 4578 13574
rect 4634 13572 4658 13574
rect 4418 13552 4714 13572
rect 4418 12540 4714 12560
rect 4474 12538 4498 12540
rect 4554 12538 4578 12540
rect 4634 12538 4658 12540
rect 4496 12486 4498 12538
rect 4560 12486 4572 12538
rect 4634 12486 4636 12538
rect 4474 12484 4498 12486
rect 4554 12484 4578 12486
rect 4634 12484 4658 12486
rect 4418 12464 4714 12484
rect 4418 11452 4714 11472
rect 4474 11450 4498 11452
rect 4554 11450 4578 11452
rect 4634 11450 4658 11452
rect 4496 11398 4498 11450
rect 4560 11398 4572 11450
rect 4634 11398 4636 11450
rect 4474 11396 4498 11398
rect 4554 11396 4578 11398
rect 4634 11396 4658 11398
rect 4418 11376 4714 11396
rect 4418 10364 4714 10384
rect 4474 10362 4498 10364
rect 4554 10362 4578 10364
rect 4634 10362 4658 10364
rect 4496 10310 4498 10362
rect 4560 10310 4572 10362
rect 4634 10310 4636 10362
rect 4474 10308 4498 10310
rect 4554 10308 4578 10310
rect 4634 10308 4658 10310
rect 4418 10288 4714 10308
rect 4418 9276 4714 9296
rect 4474 9274 4498 9276
rect 4554 9274 4578 9276
rect 4634 9274 4658 9276
rect 4496 9222 4498 9274
rect 4560 9222 4572 9274
rect 4634 9222 4636 9274
rect 4474 9220 4498 9222
rect 4554 9220 4578 9222
rect 4634 9220 4658 9222
rect 4418 9200 4714 9220
rect 4418 8188 4714 8208
rect 4474 8186 4498 8188
rect 4554 8186 4578 8188
rect 4634 8186 4658 8188
rect 4496 8134 4498 8186
rect 4560 8134 4572 8186
rect 4634 8134 4636 8186
rect 4474 8132 4498 8134
rect 4554 8132 4578 8134
rect 4634 8132 4658 8134
rect 4418 8112 4714 8132
rect 4290 8016 4342 8022
rect 4290 7958 4342 7964
rect 3286 7644 3582 7664
rect 3342 7642 3366 7644
rect 3422 7642 3446 7644
rect 3502 7642 3526 7644
rect 3364 7590 3366 7642
rect 3428 7590 3440 7642
rect 3502 7590 3504 7642
rect 3342 7588 3366 7590
rect 3422 7588 3446 7590
rect 3502 7588 3526 7590
rect 3286 7568 3582 7588
rect 3286 6556 3582 6576
rect 3342 6554 3366 6556
rect 3422 6554 3446 6556
rect 3502 6554 3526 6556
rect 3364 6502 3366 6554
rect 3428 6502 3440 6554
rect 3502 6502 3504 6554
rect 3342 6500 3366 6502
rect 3422 6500 3446 6502
rect 3502 6500 3526 6502
rect 3286 6480 3582 6500
rect 3186 6384 3238 6390
rect 3186 6326 3238 6332
rect 3646 6248 3698 6254
rect 3646 6190 3698 6196
rect 2154 6012 2450 6032
rect 2210 6010 2234 6012
rect 2290 6010 2314 6012
rect 2370 6010 2394 6012
rect 2232 5958 2234 6010
rect 2296 5958 2308 6010
rect 2370 5958 2372 6010
rect 2210 5956 2234 5958
rect 2290 5956 2314 5958
rect 2370 5956 2394 5958
rect 2154 5936 2450 5956
rect 1022 5468 1318 5488
rect 1078 5466 1102 5468
rect 1158 5466 1182 5468
rect 1238 5466 1262 5468
rect 1100 5414 1102 5466
rect 1164 5414 1176 5466
rect 1238 5414 1240 5466
rect 1078 5412 1102 5414
rect 1158 5412 1182 5414
rect 1238 5412 1262 5414
rect 1022 5392 1318 5412
rect 3286 5468 3582 5488
rect 3342 5466 3366 5468
rect 3422 5466 3446 5468
rect 3502 5466 3526 5468
rect 3364 5414 3366 5466
rect 3428 5414 3440 5466
rect 3502 5414 3504 5466
rect 3342 5412 3366 5414
rect 3422 5412 3446 5414
rect 3502 5412 3526 5414
rect 3286 5392 3582 5412
rect 2154 4924 2450 4944
rect 2210 4922 2234 4924
rect 2290 4922 2314 4924
rect 2370 4922 2394 4924
rect 2232 4870 2234 4922
rect 2296 4870 2308 4922
rect 2370 4870 2372 4922
rect 2210 4868 2234 4870
rect 2290 4868 2314 4870
rect 2370 4868 2394 4870
rect 2154 4848 2450 4868
rect 1022 4380 1318 4400
rect 1078 4378 1102 4380
rect 1158 4378 1182 4380
rect 1238 4378 1262 4380
rect 1100 4326 1102 4378
rect 1164 4326 1176 4378
rect 1238 4326 1240 4378
rect 1078 4324 1102 4326
rect 1158 4324 1182 4326
rect 1238 4324 1262 4326
rect 1022 4304 1318 4324
rect 3286 4380 3582 4400
rect 3342 4378 3366 4380
rect 3422 4378 3446 4380
rect 3502 4378 3526 4380
rect 3364 4326 3366 4378
rect 3428 4326 3440 4378
rect 3502 4326 3504 4378
rect 3342 4324 3366 4326
rect 3422 4324 3446 4326
rect 3502 4324 3526 4326
rect 3286 4304 3582 4324
rect 58 4072 110 4078
rect 58 4014 110 4020
rect 70 480 98 4014
rect 2082 4004 2134 4010
rect 2082 3946 2134 3952
rect 1022 3292 1318 3312
rect 1078 3290 1102 3292
rect 1158 3290 1182 3292
rect 1238 3290 1262 3292
rect 1100 3238 1102 3290
rect 1164 3238 1176 3290
rect 1238 3238 1240 3290
rect 1078 3236 1102 3238
rect 1158 3236 1182 3238
rect 1238 3236 1262 3238
rect 1022 3216 1318 3236
rect 1022 2204 1318 2224
rect 1078 2202 1102 2204
rect 1158 2202 1182 2204
rect 1238 2202 1262 2204
rect 1100 2150 1102 2202
rect 1164 2150 1176 2202
rect 1238 2150 1240 2202
rect 1078 2148 1102 2150
rect 1158 2148 1182 2150
rect 1238 2148 1262 2150
rect 1022 2128 1318 2148
rect 2094 1986 2122 3946
rect 3658 3942 3686 6190
rect 4302 6186 4330 7958
rect 5314 7886 5342 14334
rect 5550 14172 5846 14192
rect 5606 14170 5630 14172
rect 5686 14170 5710 14172
rect 5766 14170 5790 14172
rect 5628 14118 5630 14170
rect 5692 14118 5704 14170
rect 5766 14118 5768 14170
rect 5606 14116 5630 14118
rect 5686 14116 5710 14118
rect 5766 14116 5790 14118
rect 5550 14096 5846 14116
rect 5550 13084 5846 13104
rect 5606 13082 5630 13084
rect 5686 13082 5710 13084
rect 5766 13082 5790 13084
rect 5628 13030 5630 13082
rect 5692 13030 5704 13082
rect 5766 13030 5768 13082
rect 5606 13028 5630 13030
rect 5686 13028 5710 13030
rect 5766 13028 5790 13030
rect 5550 13008 5846 13028
rect 5550 11996 5846 12016
rect 5606 11994 5630 11996
rect 5686 11994 5710 11996
rect 5766 11994 5790 11996
rect 5628 11942 5630 11994
rect 5692 11942 5704 11994
rect 5766 11942 5768 11994
rect 5606 11940 5630 11942
rect 5686 11940 5710 11942
rect 5766 11940 5790 11942
rect 5550 11920 5846 11940
rect 5550 10908 5846 10928
rect 5606 10906 5630 10908
rect 5686 10906 5710 10908
rect 5766 10906 5790 10908
rect 5628 10854 5630 10906
rect 5692 10854 5704 10906
rect 5766 10854 5768 10906
rect 5606 10852 5630 10854
rect 5686 10852 5710 10854
rect 5766 10852 5790 10854
rect 5550 10832 5846 10852
rect 5392 10568 5448 10577
rect 5392 10503 5448 10512
rect 5406 9178 5434 10503
rect 5550 9820 5846 9840
rect 5606 9818 5630 9820
rect 5686 9818 5710 9820
rect 5766 9818 5790 9820
rect 5628 9766 5630 9818
rect 5692 9766 5704 9818
rect 5766 9766 5768 9818
rect 5606 9764 5630 9766
rect 5686 9764 5710 9766
rect 5766 9764 5790 9766
rect 5550 9744 5846 9764
rect 5394 9172 5446 9178
rect 5394 9114 5446 9120
rect 5394 9036 5446 9042
rect 5394 8978 5446 8984
rect 4750 7880 4802 7886
rect 4750 7822 4802 7828
rect 5302 7880 5354 7886
rect 5302 7822 5354 7828
rect 4418 7100 4714 7120
rect 4474 7098 4498 7100
rect 4554 7098 4578 7100
rect 4634 7098 4658 7100
rect 4496 7046 4498 7098
rect 4560 7046 4572 7098
rect 4634 7046 4636 7098
rect 4474 7044 4498 7046
rect 4554 7044 4578 7046
rect 4634 7044 4658 7046
rect 4418 7024 4714 7044
rect 4762 6361 4790 7822
rect 4748 6352 4804 6361
rect 4748 6287 4804 6296
rect 3922 6180 3974 6186
rect 3922 6122 3974 6128
rect 4290 6180 4342 6186
rect 4290 6122 4342 6128
rect 3934 5778 3962 6122
rect 4418 6012 4714 6032
rect 4474 6010 4498 6012
rect 4554 6010 4578 6012
rect 4634 6010 4658 6012
rect 4496 5958 4498 6010
rect 4560 5958 4572 6010
rect 4634 5958 4636 6010
rect 4474 5956 4498 5958
rect 4554 5956 4578 5958
rect 4634 5956 4658 5958
rect 4418 5936 4714 5956
rect 3922 5772 3974 5778
rect 3922 5714 3974 5720
rect 4750 5568 4802 5574
rect 4750 5510 4802 5516
rect 4418 4924 4714 4944
rect 4474 4922 4498 4924
rect 4554 4922 4578 4924
rect 4634 4922 4658 4924
rect 4496 4870 4498 4922
rect 4560 4870 4572 4922
rect 4634 4870 4636 4922
rect 4474 4868 4498 4870
rect 4554 4868 4578 4870
rect 4634 4868 4658 4870
rect 4418 4848 4714 4868
rect 4762 4758 4790 5510
rect 4750 4752 4802 4758
rect 5406 4706 5434 8978
rect 5550 8732 5846 8752
rect 5606 8730 5630 8732
rect 5686 8730 5710 8732
rect 5766 8730 5790 8732
rect 5628 8678 5630 8730
rect 5692 8678 5704 8730
rect 5766 8678 5768 8730
rect 5606 8676 5630 8678
rect 5686 8676 5710 8678
rect 5766 8676 5790 8678
rect 5550 8656 5846 8676
rect 5550 7644 5846 7664
rect 5606 7642 5630 7644
rect 5686 7642 5710 7644
rect 5766 7642 5790 7644
rect 5628 7590 5630 7642
rect 5692 7590 5704 7642
rect 5766 7590 5768 7642
rect 5606 7588 5630 7590
rect 5686 7588 5710 7590
rect 5766 7588 5790 7590
rect 5550 7568 5846 7588
rect 5550 6556 5846 6576
rect 5606 6554 5630 6556
rect 5686 6554 5710 6556
rect 5766 6554 5790 6556
rect 5628 6502 5630 6554
rect 5692 6502 5704 6554
rect 5766 6502 5768 6554
rect 5606 6500 5630 6502
rect 5686 6500 5710 6502
rect 5766 6500 5790 6502
rect 5550 6480 5846 6500
rect 5550 5468 5846 5488
rect 5606 5466 5630 5468
rect 5686 5466 5710 5468
rect 5766 5466 5790 5468
rect 5628 5414 5630 5466
rect 5692 5414 5704 5466
rect 5766 5414 5768 5466
rect 5606 5412 5630 5414
rect 5686 5412 5710 5414
rect 5766 5412 5790 5414
rect 5550 5392 5846 5412
rect 4750 4694 4802 4700
rect 5222 4678 5434 4706
rect 5222 4622 5250 4678
rect 5210 4616 5262 4622
rect 5210 4558 5262 4564
rect 3646 3936 3698 3942
rect 3646 3878 3698 3884
rect 4750 3936 4802 3942
rect 4750 3878 4802 3884
rect 2154 3836 2450 3856
rect 2210 3834 2234 3836
rect 2290 3834 2314 3836
rect 2370 3834 2394 3836
rect 2232 3782 2234 3834
rect 2296 3782 2308 3834
rect 2370 3782 2372 3834
rect 2210 3780 2234 3782
rect 2290 3780 2314 3782
rect 2370 3780 2394 3782
rect 2154 3760 2450 3780
rect 4418 3836 4714 3856
rect 4474 3834 4498 3836
rect 4554 3834 4578 3836
rect 4634 3834 4658 3836
rect 4496 3782 4498 3834
rect 4560 3782 4572 3834
rect 4634 3782 4636 3834
rect 4474 3780 4498 3782
rect 4554 3780 4578 3782
rect 4634 3780 4658 3782
rect 4418 3760 4714 3780
rect 3286 3292 3582 3312
rect 3342 3290 3366 3292
rect 3422 3290 3446 3292
rect 3502 3290 3526 3292
rect 3364 3238 3366 3290
rect 3428 3238 3440 3290
rect 3502 3238 3504 3290
rect 3342 3236 3366 3238
rect 3422 3236 3446 3238
rect 3502 3236 3526 3238
rect 3286 3216 3582 3236
rect 2154 2748 2450 2768
rect 2210 2746 2234 2748
rect 2290 2746 2314 2748
rect 2370 2746 2394 2748
rect 2232 2694 2234 2746
rect 2296 2694 2308 2746
rect 2370 2694 2372 2746
rect 2210 2692 2234 2694
rect 2290 2692 2314 2694
rect 2370 2692 2394 2694
rect 2154 2672 2450 2692
rect 4418 2748 4714 2768
rect 4474 2746 4498 2748
rect 4554 2746 4578 2748
rect 4634 2746 4658 2748
rect 4496 2694 4498 2746
rect 4560 2694 4572 2746
rect 4634 2694 4636 2746
rect 4474 2692 4498 2694
rect 4554 2692 4578 2694
rect 4634 2692 4658 2694
rect 4418 2672 4714 2692
rect 4762 2530 4790 3878
rect 4578 2502 4790 2530
rect 3286 2204 3582 2224
rect 3342 2202 3366 2204
rect 3422 2202 3446 2204
rect 3502 2202 3526 2204
rect 3364 2150 3366 2202
rect 3428 2150 3440 2202
rect 3502 2150 3504 2202
rect 3342 2148 3366 2150
rect 3422 2148 3446 2150
rect 3502 2148 3526 2150
rect 3286 2128 3582 2148
rect 2094 1958 2306 1986
rect 2278 480 2306 1958
rect 4578 480 4606 2502
rect 5222 2417 5250 4558
rect 6774 4548 6826 4554
rect 6774 4490 6826 4496
rect 5550 4380 5846 4400
rect 5606 4378 5630 4380
rect 5686 4378 5710 4380
rect 5766 4378 5790 4380
rect 5628 4326 5630 4378
rect 5692 4326 5704 4378
rect 5766 4326 5768 4378
rect 5606 4324 5630 4326
rect 5686 4324 5710 4326
rect 5766 4324 5790 4326
rect 5550 4304 5846 4324
rect 5550 3292 5846 3312
rect 5606 3290 5630 3292
rect 5686 3290 5710 3292
rect 5766 3290 5790 3292
rect 5628 3238 5630 3290
rect 5692 3238 5704 3290
rect 5766 3238 5768 3290
rect 5606 3236 5630 3238
rect 5686 3236 5710 3238
rect 5766 3236 5790 3238
rect 5550 3216 5846 3236
rect 5208 2408 5264 2417
rect 5208 2343 5264 2352
rect 5550 2204 5846 2224
rect 5606 2202 5630 2204
rect 5686 2202 5710 2204
rect 5766 2202 5790 2204
rect 5628 2150 5630 2202
rect 5692 2150 5704 2202
rect 5766 2150 5768 2202
rect 5606 2148 5630 2150
rect 5686 2148 5710 2150
rect 5766 2148 5790 2150
rect 5550 2128 5846 2148
rect 6786 480 6814 4490
rect 56 0 112 480
rect 2264 0 2320 480
rect 4564 0 4620 480
rect 6772 0 6828 480
<< via2 >>
rect 2154 14714 2210 14716
rect 2234 14714 2290 14716
rect 2314 14714 2370 14716
rect 2394 14714 2450 14716
rect 2154 14662 2180 14714
rect 2180 14662 2210 14714
rect 2234 14662 2244 14714
rect 2244 14662 2290 14714
rect 2314 14662 2360 14714
rect 2360 14662 2370 14714
rect 2394 14662 2424 14714
rect 2424 14662 2450 14714
rect 2154 14660 2210 14662
rect 2234 14660 2290 14662
rect 2314 14660 2370 14662
rect 2394 14660 2450 14662
rect 4418 14714 4474 14716
rect 4498 14714 4554 14716
rect 4578 14714 4634 14716
rect 4658 14714 4714 14716
rect 4418 14662 4444 14714
rect 4444 14662 4474 14714
rect 4498 14662 4508 14714
rect 4508 14662 4554 14714
rect 4578 14662 4624 14714
rect 4624 14662 4634 14714
rect 4658 14662 4688 14714
rect 4688 14662 4714 14714
rect 4418 14660 4474 14662
rect 4498 14660 4554 14662
rect 4578 14660 4634 14662
rect 4658 14660 4714 14662
rect 1022 14170 1078 14172
rect 1102 14170 1158 14172
rect 1182 14170 1238 14172
rect 1262 14170 1318 14172
rect 1022 14118 1048 14170
rect 1048 14118 1078 14170
rect 1102 14118 1112 14170
rect 1112 14118 1158 14170
rect 1182 14118 1228 14170
rect 1228 14118 1238 14170
rect 1262 14118 1292 14170
rect 1292 14118 1318 14170
rect 1022 14116 1078 14118
rect 1102 14116 1158 14118
rect 1182 14116 1238 14118
rect 1262 14116 1318 14118
rect 1022 13082 1078 13084
rect 1102 13082 1158 13084
rect 1182 13082 1238 13084
rect 1262 13082 1318 13084
rect 1022 13030 1048 13082
rect 1048 13030 1078 13082
rect 1102 13030 1112 13082
rect 1112 13030 1158 13082
rect 1182 13030 1228 13082
rect 1228 13030 1238 13082
rect 1262 13030 1292 13082
rect 1292 13030 1318 13082
rect 1022 13028 1078 13030
rect 1102 13028 1158 13030
rect 1182 13028 1238 13030
rect 1262 13028 1318 13030
rect 4288 14320 4344 14376
rect 3286 14170 3342 14172
rect 3366 14170 3422 14172
rect 3446 14170 3502 14172
rect 3526 14170 3582 14172
rect 3286 14118 3312 14170
rect 3312 14118 3342 14170
rect 3366 14118 3376 14170
rect 3376 14118 3422 14170
rect 3446 14118 3492 14170
rect 3492 14118 3502 14170
rect 3526 14118 3556 14170
rect 3556 14118 3582 14170
rect 3286 14116 3342 14118
rect 3366 14116 3422 14118
rect 3446 14116 3502 14118
rect 3526 14116 3582 14118
rect 2154 13626 2210 13628
rect 2234 13626 2290 13628
rect 2314 13626 2370 13628
rect 2394 13626 2450 13628
rect 2154 13574 2180 13626
rect 2180 13574 2210 13626
rect 2234 13574 2244 13626
rect 2244 13574 2290 13626
rect 2314 13574 2360 13626
rect 2360 13574 2370 13626
rect 2394 13574 2424 13626
rect 2424 13574 2450 13626
rect 2154 13572 2210 13574
rect 2234 13572 2290 13574
rect 2314 13572 2370 13574
rect 2394 13572 2450 13574
rect 3286 13082 3342 13084
rect 3366 13082 3422 13084
rect 3446 13082 3502 13084
rect 3526 13082 3582 13084
rect 3286 13030 3312 13082
rect 3312 13030 3342 13082
rect 3366 13030 3376 13082
rect 3376 13030 3422 13082
rect 3446 13030 3492 13082
rect 3492 13030 3502 13082
rect 3526 13030 3556 13082
rect 3556 13030 3582 13082
rect 3286 13028 3342 13030
rect 3366 13028 3422 13030
rect 3446 13028 3502 13030
rect 3526 13028 3582 13030
rect 2154 12538 2210 12540
rect 2234 12538 2290 12540
rect 2314 12538 2370 12540
rect 2394 12538 2450 12540
rect 2154 12486 2180 12538
rect 2180 12486 2210 12538
rect 2234 12486 2244 12538
rect 2244 12486 2290 12538
rect 2314 12486 2360 12538
rect 2360 12486 2370 12538
rect 2394 12486 2424 12538
rect 2424 12486 2450 12538
rect 2154 12484 2210 12486
rect 2234 12484 2290 12486
rect 2314 12484 2370 12486
rect 2394 12484 2450 12486
rect 1022 11994 1078 11996
rect 1102 11994 1158 11996
rect 1182 11994 1238 11996
rect 1262 11994 1318 11996
rect 1022 11942 1048 11994
rect 1048 11942 1078 11994
rect 1102 11942 1112 11994
rect 1112 11942 1158 11994
rect 1182 11942 1228 11994
rect 1228 11942 1238 11994
rect 1262 11942 1292 11994
rect 1292 11942 1318 11994
rect 1022 11940 1078 11942
rect 1102 11940 1158 11942
rect 1182 11940 1238 11942
rect 1262 11940 1318 11942
rect 2154 11450 2210 11452
rect 2234 11450 2290 11452
rect 2314 11450 2370 11452
rect 2394 11450 2450 11452
rect 2154 11398 2180 11450
rect 2180 11398 2210 11450
rect 2234 11398 2244 11450
rect 2244 11398 2290 11450
rect 2314 11398 2360 11450
rect 2360 11398 2370 11450
rect 2394 11398 2424 11450
rect 2424 11398 2450 11450
rect 2154 11396 2210 11398
rect 2234 11396 2290 11398
rect 2314 11396 2370 11398
rect 2394 11396 2450 11398
rect 1022 10906 1078 10908
rect 1102 10906 1158 10908
rect 1182 10906 1238 10908
rect 1262 10906 1318 10908
rect 1022 10854 1048 10906
rect 1048 10854 1078 10906
rect 1102 10854 1112 10906
rect 1112 10854 1158 10906
rect 1182 10854 1228 10906
rect 1228 10854 1238 10906
rect 1262 10854 1292 10906
rect 1292 10854 1318 10906
rect 1022 10852 1078 10854
rect 1102 10852 1158 10854
rect 1182 10852 1238 10854
rect 1262 10852 1318 10854
rect 2154 10362 2210 10364
rect 2234 10362 2290 10364
rect 2314 10362 2370 10364
rect 2394 10362 2450 10364
rect 2154 10310 2180 10362
rect 2180 10310 2210 10362
rect 2234 10310 2244 10362
rect 2244 10310 2290 10362
rect 2314 10310 2360 10362
rect 2360 10310 2370 10362
rect 2394 10310 2424 10362
rect 2424 10310 2450 10362
rect 2154 10308 2210 10310
rect 2234 10308 2290 10310
rect 2314 10308 2370 10310
rect 2394 10308 2450 10310
rect 1022 9818 1078 9820
rect 1102 9818 1158 9820
rect 1182 9818 1238 9820
rect 1262 9818 1318 9820
rect 1022 9766 1048 9818
rect 1048 9766 1078 9818
rect 1102 9766 1112 9818
rect 1112 9766 1158 9818
rect 1182 9766 1228 9818
rect 1228 9766 1238 9818
rect 1262 9766 1292 9818
rect 1292 9766 1318 9818
rect 1022 9764 1078 9766
rect 1102 9764 1158 9766
rect 1182 9764 1238 9766
rect 1262 9764 1318 9766
rect 2154 9274 2210 9276
rect 2234 9274 2290 9276
rect 2314 9274 2370 9276
rect 2394 9274 2450 9276
rect 2154 9222 2180 9274
rect 2180 9222 2210 9274
rect 2234 9222 2244 9274
rect 2244 9222 2290 9274
rect 2314 9222 2360 9274
rect 2360 9222 2370 9274
rect 2394 9222 2424 9274
rect 2424 9222 2450 9274
rect 2154 9220 2210 9222
rect 2234 9220 2290 9222
rect 2314 9220 2370 9222
rect 2394 9220 2450 9222
rect 1022 8730 1078 8732
rect 1102 8730 1158 8732
rect 1182 8730 1238 8732
rect 1262 8730 1318 8732
rect 1022 8678 1048 8730
rect 1048 8678 1078 8730
rect 1102 8678 1112 8730
rect 1112 8678 1158 8730
rect 1182 8678 1228 8730
rect 1228 8678 1238 8730
rect 1262 8678 1292 8730
rect 1292 8678 1318 8730
rect 1022 8676 1078 8678
rect 1102 8676 1158 8678
rect 1182 8676 1238 8678
rect 1262 8676 1318 8678
rect 2154 8186 2210 8188
rect 2234 8186 2290 8188
rect 2314 8186 2370 8188
rect 2394 8186 2450 8188
rect 2154 8134 2180 8186
rect 2180 8134 2210 8186
rect 2234 8134 2244 8186
rect 2244 8134 2290 8186
rect 2314 8134 2360 8186
rect 2360 8134 2370 8186
rect 2394 8134 2424 8186
rect 2424 8134 2450 8186
rect 2154 8132 2210 8134
rect 2234 8132 2290 8134
rect 2314 8132 2370 8134
rect 2394 8132 2450 8134
rect 1022 7642 1078 7644
rect 1102 7642 1158 7644
rect 1182 7642 1238 7644
rect 1262 7642 1318 7644
rect 1022 7590 1048 7642
rect 1048 7590 1078 7642
rect 1102 7590 1112 7642
rect 1112 7590 1158 7642
rect 1182 7590 1228 7642
rect 1228 7590 1238 7642
rect 1262 7590 1292 7642
rect 1292 7590 1318 7642
rect 1022 7588 1078 7590
rect 1102 7588 1158 7590
rect 1182 7588 1238 7590
rect 1262 7588 1318 7590
rect 2154 7098 2210 7100
rect 2234 7098 2290 7100
rect 2314 7098 2370 7100
rect 2394 7098 2450 7100
rect 2154 7046 2180 7098
rect 2180 7046 2210 7098
rect 2234 7046 2244 7098
rect 2244 7046 2290 7098
rect 2314 7046 2360 7098
rect 2360 7046 2370 7098
rect 2394 7046 2424 7098
rect 2424 7046 2450 7098
rect 2154 7044 2210 7046
rect 2234 7044 2290 7046
rect 2314 7044 2370 7046
rect 2394 7044 2450 7046
rect 1022 6554 1078 6556
rect 1102 6554 1158 6556
rect 1182 6554 1238 6556
rect 1262 6554 1318 6556
rect 1022 6502 1048 6554
rect 1048 6502 1078 6554
rect 1102 6502 1112 6554
rect 1112 6502 1158 6554
rect 1182 6502 1228 6554
rect 1228 6502 1238 6554
rect 1262 6502 1292 6554
rect 1292 6502 1318 6554
rect 1022 6500 1078 6502
rect 1102 6500 1158 6502
rect 1182 6500 1238 6502
rect 1262 6500 1318 6502
rect 3286 11994 3342 11996
rect 3366 11994 3422 11996
rect 3446 11994 3502 11996
rect 3526 11994 3582 11996
rect 3286 11942 3312 11994
rect 3312 11942 3342 11994
rect 3366 11942 3376 11994
rect 3376 11942 3422 11994
rect 3446 11942 3492 11994
rect 3492 11942 3502 11994
rect 3526 11942 3556 11994
rect 3556 11942 3582 11994
rect 3286 11940 3342 11942
rect 3366 11940 3422 11942
rect 3446 11940 3502 11942
rect 3526 11940 3582 11942
rect 3286 10906 3342 10908
rect 3366 10906 3422 10908
rect 3446 10906 3502 10908
rect 3526 10906 3582 10908
rect 3286 10854 3312 10906
rect 3312 10854 3342 10906
rect 3366 10854 3376 10906
rect 3376 10854 3422 10906
rect 3446 10854 3492 10906
rect 3492 10854 3502 10906
rect 3526 10854 3556 10906
rect 3556 10854 3582 10906
rect 3286 10852 3342 10854
rect 3366 10852 3422 10854
rect 3446 10852 3502 10854
rect 3526 10852 3582 10854
rect 3286 9818 3342 9820
rect 3366 9818 3422 9820
rect 3446 9818 3502 9820
rect 3526 9818 3582 9820
rect 3286 9766 3312 9818
rect 3312 9766 3342 9818
rect 3366 9766 3376 9818
rect 3376 9766 3422 9818
rect 3446 9766 3492 9818
rect 3492 9766 3502 9818
rect 3526 9766 3556 9818
rect 3556 9766 3582 9818
rect 3286 9764 3342 9766
rect 3366 9764 3422 9766
rect 3446 9764 3502 9766
rect 3526 9764 3582 9766
rect 3286 8730 3342 8732
rect 3366 8730 3422 8732
rect 3446 8730 3502 8732
rect 3526 8730 3582 8732
rect 3286 8678 3312 8730
rect 3312 8678 3342 8730
rect 3366 8678 3376 8730
rect 3376 8678 3422 8730
rect 3446 8678 3492 8730
rect 3492 8678 3502 8730
rect 3526 8678 3556 8730
rect 3556 8678 3582 8730
rect 3286 8676 3342 8678
rect 3366 8676 3422 8678
rect 3446 8676 3502 8678
rect 3526 8676 3582 8678
rect 4418 13626 4474 13628
rect 4498 13626 4554 13628
rect 4578 13626 4634 13628
rect 4658 13626 4714 13628
rect 4418 13574 4444 13626
rect 4444 13574 4474 13626
rect 4498 13574 4508 13626
rect 4508 13574 4554 13626
rect 4578 13574 4624 13626
rect 4624 13574 4634 13626
rect 4658 13574 4688 13626
rect 4688 13574 4714 13626
rect 4418 13572 4474 13574
rect 4498 13572 4554 13574
rect 4578 13572 4634 13574
rect 4658 13572 4714 13574
rect 4418 12538 4474 12540
rect 4498 12538 4554 12540
rect 4578 12538 4634 12540
rect 4658 12538 4714 12540
rect 4418 12486 4444 12538
rect 4444 12486 4474 12538
rect 4498 12486 4508 12538
rect 4508 12486 4554 12538
rect 4578 12486 4624 12538
rect 4624 12486 4634 12538
rect 4658 12486 4688 12538
rect 4688 12486 4714 12538
rect 4418 12484 4474 12486
rect 4498 12484 4554 12486
rect 4578 12484 4634 12486
rect 4658 12484 4714 12486
rect 4418 11450 4474 11452
rect 4498 11450 4554 11452
rect 4578 11450 4634 11452
rect 4658 11450 4714 11452
rect 4418 11398 4444 11450
rect 4444 11398 4474 11450
rect 4498 11398 4508 11450
rect 4508 11398 4554 11450
rect 4578 11398 4624 11450
rect 4624 11398 4634 11450
rect 4658 11398 4688 11450
rect 4688 11398 4714 11450
rect 4418 11396 4474 11398
rect 4498 11396 4554 11398
rect 4578 11396 4634 11398
rect 4658 11396 4714 11398
rect 4418 10362 4474 10364
rect 4498 10362 4554 10364
rect 4578 10362 4634 10364
rect 4658 10362 4714 10364
rect 4418 10310 4444 10362
rect 4444 10310 4474 10362
rect 4498 10310 4508 10362
rect 4508 10310 4554 10362
rect 4578 10310 4624 10362
rect 4624 10310 4634 10362
rect 4658 10310 4688 10362
rect 4688 10310 4714 10362
rect 4418 10308 4474 10310
rect 4498 10308 4554 10310
rect 4578 10308 4634 10310
rect 4658 10308 4714 10310
rect 4418 9274 4474 9276
rect 4498 9274 4554 9276
rect 4578 9274 4634 9276
rect 4658 9274 4714 9276
rect 4418 9222 4444 9274
rect 4444 9222 4474 9274
rect 4498 9222 4508 9274
rect 4508 9222 4554 9274
rect 4578 9222 4624 9274
rect 4624 9222 4634 9274
rect 4658 9222 4688 9274
rect 4688 9222 4714 9274
rect 4418 9220 4474 9222
rect 4498 9220 4554 9222
rect 4578 9220 4634 9222
rect 4658 9220 4714 9222
rect 4418 8186 4474 8188
rect 4498 8186 4554 8188
rect 4578 8186 4634 8188
rect 4658 8186 4714 8188
rect 4418 8134 4444 8186
rect 4444 8134 4474 8186
rect 4498 8134 4508 8186
rect 4508 8134 4554 8186
rect 4578 8134 4624 8186
rect 4624 8134 4634 8186
rect 4658 8134 4688 8186
rect 4688 8134 4714 8186
rect 4418 8132 4474 8134
rect 4498 8132 4554 8134
rect 4578 8132 4634 8134
rect 4658 8132 4714 8134
rect 3286 7642 3342 7644
rect 3366 7642 3422 7644
rect 3446 7642 3502 7644
rect 3526 7642 3582 7644
rect 3286 7590 3312 7642
rect 3312 7590 3342 7642
rect 3366 7590 3376 7642
rect 3376 7590 3422 7642
rect 3446 7590 3492 7642
rect 3492 7590 3502 7642
rect 3526 7590 3556 7642
rect 3556 7590 3582 7642
rect 3286 7588 3342 7590
rect 3366 7588 3422 7590
rect 3446 7588 3502 7590
rect 3526 7588 3582 7590
rect 3286 6554 3342 6556
rect 3366 6554 3422 6556
rect 3446 6554 3502 6556
rect 3526 6554 3582 6556
rect 3286 6502 3312 6554
rect 3312 6502 3342 6554
rect 3366 6502 3376 6554
rect 3376 6502 3422 6554
rect 3446 6502 3492 6554
rect 3492 6502 3502 6554
rect 3526 6502 3556 6554
rect 3556 6502 3582 6554
rect 3286 6500 3342 6502
rect 3366 6500 3422 6502
rect 3446 6500 3502 6502
rect 3526 6500 3582 6502
rect 2154 6010 2210 6012
rect 2234 6010 2290 6012
rect 2314 6010 2370 6012
rect 2394 6010 2450 6012
rect 2154 5958 2180 6010
rect 2180 5958 2210 6010
rect 2234 5958 2244 6010
rect 2244 5958 2290 6010
rect 2314 5958 2360 6010
rect 2360 5958 2370 6010
rect 2394 5958 2424 6010
rect 2424 5958 2450 6010
rect 2154 5956 2210 5958
rect 2234 5956 2290 5958
rect 2314 5956 2370 5958
rect 2394 5956 2450 5958
rect 1022 5466 1078 5468
rect 1102 5466 1158 5468
rect 1182 5466 1238 5468
rect 1262 5466 1318 5468
rect 1022 5414 1048 5466
rect 1048 5414 1078 5466
rect 1102 5414 1112 5466
rect 1112 5414 1158 5466
rect 1182 5414 1228 5466
rect 1228 5414 1238 5466
rect 1262 5414 1292 5466
rect 1292 5414 1318 5466
rect 1022 5412 1078 5414
rect 1102 5412 1158 5414
rect 1182 5412 1238 5414
rect 1262 5412 1318 5414
rect 3286 5466 3342 5468
rect 3366 5466 3422 5468
rect 3446 5466 3502 5468
rect 3526 5466 3582 5468
rect 3286 5414 3312 5466
rect 3312 5414 3342 5466
rect 3366 5414 3376 5466
rect 3376 5414 3422 5466
rect 3446 5414 3492 5466
rect 3492 5414 3502 5466
rect 3526 5414 3556 5466
rect 3556 5414 3582 5466
rect 3286 5412 3342 5414
rect 3366 5412 3422 5414
rect 3446 5412 3502 5414
rect 3526 5412 3582 5414
rect 2154 4922 2210 4924
rect 2234 4922 2290 4924
rect 2314 4922 2370 4924
rect 2394 4922 2450 4924
rect 2154 4870 2180 4922
rect 2180 4870 2210 4922
rect 2234 4870 2244 4922
rect 2244 4870 2290 4922
rect 2314 4870 2360 4922
rect 2360 4870 2370 4922
rect 2394 4870 2424 4922
rect 2424 4870 2450 4922
rect 2154 4868 2210 4870
rect 2234 4868 2290 4870
rect 2314 4868 2370 4870
rect 2394 4868 2450 4870
rect 1022 4378 1078 4380
rect 1102 4378 1158 4380
rect 1182 4378 1238 4380
rect 1262 4378 1318 4380
rect 1022 4326 1048 4378
rect 1048 4326 1078 4378
rect 1102 4326 1112 4378
rect 1112 4326 1158 4378
rect 1182 4326 1228 4378
rect 1228 4326 1238 4378
rect 1262 4326 1292 4378
rect 1292 4326 1318 4378
rect 1022 4324 1078 4326
rect 1102 4324 1158 4326
rect 1182 4324 1238 4326
rect 1262 4324 1318 4326
rect 3286 4378 3342 4380
rect 3366 4378 3422 4380
rect 3446 4378 3502 4380
rect 3526 4378 3582 4380
rect 3286 4326 3312 4378
rect 3312 4326 3342 4378
rect 3366 4326 3376 4378
rect 3376 4326 3422 4378
rect 3446 4326 3492 4378
rect 3492 4326 3502 4378
rect 3526 4326 3556 4378
rect 3556 4326 3582 4378
rect 3286 4324 3342 4326
rect 3366 4324 3422 4326
rect 3446 4324 3502 4326
rect 3526 4324 3582 4326
rect 1022 3290 1078 3292
rect 1102 3290 1158 3292
rect 1182 3290 1238 3292
rect 1262 3290 1318 3292
rect 1022 3238 1048 3290
rect 1048 3238 1078 3290
rect 1102 3238 1112 3290
rect 1112 3238 1158 3290
rect 1182 3238 1228 3290
rect 1228 3238 1238 3290
rect 1262 3238 1292 3290
rect 1292 3238 1318 3290
rect 1022 3236 1078 3238
rect 1102 3236 1158 3238
rect 1182 3236 1238 3238
rect 1262 3236 1318 3238
rect 1022 2202 1078 2204
rect 1102 2202 1158 2204
rect 1182 2202 1238 2204
rect 1262 2202 1318 2204
rect 1022 2150 1048 2202
rect 1048 2150 1078 2202
rect 1102 2150 1112 2202
rect 1112 2150 1158 2202
rect 1182 2150 1228 2202
rect 1228 2150 1238 2202
rect 1262 2150 1292 2202
rect 1292 2150 1318 2202
rect 1022 2148 1078 2150
rect 1102 2148 1158 2150
rect 1182 2148 1238 2150
rect 1262 2148 1318 2150
rect 5550 14170 5606 14172
rect 5630 14170 5686 14172
rect 5710 14170 5766 14172
rect 5790 14170 5846 14172
rect 5550 14118 5576 14170
rect 5576 14118 5606 14170
rect 5630 14118 5640 14170
rect 5640 14118 5686 14170
rect 5710 14118 5756 14170
rect 5756 14118 5766 14170
rect 5790 14118 5820 14170
rect 5820 14118 5846 14170
rect 5550 14116 5606 14118
rect 5630 14116 5686 14118
rect 5710 14116 5766 14118
rect 5790 14116 5846 14118
rect 5550 13082 5606 13084
rect 5630 13082 5686 13084
rect 5710 13082 5766 13084
rect 5790 13082 5846 13084
rect 5550 13030 5576 13082
rect 5576 13030 5606 13082
rect 5630 13030 5640 13082
rect 5640 13030 5686 13082
rect 5710 13030 5756 13082
rect 5756 13030 5766 13082
rect 5790 13030 5820 13082
rect 5820 13030 5846 13082
rect 5550 13028 5606 13030
rect 5630 13028 5686 13030
rect 5710 13028 5766 13030
rect 5790 13028 5846 13030
rect 5550 11994 5606 11996
rect 5630 11994 5686 11996
rect 5710 11994 5766 11996
rect 5790 11994 5846 11996
rect 5550 11942 5576 11994
rect 5576 11942 5606 11994
rect 5630 11942 5640 11994
rect 5640 11942 5686 11994
rect 5710 11942 5756 11994
rect 5756 11942 5766 11994
rect 5790 11942 5820 11994
rect 5820 11942 5846 11994
rect 5550 11940 5606 11942
rect 5630 11940 5686 11942
rect 5710 11940 5766 11942
rect 5790 11940 5846 11942
rect 5550 10906 5606 10908
rect 5630 10906 5686 10908
rect 5710 10906 5766 10908
rect 5790 10906 5846 10908
rect 5550 10854 5576 10906
rect 5576 10854 5606 10906
rect 5630 10854 5640 10906
rect 5640 10854 5686 10906
rect 5710 10854 5756 10906
rect 5756 10854 5766 10906
rect 5790 10854 5820 10906
rect 5820 10854 5846 10906
rect 5550 10852 5606 10854
rect 5630 10852 5686 10854
rect 5710 10852 5766 10854
rect 5790 10852 5846 10854
rect 5392 10512 5448 10568
rect 5550 9818 5606 9820
rect 5630 9818 5686 9820
rect 5710 9818 5766 9820
rect 5790 9818 5846 9820
rect 5550 9766 5576 9818
rect 5576 9766 5606 9818
rect 5630 9766 5640 9818
rect 5640 9766 5686 9818
rect 5710 9766 5756 9818
rect 5756 9766 5766 9818
rect 5790 9766 5820 9818
rect 5820 9766 5846 9818
rect 5550 9764 5606 9766
rect 5630 9764 5686 9766
rect 5710 9764 5766 9766
rect 5790 9764 5846 9766
rect 4418 7098 4474 7100
rect 4498 7098 4554 7100
rect 4578 7098 4634 7100
rect 4658 7098 4714 7100
rect 4418 7046 4444 7098
rect 4444 7046 4474 7098
rect 4498 7046 4508 7098
rect 4508 7046 4554 7098
rect 4578 7046 4624 7098
rect 4624 7046 4634 7098
rect 4658 7046 4688 7098
rect 4688 7046 4714 7098
rect 4418 7044 4474 7046
rect 4498 7044 4554 7046
rect 4578 7044 4634 7046
rect 4658 7044 4714 7046
rect 4748 6296 4804 6352
rect 4418 6010 4474 6012
rect 4498 6010 4554 6012
rect 4578 6010 4634 6012
rect 4658 6010 4714 6012
rect 4418 5958 4444 6010
rect 4444 5958 4474 6010
rect 4498 5958 4508 6010
rect 4508 5958 4554 6010
rect 4578 5958 4624 6010
rect 4624 5958 4634 6010
rect 4658 5958 4688 6010
rect 4688 5958 4714 6010
rect 4418 5956 4474 5958
rect 4498 5956 4554 5958
rect 4578 5956 4634 5958
rect 4658 5956 4714 5958
rect 4418 4922 4474 4924
rect 4498 4922 4554 4924
rect 4578 4922 4634 4924
rect 4658 4922 4714 4924
rect 4418 4870 4444 4922
rect 4444 4870 4474 4922
rect 4498 4870 4508 4922
rect 4508 4870 4554 4922
rect 4578 4870 4624 4922
rect 4624 4870 4634 4922
rect 4658 4870 4688 4922
rect 4688 4870 4714 4922
rect 4418 4868 4474 4870
rect 4498 4868 4554 4870
rect 4578 4868 4634 4870
rect 4658 4868 4714 4870
rect 5550 8730 5606 8732
rect 5630 8730 5686 8732
rect 5710 8730 5766 8732
rect 5790 8730 5846 8732
rect 5550 8678 5576 8730
rect 5576 8678 5606 8730
rect 5630 8678 5640 8730
rect 5640 8678 5686 8730
rect 5710 8678 5756 8730
rect 5756 8678 5766 8730
rect 5790 8678 5820 8730
rect 5820 8678 5846 8730
rect 5550 8676 5606 8678
rect 5630 8676 5686 8678
rect 5710 8676 5766 8678
rect 5790 8676 5846 8678
rect 5550 7642 5606 7644
rect 5630 7642 5686 7644
rect 5710 7642 5766 7644
rect 5790 7642 5846 7644
rect 5550 7590 5576 7642
rect 5576 7590 5606 7642
rect 5630 7590 5640 7642
rect 5640 7590 5686 7642
rect 5710 7590 5756 7642
rect 5756 7590 5766 7642
rect 5790 7590 5820 7642
rect 5820 7590 5846 7642
rect 5550 7588 5606 7590
rect 5630 7588 5686 7590
rect 5710 7588 5766 7590
rect 5790 7588 5846 7590
rect 5550 6554 5606 6556
rect 5630 6554 5686 6556
rect 5710 6554 5766 6556
rect 5790 6554 5846 6556
rect 5550 6502 5576 6554
rect 5576 6502 5606 6554
rect 5630 6502 5640 6554
rect 5640 6502 5686 6554
rect 5710 6502 5756 6554
rect 5756 6502 5766 6554
rect 5790 6502 5820 6554
rect 5820 6502 5846 6554
rect 5550 6500 5606 6502
rect 5630 6500 5686 6502
rect 5710 6500 5766 6502
rect 5790 6500 5846 6502
rect 5550 5466 5606 5468
rect 5630 5466 5686 5468
rect 5710 5466 5766 5468
rect 5790 5466 5846 5468
rect 5550 5414 5576 5466
rect 5576 5414 5606 5466
rect 5630 5414 5640 5466
rect 5640 5414 5686 5466
rect 5710 5414 5756 5466
rect 5756 5414 5766 5466
rect 5790 5414 5820 5466
rect 5820 5414 5846 5466
rect 5550 5412 5606 5414
rect 5630 5412 5686 5414
rect 5710 5412 5766 5414
rect 5790 5412 5846 5414
rect 2154 3834 2210 3836
rect 2234 3834 2290 3836
rect 2314 3834 2370 3836
rect 2394 3834 2450 3836
rect 2154 3782 2180 3834
rect 2180 3782 2210 3834
rect 2234 3782 2244 3834
rect 2244 3782 2290 3834
rect 2314 3782 2360 3834
rect 2360 3782 2370 3834
rect 2394 3782 2424 3834
rect 2424 3782 2450 3834
rect 2154 3780 2210 3782
rect 2234 3780 2290 3782
rect 2314 3780 2370 3782
rect 2394 3780 2450 3782
rect 4418 3834 4474 3836
rect 4498 3834 4554 3836
rect 4578 3834 4634 3836
rect 4658 3834 4714 3836
rect 4418 3782 4444 3834
rect 4444 3782 4474 3834
rect 4498 3782 4508 3834
rect 4508 3782 4554 3834
rect 4578 3782 4624 3834
rect 4624 3782 4634 3834
rect 4658 3782 4688 3834
rect 4688 3782 4714 3834
rect 4418 3780 4474 3782
rect 4498 3780 4554 3782
rect 4578 3780 4634 3782
rect 4658 3780 4714 3782
rect 3286 3290 3342 3292
rect 3366 3290 3422 3292
rect 3446 3290 3502 3292
rect 3526 3290 3582 3292
rect 3286 3238 3312 3290
rect 3312 3238 3342 3290
rect 3366 3238 3376 3290
rect 3376 3238 3422 3290
rect 3446 3238 3492 3290
rect 3492 3238 3502 3290
rect 3526 3238 3556 3290
rect 3556 3238 3582 3290
rect 3286 3236 3342 3238
rect 3366 3236 3422 3238
rect 3446 3236 3502 3238
rect 3526 3236 3582 3238
rect 2154 2746 2210 2748
rect 2234 2746 2290 2748
rect 2314 2746 2370 2748
rect 2394 2746 2450 2748
rect 2154 2694 2180 2746
rect 2180 2694 2210 2746
rect 2234 2694 2244 2746
rect 2244 2694 2290 2746
rect 2314 2694 2360 2746
rect 2360 2694 2370 2746
rect 2394 2694 2424 2746
rect 2424 2694 2450 2746
rect 2154 2692 2210 2694
rect 2234 2692 2290 2694
rect 2314 2692 2370 2694
rect 2394 2692 2450 2694
rect 4418 2746 4474 2748
rect 4498 2746 4554 2748
rect 4578 2746 4634 2748
rect 4658 2746 4714 2748
rect 4418 2694 4444 2746
rect 4444 2694 4474 2746
rect 4498 2694 4508 2746
rect 4508 2694 4554 2746
rect 4578 2694 4624 2746
rect 4624 2694 4634 2746
rect 4658 2694 4688 2746
rect 4688 2694 4714 2746
rect 4418 2692 4474 2694
rect 4498 2692 4554 2694
rect 4578 2692 4634 2694
rect 4658 2692 4714 2694
rect 3286 2202 3342 2204
rect 3366 2202 3422 2204
rect 3446 2202 3502 2204
rect 3526 2202 3582 2204
rect 3286 2150 3312 2202
rect 3312 2150 3342 2202
rect 3366 2150 3376 2202
rect 3376 2150 3422 2202
rect 3446 2150 3492 2202
rect 3492 2150 3502 2202
rect 3526 2150 3556 2202
rect 3556 2150 3582 2202
rect 3286 2148 3342 2150
rect 3366 2148 3422 2150
rect 3446 2148 3502 2150
rect 3526 2148 3582 2150
rect 5550 4378 5606 4380
rect 5630 4378 5686 4380
rect 5710 4378 5766 4380
rect 5790 4378 5846 4380
rect 5550 4326 5576 4378
rect 5576 4326 5606 4378
rect 5630 4326 5640 4378
rect 5640 4326 5686 4378
rect 5710 4326 5756 4378
rect 5756 4326 5766 4378
rect 5790 4326 5820 4378
rect 5820 4326 5846 4378
rect 5550 4324 5606 4326
rect 5630 4324 5686 4326
rect 5710 4324 5766 4326
rect 5790 4324 5846 4326
rect 5550 3290 5606 3292
rect 5630 3290 5686 3292
rect 5710 3290 5766 3292
rect 5790 3290 5846 3292
rect 5550 3238 5576 3290
rect 5576 3238 5606 3290
rect 5630 3238 5640 3290
rect 5640 3238 5686 3290
rect 5710 3238 5756 3290
rect 5756 3238 5766 3290
rect 5790 3238 5820 3290
rect 5820 3238 5846 3290
rect 5550 3236 5606 3238
rect 5630 3236 5686 3238
rect 5710 3236 5766 3238
rect 5790 3236 5846 3238
rect 5208 2352 5264 2408
rect 5550 2202 5606 2204
rect 5630 2202 5686 2204
rect 5710 2202 5766 2204
rect 5790 2202 5846 2204
rect 5550 2150 5576 2202
rect 5576 2150 5606 2202
rect 5630 2150 5640 2202
rect 5640 2150 5686 2202
rect 5710 2150 5756 2202
rect 5756 2150 5766 2202
rect 5790 2150 5820 2202
rect 5820 2150 5846 2202
rect 5550 2148 5606 2150
rect 5630 2148 5686 2150
rect 5710 2148 5766 2150
rect 5790 2148 5846 2150
<< metal3 >>
rect 7454 14786 7934 14816
rect 4884 14726 7934 14786
rect 2142 14720 2462 14721
rect 2142 14656 2150 14720
rect 2214 14656 2230 14720
rect 2294 14656 2310 14720
rect 2374 14656 2390 14720
rect 2454 14656 2462 14720
rect 2142 14655 2462 14656
rect 4406 14720 4726 14721
rect 4406 14656 4414 14720
rect 4478 14656 4494 14720
rect 4558 14656 4574 14720
rect 4638 14656 4654 14720
rect 4718 14656 4726 14720
rect 4406 14655 4726 14656
rect 4283 14378 4349 14381
rect 4884 14378 4944 14726
rect 7454 14696 7934 14726
rect 4283 14376 4944 14378
rect 4283 14320 4288 14376
rect 4344 14320 4944 14376
rect 4283 14318 4944 14320
rect 4283 14315 4349 14318
rect 1010 14176 1330 14177
rect 1010 14112 1018 14176
rect 1082 14112 1098 14176
rect 1162 14112 1178 14176
rect 1242 14112 1258 14176
rect 1322 14112 1330 14176
rect 1010 14111 1330 14112
rect 3274 14176 3594 14177
rect 3274 14112 3282 14176
rect 3346 14112 3362 14176
rect 3426 14112 3442 14176
rect 3506 14112 3522 14176
rect 3586 14112 3594 14176
rect 3274 14111 3594 14112
rect 5538 14176 5858 14177
rect 5538 14112 5546 14176
rect 5610 14112 5626 14176
rect 5690 14112 5706 14176
rect 5770 14112 5786 14176
rect 5850 14112 5858 14176
rect 5538 14111 5858 14112
rect 2142 13632 2462 13633
rect 2142 13568 2150 13632
rect 2214 13568 2230 13632
rect 2294 13568 2310 13632
rect 2374 13568 2390 13632
rect 2454 13568 2462 13632
rect 2142 13567 2462 13568
rect 4406 13632 4726 13633
rect 4406 13568 4414 13632
rect 4478 13568 4494 13632
rect 4558 13568 4574 13632
rect 4638 13568 4654 13632
rect 4718 13568 4726 13632
rect 4406 13567 4726 13568
rect 1010 13088 1330 13089
rect 1010 13024 1018 13088
rect 1082 13024 1098 13088
rect 1162 13024 1178 13088
rect 1242 13024 1258 13088
rect 1322 13024 1330 13088
rect 1010 13023 1330 13024
rect 3274 13088 3594 13089
rect 3274 13024 3282 13088
rect 3346 13024 3362 13088
rect 3426 13024 3442 13088
rect 3506 13024 3522 13088
rect 3586 13024 3594 13088
rect 3274 13023 3594 13024
rect 5538 13088 5858 13089
rect 5538 13024 5546 13088
rect 5610 13024 5626 13088
rect 5690 13024 5706 13088
rect 5770 13024 5786 13088
rect 5850 13024 5858 13088
rect 5538 13023 5858 13024
rect 2142 12544 2462 12545
rect 2142 12480 2150 12544
rect 2214 12480 2230 12544
rect 2294 12480 2310 12544
rect 2374 12480 2390 12544
rect 2454 12480 2462 12544
rect 2142 12479 2462 12480
rect 4406 12544 4726 12545
rect 4406 12480 4414 12544
rect 4478 12480 4494 12544
rect 4558 12480 4574 12544
rect 4638 12480 4654 12544
rect 4718 12480 4726 12544
rect 4406 12479 4726 12480
rect 1010 12000 1330 12001
rect 1010 11936 1018 12000
rect 1082 11936 1098 12000
rect 1162 11936 1178 12000
rect 1242 11936 1258 12000
rect 1322 11936 1330 12000
rect 1010 11935 1330 11936
rect 3274 12000 3594 12001
rect 3274 11936 3282 12000
rect 3346 11936 3362 12000
rect 3426 11936 3442 12000
rect 3506 11936 3522 12000
rect 3586 11936 3594 12000
rect 3274 11935 3594 11936
rect 5538 12000 5858 12001
rect 5538 11936 5546 12000
rect 5610 11936 5626 12000
rect 5690 11936 5706 12000
rect 5770 11936 5786 12000
rect 5850 11936 5858 12000
rect 5538 11935 5858 11936
rect 2142 11456 2462 11457
rect 2142 11392 2150 11456
rect 2214 11392 2230 11456
rect 2294 11392 2310 11456
rect 2374 11392 2390 11456
rect 2454 11392 2462 11456
rect 2142 11391 2462 11392
rect 4406 11456 4726 11457
rect 4406 11392 4414 11456
rect 4478 11392 4494 11456
rect 4558 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4726 11456
rect 4406 11391 4726 11392
rect 1010 10912 1330 10913
rect 1010 10848 1018 10912
rect 1082 10848 1098 10912
rect 1162 10848 1178 10912
rect 1242 10848 1258 10912
rect 1322 10848 1330 10912
rect 1010 10847 1330 10848
rect 3274 10912 3594 10913
rect 3274 10848 3282 10912
rect 3346 10848 3362 10912
rect 3426 10848 3442 10912
rect 3506 10848 3522 10912
rect 3586 10848 3594 10912
rect 3274 10847 3594 10848
rect 5538 10912 5858 10913
rect 5538 10848 5546 10912
rect 5610 10848 5626 10912
rect 5690 10848 5706 10912
rect 5770 10848 5786 10912
rect 5850 10848 5858 10912
rect 5538 10847 5858 10848
rect 5387 10570 5453 10573
rect 7454 10570 7934 10600
rect 5387 10568 7934 10570
rect 5387 10512 5392 10568
rect 5448 10512 7934 10568
rect 5387 10510 7934 10512
rect 5387 10507 5453 10510
rect 7454 10480 7934 10510
rect 2142 10368 2462 10369
rect 2142 10304 2150 10368
rect 2214 10304 2230 10368
rect 2294 10304 2310 10368
rect 2374 10304 2390 10368
rect 2454 10304 2462 10368
rect 2142 10303 2462 10304
rect 4406 10368 4726 10369
rect 4406 10304 4414 10368
rect 4478 10304 4494 10368
rect 4558 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4726 10368
rect 4406 10303 4726 10304
rect 1010 9824 1330 9825
rect 1010 9760 1018 9824
rect 1082 9760 1098 9824
rect 1162 9760 1178 9824
rect 1242 9760 1258 9824
rect 1322 9760 1330 9824
rect 1010 9759 1330 9760
rect 3274 9824 3594 9825
rect 3274 9760 3282 9824
rect 3346 9760 3362 9824
rect 3426 9760 3442 9824
rect 3506 9760 3522 9824
rect 3586 9760 3594 9824
rect 3274 9759 3594 9760
rect 5538 9824 5858 9825
rect 5538 9760 5546 9824
rect 5610 9760 5626 9824
rect 5690 9760 5706 9824
rect 5770 9760 5786 9824
rect 5850 9760 5858 9824
rect 5538 9759 5858 9760
rect 2142 9280 2462 9281
rect 2142 9216 2150 9280
rect 2214 9216 2230 9280
rect 2294 9216 2310 9280
rect 2374 9216 2390 9280
rect 2454 9216 2462 9280
rect 2142 9215 2462 9216
rect 4406 9280 4726 9281
rect 4406 9216 4414 9280
rect 4478 9216 4494 9280
rect 4558 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4726 9280
rect 4406 9215 4726 9216
rect 1010 8736 1330 8737
rect 1010 8672 1018 8736
rect 1082 8672 1098 8736
rect 1162 8672 1178 8736
rect 1242 8672 1258 8736
rect 1322 8672 1330 8736
rect 1010 8671 1330 8672
rect 3274 8736 3594 8737
rect 3274 8672 3282 8736
rect 3346 8672 3362 8736
rect 3426 8672 3442 8736
rect 3506 8672 3522 8736
rect 3586 8672 3594 8736
rect 3274 8671 3594 8672
rect 5538 8736 5858 8737
rect 5538 8672 5546 8736
rect 5610 8672 5626 8736
rect 5690 8672 5706 8736
rect 5770 8672 5786 8736
rect 5850 8672 5858 8736
rect 5538 8671 5858 8672
rect 2142 8192 2462 8193
rect 2142 8128 2150 8192
rect 2214 8128 2230 8192
rect 2294 8128 2310 8192
rect 2374 8128 2390 8192
rect 2454 8128 2462 8192
rect 2142 8127 2462 8128
rect 4406 8192 4726 8193
rect 4406 8128 4414 8192
rect 4478 8128 4494 8192
rect 4558 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4726 8192
rect 4406 8127 4726 8128
rect 1010 7648 1330 7649
rect 1010 7584 1018 7648
rect 1082 7584 1098 7648
rect 1162 7584 1178 7648
rect 1242 7584 1258 7648
rect 1322 7584 1330 7648
rect 1010 7583 1330 7584
rect 3274 7648 3594 7649
rect 3274 7584 3282 7648
rect 3346 7584 3362 7648
rect 3426 7584 3442 7648
rect 3506 7584 3522 7648
rect 3586 7584 3594 7648
rect 3274 7583 3594 7584
rect 5538 7648 5858 7649
rect 5538 7584 5546 7648
rect 5610 7584 5626 7648
rect 5690 7584 5706 7648
rect 5770 7584 5786 7648
rect 5850 7584 5858 7648
rect 5538 7583 5858 7584
rect 2142 7104 2462 7105
rect 2142 7040 2150 7104
rect 2214 7040 2230 7104
rect 2294 7040 2310 7104
rect 2374 7040 2390 7104
rect 2454 7040 2462 7104
rect 2142 7039 2462 7040
rect 4406 7104 4726 7105
rect 4406 7040 4414 7104
rect 4478 7040 4494 7104
rect 4558 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4726 7104
rect 4406 7039 4726 7040
rect 1010 6560 1330 6561
rect 1010 6496 1018 6560
rect 1082 6496 1098 6560
rect 1162 6496 1178 6560
rect 1242 6496 1258 6560
rect 1322 6496 1330 6560
rect 1010 6495 1330 6496
rect 3274 6560 3594 6561
rect 3274 6496 3282 6560
rect 3346 6496 3362 6560
rect 3426 6496 3442 6560
rect 3506 6496 3522 6560
rect 3586 6496 3594 6560
rect 3274 6495 3594 6496
rect 5538 6560 5858 6561
rect 5538 6496 5546 6560
rect 5610 6496 5626 6560
rect 5690 6496 5706 6560
rect 5770 6496 5786 6560
rect 5850 6496 5858 6560
rect 5538 6495 5858 6496
rect 4743 6354 4809 6357
rect 7454 6354 7934 6384
rect 4743 6352 7934 6354
rect 4743 6296 4748 6352
rect 4804 6296 7934 6352
rect 4743 6294 7934 6296
rect 4743 6291 4809 6294
rect 7454 6264 7934 6294
rect 2142 6016 2462 6017
rect 2142 5952 2150 6016
rect 2214 5952 2230 6016
rect 2294 5952 2310 6016
rect 2374 5952 2390 6016
rect 2454 5952 2462 6016
rect 2142 5951 2462 5952
rect 4406 6016 4726 6017
rect 4406 5952 4414 6016
rect 4478 5952 4494 6016
rect 4558 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4726 6016
rect 4406 5951 4726 5952
rect 1010 5472 1330 5473
rect 1010 5408 1018 5472
rect 1082 5408 1098 5472
rect 1162 5408 1178 5472
rect 1242 5408 1258 5472
rect 1322 5408 1330 5472
rect 1010 5407 1330 5408
rect 3274 5472 3594 5473
rect 3274 5408 3282 5472
rect 3346 5408 3362 5472
rect 3426 5408 3442 5472
rect 3506 5408 3522 5472
rect 3586 5408 3594 5472
rect 3274 5407 3594 5408
rect 5538 5472 5858 5473
rect 5538 5408 5546 5472
rect 5610 5408 5626 5472
rect 5690 5408 5706 5472
rect 5770 5408 5786 5472
rect 5850 5408 5858 5472
rect 5538 5407 5858 5408
rect 2142 4928 2462 4929
rect 2142 4864 2150 4928
rect 2214 4864 2230 4928
rect 2294 4864 2310 4928
rect 2374 4864 2390 4928
rect 2454 4864 2462 4928
rect 2142 4863 2462 4864
rect 4406 4928 4726 4929
rect 4406 4864 4414 4928
rect 4478 4864 4494 4928
rect 4558 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4726 4928
rect 4406 4863 4726 4864
rect 1010 4384 1330 4385
rect 1010 4320 1018 4384
rect 1082 4320 1098 4384
rect 1162 4320 1178 4384
rect 1242 4320 1258 4384
rect 1322 4320 1330 4384
rect 1010 4319 1330 4320
rect 3274 4384 3594 4385
rect 3274 4320 3282 4384
rect 3346 4320 3362 4384
rect 3426 4320 3442 4384
rect 3506 4320 3522 4384
rect 3586 4320 3594 4384
rect 3274 4319 3594 4320
rect 5538 4384 5858 4385
rect 5538 4320 5546 4384
rect 5610 4320 5626 4384
rect 5690 4320 5706 4384
rect 5770 4320 5786 4384
rect 5850 4320 5858 4384
rect 5538 4319 5858 4320
rect 2142 3840 2462 3841
rect 2142 3776 2150 3840
rect 2214 3776 2230 3840
rect 2294 3776 2310 3840
rect 2374 3776 2390 3840
rect 2454 3776 2462 3840
rect 2142 3775 2462 3776
rect 4406 3840 4726 3841
rect 4406 3776 4414 3840
rect 4478 3776 4494 3840
rect 4558 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4726 3840
rect 4406 3775 4726 3776
rect 1010 3296 1330 3297
rect 1010 3232 1018 3296
rect 1082 3232 1098 3296
rect 1162 3232 1178 3296
rect 1242 3232 1258 3296
rect 1322 3232 1330 3296
rect 1010 3231 1330 3232
rect 3274 3296 3594 3297
rect 3274 3232 3282 3296
rect 3346 3232 3362 3296
rect 3426 3232 3442 3296
rect 3506 3232 3522 3296
rect 3586 3232 3594 3296
rect 3274 3231 3594 3232
rect 5538 3296 5858 3297
rect 5538 3232 5546 3296
rect 5610 3232 5626 3296
rect 5690 3232 5706 3296
rect 5770 3232 5786 3296
rect 5850 3232 5858 3296
rect 5538 3231 5858 3232
rect 2142 2752 2462 2753
rect 2142 2688 2150 2752
rect 2214 2688 2230 2752
rect 2294 2688 2310 2752
rect 2374 2688 2390 2752
rect 2454 2688 2462 2752
rect 2142 2687 2462 2688
rect 4406 2752 4726 2753
rect 4406 2688 4414 2752
rect 4478 2688 4494 2752
rect 4558 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4726 2752
rect 4406 2687 4726 2688
rect 5203 2410 5269 2413
rect 5203 2408 6600 2410
rect 5203 2352 5208 2408
rect 5264 2352 6600 2408
rect 5203 2350 6600 2352
rect 5203 2347 5269 2350
rect 1010 2208 1330 2209
rect 1010 2144 1018 2208
rect 1082 2144 1098 2208
rect 1162 2144 1178 2208
rect 1242 2144 1258 2208
rect 1322 2144 1330 2208
rect 1010 2143 1330 2144
rect 3274 2208 3594 2209
rect 3274 2144 3282 2208
rect 3346 2144 3362 2208
rect 3426 2144 3442 2208
rect 3506 2144 3522 2208
rect 3586 2144 3594 2208
rect 3274 2143 3594 2144
rect 5538 2208 5858 2209
rect 5538 2144 5546 2208
rect 5610 2144 5626 2208
rect 5690 2144 5706 2208
rect 5770 2144 5786 2208
rect 5850 2144 5858 2208
rect 5538 2143 5858 2144
rect 6540 2138 6600 2350
rect 7454 2138 7934 2168
rect 6540 2078 7934 2138
rect 7454 2048 7934 2078
<< via3 >>
rect 2150 14716 2214 14720
rect 2150 14660 2154 14716
rect 2154 14660 2210 14716
rect 2210 14660 2214 14716
rect 2150 14656 2214 14660
rect 2230 14716 2294 14720
rect 2230 14660 2234 14716
rect 2234 14660 2290 14716
rect 2290 14660 2294 14716
rect 2230 14656 2294 14660
rect 2310 14716 2374 14720
rect 2310 14660 2314 14716
rect 2314 14660 2370 14716
rect 2370 14660 2374 14716
rect 2310 14656 2374 14660
rect 2390 14716 2454 14720
rect 2390 14660 2394 14716
rect 2394 14660 2450 14716
rect 2450 14660 2454 14716
rect 2390 14656 2454 14660
rect 4414 14716 4478 14720
rect 4414 14660 4418 14716
rect 4418 14660 4474 14716
rect 4474 14660 4478 14716
rect 4414 14656 4478 14660
rect 4494 14716 4558 14720
rect 4494 14660 4498 14716
rect 4498 14660 4554 14716
rect 4554 14660 4558 14716
rect 4494 14656 4558 14660
rect 4574 14716 4638 14720
rect 4574 14660 4578 14716
rect 4578 14660 4634 14716
rect 4634 14660 4638 14716
rect 4574 14656 4638 14660
rect 4654 14716 4718 14720
rect 4654 14660 4658 14716
rect 4658 14660 4714 14716
rect 4714 14660 4718 14716
rect 4654 14656 4718 14660
rect 1018 14172 1082 14176
rect 1018 14116 1022 14172
rect 1022 14116 1078 14172
rect 1078 14116 1082 14172
rect 1018 14112 1082 14116
rect 1098 14172 1162 14176
rect 1098 14116 1102 14172
rect 1102 14116 1158 14172
rect 1158 14116 1162 14172
rect 1098 14112 1162 14116
rect 1178 14172 1242 14176
rect 1178 14116 1182 14172
rect 1182 14116 1238 14172
rect 1238 14116 1242 14172
rect 1178 14112 1242 14116
rect 1258 14172 1322 14176
rect 1258 14116 1262 14172
rect 1262 14116 1318 14172
rect 1318 14116 1322 14172
rect 1258 14112 1322 14116
rect 3282 14172 3346 14176
rect 3282 14116 3286 14172
rect 3286 14116 3342 14172
rect 3342 14116 3346 14172
rect 3282 14112 3346 14116
rect 3362 14172 3426 14176
rect 3362 14116 3366 14172
rect 3366 14116 3422 14172
rect 3422 14116 3426 14172
rect 3362 14112 3426 14116
rect 3442 14172 3506 14176
rect 3442 14116 3446 14172
rect 3446 14116 3502 14172
rect 3502 14116 3506 14172
rect 3442 14112 3506 14116
rect 3522 14172 3586 14176
rect 3522 14116 3526 14172
rect 3526 14116 3582 14172
rect 3582 14116 3586 14172
rect 3522 14112 3586 14116
rect 5546 14172 5610 14176
rect 5546 14116 5550 14172
rect 5550 14116 5606 14172
rect 5606 14116 5610 14172
rect 5546 14112 5610 14116
rect 5626 14172 5690 14176
rect 5626 14116 5630 14172
rect 5630 14116 5686 14172
rect 5686 14116 5690 14172
rect 5626 14112 5690 14116
rect 5706 14172 5770 14176
rect 5706 14116 5710 14172
rect 5710 14116 5766 14172
rect 5766 14116 5770 14172
rect 5706 14112 5770 14116
rect 5786 14172 5850 14176
rect 5786 14116 5790 14172
rect 5790 14116 5846 14172
rect 5846 14116 5850 14172
rect 5786 14112 5850 14116
rect 2150 13628 2214 13632
rect 2150 13572 2154 13628
rect 2154 13572 2210 13628
rect 2210 13572 2214 13628
rect 2150 13568 2214 13572
rect 2230 13628 2294 13632
rect 2230 13572 2234 13628
rect 2234 13572 2290 13628
rect 2290 13572 2294 13628
rect 2230 13568 2294 13572
rect 2310 13628 2374 13632
rect 2310 13572 2314 13628
rect 2314 13572 2370 13628
rect 2370 13572 2374 13628
rect 2310 13568 2374 13572
rect 2390 13628 2454 13632
rect 2390 13572 2394 13628
rect 2394 13572 2450 13628
rect 2450 13572 2454 13628
rect 2390 13568 2454 13572
rect 4414 13628 4478 13632
rect 4414 13572 4418 13628
rect 4418 13572 4474 13628
rect 4474 13572 4478 13628
rect 4414 13568 4478 13572
rect 4494 13628 4558 13632
rect 4494 13572 4498 13628
rect 4498 13572 4554 13628
rect 4554 13572 4558 13628
rect 4494 13568 4558 13572
rect 4574 13628 4638 13632
rect 4574 13572 4578 13628
rect 4578 13572 4634 13628
rect 4634 13572 4638 13628
rect 4574 13568 4638 13572
rect 4654 13628 4718 13632
rect 4654 13572 4658 13628
rect 4658 13572 4714 13628
rect 4714 13572 4718 13628
rect 4654 13568 4718 13572
rect 1018 13084 1082 13088
rect 1018 13028 1022 13084
rect 1022 13028 1078 13084
rect 1078 13028 1082 13084
rect 1018 13024 1082 13028
rect 1098 13084 1162 13088
rect 1098 13028 1102 13084
rect 1102 13028 1158 13084
rect 1158 13028 1162 13084
rect 1098 13024 1162 13028
rect 1178 13084 1242 13088
rect 1178 13028 1182 13084
rect 1182 13028 1238 13084
rect 1238 13028 1242 13084
rect 1178 13024 1242 13028
rect 1258 13084 1322 13088
rect 1258 13028 1262 13084
rect 1262 13028 1318 13084
rect 1318 13028 1322 13084
rect 1258 13024 1322 13028
rect 3282 13084 3346 13088
rect 3282 13028 3286 13084
rect 3286 13028 3342 13084
rect 3342 13028 3346 13084
rect 3282 13024 3346 13028
rect 3362 13084 3426 13088
rect 3362 13028 3366 13084
rect 3366 13028 3422 13084
rect 3422 13028 3426 13084
rect 3362 13024 3426 13028
rect 3442 13084 3506 13088
rect 3442 13028 3446 13084
rect 3446 13028 3502 13084
rect 3502 13028 3506 13084
rect 3442 13024 3506 13028
rect 3522 13084 3586 13088
rect 3522 13028 3526 13084
rect 3526 13028 3582 13084
rect 3582 13028 3586 13084
rect 3522 13024 3586 13028
rect 5546 13084 5610 13088
rect 5546 13028 5550 13084
rect 5550 13028 5606 13084
rect 5606 13028 5610 13084
rect 5546 13024 5610 13028
rect 5626 13084 5690 13088
rect 5626 13028 5630 13084
rect 5630 13028 5686 13084
rect 5686 13028 5690 13084
rect 5626 13024 5690 13028
rect 5706 13084 5770 13088
rect 5706 13028 5710 13084
rect 5710 13028 5766 13084
rect 5766 13028 5770 13084
rect 5706 13024 5770 13028
rect 5786 13084 5850 13088
rect 5786 13028 5790 13084
rect 5790 13028 5846 13084
rect 5846 13028 5850 13084
rect 5786 13024 5850 13028
rect 2150 12540 2214 12544
rect 2150 12484 2154 12540
rect 2154 12484 2210 12540
rect 2210 12484 2214 12540
rect 2150 12480 2214 12484
rect 2230 12540 2294 12544
rect 2230 12484 2234 12540
rect 2234 12484 2290 12540
rect 2290 12484 2294 12540
rect 2230 12480 2294 12484
rect 2310 12540 2374 12544
rect 2310 12484 2314 12540
rect 2314 12484 2370 12540
rect 2370 12484 2374 12540
rect 2310 12480 2374 12484
rect 2390 12540 2454 12544
rect 2390 12484 2394 12540
rect 2394 12484 2450 12540
rect 2450 12484 2454 12540
rect 2390 12480 2454 12484
rect 4414 12540 4478 12544
rect 4414 12484 4418 12540
rect 4418 12484 4474 12540
rect 4474 12484 4478 12540
rect 4414 12480 4478 12484
rect 4494 12540 4558 12544
rect 4494 12484 4498 12540
rect 4498 12484 4554 12540
rect 4554 12484 4558 12540
rect 4494 12480 4558 12484
rect 4574 12540 4638 12544
rect 4574 12484 4578 12540
rect 4578 12484 4634 12540
rect 4634 12484 4638 12540
rect 4574 12480 4638 12484
rect 4654 12540 4718 12544
rect 4654 12484 4658 12540
rect 4658 12484 4714 12540
rect 4714 12484 4718 12540
rect 4654 12480 4718 12484
rect 1018 11996 1082 12000
rect 1018 11940 1022 11996
rect 1022 11940 1078 11996
rect 1078 11940 1082 11996
rect 1018 11936 1082 11940
rect 1098 11996 1162 12000
rect 1098 11940 1102 11996
rect 1102 11940 1158 11996
rect 1158 11940 1162 11996
rect 1098 11936 1162 11940
rect 1178 11996 1242 12000
rect 1178 11940 1182 11996
rect 1182 11940 1238 11996
rect 1238 11940 1242 11996
rect 1178 11936 1242 11940
rect 1258 11996 1322 12000
rect 1258 11940 1262 11996
rect 1262 11940 1318 11996
rect 1318 11940 1322 11996
rect 1258 11936 1322 11940
rect 3282 11996 3346 12000
rect 3282 11940 3286 11996
rect 3286 11940 3342 11996
rect 3342 11940 3346 11996
rect 3282 11936 3346 11940
rect 3362 11996 3426 12000
rect 3362 11940 3366 11996
rect 3366 11940 3422 11996
rect 3422 11940 3426 11996
rect 3362 11936 3426 11940
rect 3442 11996 3506 12000
rect 3442 11940 3446 11996
rect 3446 11940 3502 11996
rect 3502 11940 3506 11996
rect 3442 11936 3506 11940
rect 3522 11996 3586 12000
rect 3522 11940 3526 11996
rect 3526 11940 3582 11996
rect 3582 11940 3586 11996
rect 3522 11936 3586 11940
rect 5546 11996 5610 12000
rect 5546 11940 5550 11996
rect 5550 11940 5606 11996
rect 5606 11940 5610 11996
rect 5546 11936 5610 11940
rect 5626 11996 5690 12000
rect 5626 11940 5630 11996
rect 5630 11940 5686 11996
rect 5686 11940 5690 11996
rect 5626 11936 5690 11940
rect 5706 11996 5770 12000
rect 5706 11940 5710 11996
rect 5710 11940 5766 11996
rect 5766 11940 5770 11996
rect 5706 11936 5770 11940
rect 5786 11996 5850 12000
rect 5786 11940 5790 11996
rect 5790 11940 5846 11996
rect 5846 11940 5850 11996
rect 5786 11936 5850 11940
rect 2150 11452 2214 11456
rect 2150 11396 2154 11452
rect 2154 11396 2210 11452
rect 2210 11396 2214 11452
rect 2150 11392 2214 11396
rect 2230 11452 2294 11456
rect 2230 11396 2234 11452
rect 2234 11396 2290 11452
rect 2290 11396 2294 11452
rect 2230 11392 2294 11396
rect 2310 11452 2374 11456
rect 2310 11396 2314 11452
rect 2314 11396 2370 11452
rect 2370 11396 2374 11452
rect 2310 11392 2374 11396
rect 2390 11452 2454 11456
rect 2390 11396 2394 11452
rect 2394 11396 2450 11452
rect 2450 11396 2454 11452
rect 2390 11392 2454 11396
rect 4414 11452 4478 11456
rect 4414 11396 4418 11452
rect 4418 11396 4474 11452
rect 4474 11396 4478 11452
rect 4414 11392 4478 11396
rect 4494 11452 4558 11456
rect 4494 11396 4498 11452
rect 4498 11396 4554 11452
rect 4554 11396 4558 11452
rect 4494 11392 4558 11396
rect 4574 11452 4638 11456
rect 4574 11396 4578 11452
rect 4578 11396 4634 11452
rect 4634 11396 4638 11452
rect 4574 11392 4638 11396
rect 4654 11452 4718 11456
rect 4654 11396 4658 11452
rect 4658 11396 4714 11452
rect 4714 11396 4718 11452
rect 4654 11392 4718 11396
rect 1018 10908 1082 10912
rect 1018 10852 1022 10908
rect 1022 10852 1078 10908
rect 1078 10852 1082 10908
rect 1018 10848 1082 10852
rect 1098 10908 1162 10912
rect 1098 10852 1102 10908
rect 1102 10852 1158 10908
rect 1158 10852 1162 10908
rect 1098 10848 1162 10852
rect 1178 10908 1242 10912
rect 1178 10852 1182 10908
rect 1182 10852 1238 10908
rect 1238 10852 1242 10908
rect 1178 10848 1242 10852
rect 1258 10908 1322 10912
rect 1258 10852 1262 10908
rect 1262 10852 1318 10908
rect 1318 10852 1322 10908
rect 1258 10848 1322 10852
rect 3282 10908 3346 10912
rect 3282 10852 3286 10908
rect 3286 10852 3342 10908
rect 3342 10852 3346 10908
rect 3282 10848 3346 10852
rect 3362 10908 3426 10912
rect 3362 10852 3366 10908
rect 3366 10852 3422 10908
rect 3422 10852 3426 10908
rect 3362 10848 3426 10852
rect 3442 10908 3506 10912
rect 3442 10852 3446 10908
rect 3446 10852 3502 10908
rect 3502 10852 3506 10908
rect 3442 10848 3506 10852
rect 3522 10908 3586 10912
rect 3522 10852 3526 10908
rect 3526 10852 3582 10908
rect 3582 10852 3586 10908
rect 3522 10848 3586 10852
rect 5546 10908 5610 10912
rect 5546 10852 5550 10908
rect 5550 10852 5606 10908
rect 5606 10852 5610 10908
rect 5546 10848 5610 10852
rect 5626 10908 5690 10912
rect 5626 10852 5630 10908
rect 5630 10852 5686 10908
rect 5686 10852 5690 10908
rect 5626 10848 5690 10852
rect 5706 10908 5770 10912
rect 5706 10852 5710 10908
rect 5710 10852 5766 10908
rect 5766 10852 5770 10908
rect 5706 10848 5770 10852
rect 5786 10908 5850 10912
rect 5786 10852 5790 10908
rect 5790 10852 5846 10908
rect 5846 10852 5850 10908
rect 5786 10848 5850 10852
rect 2150 10364 2214 10368
rect 2150 10308 2154 10364
rect 2154 10308 2210 10364
rect 2210 10308 2214 10364
rect 2150 10304 2214 10308
rect 2230 10364 2294 10368
rect 2230 10308 2234 10364
rect 2234 10308 2290 10364
rect 2290 10308 2294 10364
rect 2230 10304 2294 10308
rect 2310 10364 2374 10368
rect 2310 10308 2314 10364
rect 2314 10308 2370 10364
rect 2370 10308 2374 10364
rect 2310 10304 2374 10308
rect 2390 10364 2454 10368
rect 2390 10308 2394 10364
rect 2394 10308 2450 10364
rect 2450 10308 2454 10364
rect 2390 10304 2454 10308
rect 4414 10364 4478 10368
rect 4414 10308 4418 10364
rect 4418 10308 4474 10364
rect 4474 10308 4478 10364
rect 4414 10304 4478 10308
rect 4494 10364 4558 10368
rect 4494 10308 4498 10364
rect 4498 10308 4554 10364
rect 4554 10308 4558 10364
rect 4494 10304 4558 10308
rect 4574 10364 4638 10368
rect 4574 10308 4578 10364
rect 4578 10308 4634 10364
rect 4634 10308 4638 10364
rect 4574 10304 4638 10308
rect 4654 10364 4718 10368
rect 4654 10308 4658 10364
rect 4658 10308 4714 10364
rect 4714 10308 4718 10364
rect 4654 10304 4718 10308
rect 1018 9820 1082 9824
rect 1018 9764 1022 9820
rect 1022 9764 1078 9820
rect 1078 9764 1082 9820
rect 1018 9760 1082 9764
rect 1098 9820 1162 9824
rect 1098 9764 1102 9820
rect 1102 9764 1158 9820
rect 1158 9764 1162 9820
rect 1098 9760 1162 9764
rect 1178 9820 1242 9824
rect 1178 9764 1182 9820
rect 1182 9764 1238 9820
rect 1238 9764 1242 9820
rect 1178 9760 1242 9764
rect 1258 9820 1322 9824
rect 1258 9764 1262 9820
rect 1262 9764 1318 9820
rect 1318 9764 1322 9820
rect 1258 9760 1322 9764
rect 3282 9820 3346 9824
rect 3282 9764 3286 9820
rect 3286 9764 3342 9820
rect 3342 9764 3346 9820
rect 3282 9760 3346 9764
rect 3362 9820 3426 9824
rect 3362 9764 3366 9820
rect 3366 9764 3422 9820
rect 3422 9764 3426 9820
rect 3362 9760 3426 9764
rect 3442 9820 3506 9824
rect 3442 9764 3446 9820
rect 3446 9764 3502 9820
rect 3502 9764 3506 9820
rect 3442 9760 3506 9764
rect 3522 9820 3586 9824
rect 3522 9764 3526 9820
rect 3526 9764 3582 9820
rect 3582 9764 3586 9820
rect 3522 9760 3586 9764
rect 5546 9820 5610 9824
rect 5546 9764 5550 9820
rect 5550 9764 5606 9820
rect 5606 9764 5610 9820
rect 5546 9760 5610 9764
rect 5626 9820 5690 9824
rect 5626 9764 5630 9820
rect 5630 9764 5686 9820
rect 5686 9764 5690 9820
rect 5626 9760 5690 9764
rect 5706 9820 5770 9824
rect 5706 9764 5710 9820
rect 5710 9764 5766 9820
rect 5766 9764 5770 9820
rect 5706 9760 5770 9764
rect 5786 9820 5850 9824
rect 5786 9764 5790 9820
rect 5790 9764 5846 9820
rect 5846 9764 5850 9820
rect 5786 9760 5850 9764
rect 2150 9276 2214 9280
rect 2150 9220 2154 9276
rect 2154 9220 2210 9276
rect 2210 9220 2214 9276
rect 2150 9216 2214 9220
rect 2230 9276 2294 9280
rect 2230 9220 2234 9276
rect 2234 9220 2290 9276
rect 2290 9220 2294 9276
rect 2230 9216 2294 9220
rect 2310 9276 2374 9280
rect 2310 9220 2314 9276
rect 2314 9220 2370 9276
rect 2370 9220 2374 9276
rect 2310 9216 2374 9220
rect 2390 9276 2454 9280
rect 2390 9220 2394 9276
rect 2394 9220 2450 9276
rect 2450 9220 2454 9276
rect 2390 9216 2454 9220
rect 4414 9276 4478 9280
rect 4414 9220 4418 9276
rect 4418 9220 4474 9276
rect 4474 9220 4478 9276
rect 4414 9216 4478 9220
rect 4494 9276 4558 9280
rect 4494 9220 4498 9276
rect 4498 9220 4554 9276
rect 4554 9220 4558 9276
rect 4494 9216 4558 9220
rect 4574 9276 4638 9280
rect 4574 9220 4578 9276
rect 4578 9220 4634 9276
rect 4634 9220 4638 9276
rect 4574 9216 4638 9220
rect 4654 9276 4718 9280
rect 4654 9220 4658 9276
rect 4658 9220 4714 9276
rect 4714 9220 4718 9276
rect 4654 9216 4718 9220
rect 1018 8732 1082 8736
rect 1018 8676 1022 8732
rect 1022 8676 1078 8732
rect 1078 8676 1082 8732
rect 1018 8672 1082 8676
rect 1098 8732 1162 8736
rect 1098 8676 1102 8732
rect 1102 8676 1158 8732
rect 1158 8676 1162 8732
rect 1098 8672 1162 8676
rect 1178 8732 1242 8736
rect 1178 8676 1182 8732
rect 1182 8676 1238 8732
rect 1238 8676 1242 8732
rect 1178 8672 1242 8676
rect 1258 8732 1322 8736
rect 1258 8676 1262 8732
rect 1262 8676 1318 8732
rect 1318 8676 1322 8732
rect 1258 8672 1322 8676
rect 3282 8732 3346 8736
rect 3282 8676 3286 8732
rect 3286 8676 3342 8732
rect 3342 8676 3346 8732
rect 3282 8672 3346 8676
rect 3362 8732 3426 8736
rect 3362 8676 3366 8732
rect 3366 8676 3422 8732
rect 3422 8676 3426 8732
rect 3362 8672 3426 8676
rect 3442 8732 3506 8736
rect 3442 8676 3446 8732
rect 3446 8676 3502 8732
rect 3502 8676 3506 8732
rect 3442 8672 3506 8676
rect 3522 8732 3586 8736
rect 3522 8676 3526 8732
rect 3526 8676 3582 8732
rect 3582 8676 3586 8732
rect 3522 8672 3586 8676
rect 5546 8732 5610 8736
rect 5546 8676 5550 8732
rect 5550 8676 5606 8732
rect 5606 8676 5610 8732
rect 5546 8672 5610 8676
rect 5626 8732 5690 8736
rect 5626 8676 5630 8732
rect 5630 8676 5686 8732
rect 5686 8676 5690 8732
rect 5626 8672 5690 8676
rect 5706 8732 5770 8736
rect 5706 8676 5710 8732
rect 5710 8676 5766 8732
rect 5766 8676 5770 8732
rect 5706 8672 5770 8676
rect 5786 8732 5850 8736
rect 5786 8676 5790 8732
rect 5790 8676 5846 8732
rect 5846 8676 5850 8732
rect 5786 8672 5850 8676
rect 2150 8188 2214 8192
rect 2150 8132 2154 8188
rect 2154 8132 2210 8188
rect 2210 8132 2214 8188
rect 2150 8128 2214 8132
rect 2230 8188 2294 8192
rect 2230 8132 2234 8188
rect 2234 8132 2290 8188
rect 2290 8132 2294 8188
rect 2230 8128 2294 8132
rect 2310 8188 2374 8192
rect 2310 8132 2314 8188
rect 2314 8132 2370 8188
rect 2370 8132 2374 8188
rect 2310 8128 2374 8132
rect 2390 8188 2454 8192
rect 2390 8132 2394 8188
rect 2394 8132 2450 8188
rect 2450 8132 2454 8188
rect 2390 8128 2454 8132
rect 4414 8188 4478 8192
rect 4414 8132 4418 8188
rect 4418 8132 4474 8188
rect 4474 8132 4478 8188
rect 4414 8128 4478 8132
rect 4494 8188 4558 8192
rect 4494 8132 4498 8188
rect 4498 8132 4554 8188
rect 4554 8132 4558 8188
rect 4494 8128 4558 8132
rect 4574 8188 4638 8192
rect 4574 8132 4578 8188
rect 4578 8132 4634 8188
rect 4634 8132 4638 8188
rect 4574 8128 4638 8132
rect 4654 8188 4718 8192
rect 4654 8132 4658 8188
rect 4658 8132 4714 8188
rect 4714 8132 4718 8188
rect 4654 8128 4718 8132
rect 1018 7644 1082 7648
rect 1018 7588 1022 7644
rect 1022 7588 1078 7644
rect 1078 7588 1082 7644
rect 1018 7584 1082 7588
rect 1098 7644 1162 7648
rect 1098 7588 1102 7644
rect 1102 7588 1158 7644
rect 1158 7588 1162 7644
rect 1098 7584 1162 7588
rect 1178 7644 1242 7648
rect 1178 7588 1182 7644
rect 1182 7588 1238 7644
rect 1238 7588 1242 7644
rect 1178 7584 1242 7588
rect 1258 7644 1322 7648
rect 1258 7588 1262 7644
rect 1262 7588 1318 7644
rect 1318 7588 1322 7644
rect 1258 7584 1322 7588
rect 3282 7644 3346 7648
rect 3282 7588 3286 7644
rect 3286 7588 3342 7644
rect 3342 7588 3346 7644
rect 3282 7584 3346 7588
rect 3362 7644 3426 7648
rect 3362 7588 3366 7644
rect 3366 7588 3422 7644
rect 3422 7588 3426 7644
rect 3362 7584 3426 7588
rect 3442 7644 3506 7648
rect 3442 7588 3446 7644
rect 3446 7588 3502 7644
rect 3502 7588 3506 7644
rect 3442 7584 3506 7588
rect 3522 7644 3586 7648
rect 3522 7588 3526 7644
rect 3526 7588 3582 7644
rect 3582 7588 3586 7644
rect 3522 7584 3586 7588
rect 5546 7644 5610 7648
rect 5546 7588 5550 7644
rect 5550 7588 5606 7644
rect 5606 7588 5610 7644
rect 5546 7584 5610 7588
rect 5626 7644 5690 7648
rect 5626 7588 5630 7644
rect 5630 7588 5686 7644
rect 5686 7588 5690 7644
rect 5626 7584 5690 7588
rect 5706 7644 5770 7648
rect 5706 7588 5710 7644
rect 5710 7588 5766 7644
rect 5766 7588 5770 7644
rect 5706 7584 5770 7588
rect 5786 7644 5850 7648
rect 5786 7588 5790 7644
rect 5790 7588 5846 7644
rect 5846 7588 5850 7644
rect 5786 7584 5850 7588
rect 2150 7100 2214 7104
rect 2150 7044 2154 7100
rect 2154 7044 2210 7100
rect 2210 7044 2214 7100
rect 2150 7040 2214 7044
rect 2230 7100 2294 7104
rect 2230 7044 2234 7100
rect 2234 7044 2290 7100
rect 2290 7044 2294 7100
rect 2230 7040 2294 7044
rect 2310 7100 2374 7104
rect 2310 7044 2314 7100
rect 2314 7044 2370 7100
rect 2370 7044 2374 7100
rect 2310 7040 2374 7044
rect 2390 7100 2454 7104
rect 2390 7044 2394 7100
rect 2394 7044 2450 7100
rect 2450 7044 2454 7100
rect 2390 7040 2454 7044
rect 4414 7100 4478 7104
rect 4414 7044 4418 7100
rect 4418 7044 4474 7100
rect 4474 7044 4478 7100
rect 4414 7040 4478 7044
rect 4494 7100 4558 7104
rect 4494 7044 4498 7100
rect 4498 7044 4554 7100
rect 4554 7044 4558 7100
rect 4494 7040 4558 7044
rect 4574 7100 4638 7104
rect 4574 7044 4578 7100
rect 4578 7044 4634 7100
rect 4634 7044 4638 7100
rect 4574 7040 4638 7044
rect 4654 7100 4718 7104
rect 4654 7044 4658 7100
rect 4658 7044 4714 7100
rect 4714 7044 4718 7100
rect 4654 7040 4718 7044
rect 1018 6556 1082 6560
rect 1018 6500 1022 6556
rect 1022 6500 1078 6556
rect 1078 6500 1082 6556
rect 1018 6496 1082 6500
rect 1098 6556 1162 6560
rect 1098 6500 1102 6556
rect 1102 6500 1158 6556
rect 1158 6500 1162 6556
rect 1098 6496 1162 6500
rect 1178 6556 1242 6560
rect 1178 6500 1182 6556
rect 1182 6500 1238 6556
rect 1238 6500 1242 6556
rect 1178 6496 1242 6500
rect 1258 6556 1322 6560
rect 1258 6500 1262 6556
rect 1262 6500 1318 6556
rect 1318 6500 1322 6556
rect 1258 6496 1322 6500
rect 3282 6556 3346 6560
rect 3282 6500 3286 6556
rect 3286 6500 3342 6556
rect 3342 6500 3346 6556
rect 3282 6496 3346 6500
rect 3362 6556 3426 6560
rect 3362 6500 3366 6556
rect 3366 6500 3422 6556
rect 3422 6500 3426 6556
rect 3362 6496 3426 6500
rect 3442 6556 3506 6560
rect 3442 6500 3446 6556
rect 3446 6500 3502 6556
rect 3502 6500 3506 6556
rect 3442 6496 3506 6500
rect 3522 6556 3586 6560
rect 3522 6500 3526 6556
rect 3526 6500 3582 6556
rect 3582 6500 3586 6556
rect 3522 6496 3586 6500
rect 5546 6556 5610 6560
rect 5546 6500 5550 6556
rect 5550 6500 5606 6556
rect 5606 6500 5610 6556
rect 5546 6496 5610 6500
rect 5626 6556 5690 6560
rect 5626 6500 5630 6556
rect 5630 6500 5686 6556
rect 5686 6500 5690 6556
rect 5626 6496 5690 6500
rect 5706 6556 5770 6560
rect 5706 6500 5710 6556
rect 5710 6500 5766 6556
rect 5766 6500 5770 6556
rect 5706 6496 5770 6500
rect 5786 6556 5850 6560
rect 5786 6500 5790 6556
rect 5790 6500 5846 6556
rect 5846 6500 5850 6556
rect 5786 6496 5850 6500
rect 2150 6012 2214 6016
rect 2150 5956 2154 6012
rect 2154 5956 2210 6012
rect 2210 5956 2214 6012
rect 2150 5952 2214 5956
rect 2230 6012 2294 6016
rect 2230 5956 2234 6012
rect 2234 5956 2290 6012
rect 2290 5956 2294 6012
rect 2230 5952 2294 5956
rect 2310 6012 2374 6016
rect 2310 5956 2314 6012
rect 2314 5956 2370 6012
rect 2370 5956 2374 6012
rect 2310 5952 2374 5956
rect 2390 6012 2454 6016
rect 2390 5956 2394 6012
rect 2394 5956 2450 6012
rect 2450 5956 2454 6012
rect 2390 5952 2454 5956
rect 4414 6012 4478 6016
rect 4414 5956 4418 6012
rect 4418 5956 4474 6012
rect 4474 5956 4478 6012
rect 4414 5952 4478 5956
rect 4494 6012 4558 6016
rect 4494 5956 4498 6012
rect 4498 5956 4554 6012
rect 4554 5956 4558 6012
rect 4494 5952 4558 5956
rect 4574 6012 4638 6016
rect 4574 5956 4578 6012
rect 4578 5956 4634 6012
rect 4634 5956 4638 6012
rect 4574 5952 4638 5956
rect 4654 6012 4718 6016
rect 4654 5956 4658 6012
rect 4658 5956 4714 6012
rect 4714 5956 4718 6012
rect 4654 5952 4718 5956
rect 1018 5468 1082 5472
rect 1018 5412 1022 5468
rect 1022 5412 1078 5468
rect 1078 5412 1082 5468
rect 1018 5408 1082 5412
rect 1098 5468 1162 5472
rect 1098 5412 1102 5468
rect 1102 5412 1158 5468
rect 1158 5412 1162 5468
rect 1098 5408 1162 5412
rect 1178 5468 1242 5472
rect 1178 5412 1182 5468
rect 1182 5412 1238 5468
rect 1238 5412 1242 5468
rect 1178 5408 1242 5412
rect 1258 5468 1322 5472
rect 1258 5412 1262 5468
rect 1262 5412 1318 5468
rect 1318 5412 1322 5468
rect 1258 5408 1322 5412
rect 3282 5468 3346 5472
rect 3282 5412 3286 5468
rect 3286 5412 3342 5468
rect 3342 5412 3346 5468
rect 3282 5408 3346 5412
rect 3362 5468 3426 5472
rect 3362 5412 3366 5468
rect 3366 5412 3422 5468
rect 3422 5412 3426 5468
rect 3362 5408 3426 5412
rect 3442 5468 3506 5472
rect 3442 5412 3446 5468
rect 3446 5412 3502 5468
rect 3502 5412 3506 5468
rect 3442 5408 3506 5412
rect 3522 5468 3586 5472
rect 3522 5412 3526 5468
rect 3526 5412 3582 5468
rect 3582 5412 3586 5468
rect 3522 5408 3586 5412
rect 5546 5468 5610 5472
rect 5546 5412 5550 5468
rect 5550 5412 5606 5468
rect 5606 5412 5610 5468
rect 5546 5408 5610 5412
rect 5626 5468 5690 5472
rect 5626 5412 5630 5468
rect 5630 5412 5686 5468
rect 5686 5412 5690 5468
rect 5626 5408 5690 5412
rect 5706 5468 5770 5472
rect 5706 5412 5710 5468
rect 5710 5412 5766 5468
rect 5766 5412 5770 5468
rect 5706 5408 5770 5412
rect 5786 5468 5850 5472
rect 5786 5412 5790 5468
rect 5790 5412 5846 5468
rect 5846 5412 5850 5468
rect 5786 5408 5850 5412
rect 2150 4924 2214 4928
rect 2150 4868 2154 4924
rect 2154 4868 2210 4924
rect 2210 4868 2214 4924
rect 2150 4864 2214 4868
rect 2230 4924 2294 4928
rect 2230 4868 2234 4924
rect 2234 4868 2290 4924
rect 2290 4868 2294 4924
rect 2230 4864 2294 4868
rect 2310 4924 2374 4928
rect 2310 4868 2314 4924
rect 2314 4868 2370 4924
rect 2370 4868 2374 4924
rect 2310 4864 2374 4868
rect 2390 4924 2454 4928
rect 2390 4868 2394 4924
rect 2394 4868 2450 4924
rect 2450 4868 2454 4924
rect 2390 4864 2454 4868
rect 4414 4924 4478 4928
rect 4414 4868 4418 4924
rect 4418 4868 4474 4924
rect 4474 4868 4478 4924
rect 4414 4864 4478 4868
rect 4494 4924 4558 4928
rect 4494 4868 4498 4924
rect 4498 4868 4554 4924
rect 4554 4868 4558 4924
rect 4494 4864 4558 4868
rect 4574 4924 4638 4928
rect 4574 4868 4578 4924
rect 4578 4868 4634 4924
rect 4634 4868 4638 4924
rect 4574 4864 4638 4868
rect 4654 4924 4718 4928
rect 4654 4868 4658 4924
rect 4658 4868 4714 4924
rect 4714 4868 4718 4924
rect 4654 4864 4718 4868
rect 1018 4380 1082 4384
rect 1018 4324 1022 4380
rect 1022 4324 1078 4380
rect 1078 4324 1082 4380
rect 1018 4320 1082 4324
rect 1098 4380 1162 4384
rect 1098 4324 1102 4380
rect 1102 4324 1158 4380
rect 1158 4324 1162 4380
rect 1098 4320 1162 4324
rect 1178 4380 1242 4384
rect 1178 4324 1182 4380
rect 1182 4324 1238 4380
rect 1238 4324 1242 4380
rect 1178 4320 1242 4324
rect 1258 4380 1322 4384
rect 1258 4324 1262 4380
rect 1262 4324 1318 4380
rect 1318 4324 1322 4380
rect 1258 4320 1322 4324
rect 3282 4380 3346 4384
rect 3282 4324 3286 4380
rect 3286 4324 3342 4380
rect 3342 4324 3346 4380
rect 3282 4320 3346 4324
rect 3362 4380 3426 4384
rect 3362 4324 3366 4380
rect 3366 4324 3422 4380
rect 3422 4324 3426 4380
rect 3362 4320 3426 4324
rect 3442 4380 3506 4384
rect 3442 4324 3446 4380
rect 3446 4324 3502 4380
rect 3502 4324 3506 4380
rect 3442 4320 3506 4324
rect 3522 4380 3586 4384
rect 3522 4324 3526 4380
rect 3526 4324 3582 4380
rect 3582 4324 3586 4380
rect 3522 4320 3586 4324
rect 5546 4380 5610 4384
rect 5546 4324 5550 4380
rect 5550 4324 5606 4380
rect 5606 4324 5610 4380
rect 5546 4320 5610 4324
rect 5626 4380 5690 4384
rect 5626 4324 5630 4380
rect 5630 4324 5686 4380
rect 5686 4324 5690 4380
rect 5626 4320 5690 4324
rect 5706 4380 5770 4384
rect 5706 4324 5710 4380
rect 5710 4324 5766 4380
rect 5766 4324 5770 4380
rect 5706 4320 5770 4324
rect 5786 4380 5850 4384
rect 5786 4324 5790 4380
rect 5790 4324 5846 4380
rect 5846 4324 5850 4380
rect 5786 4320 5850 4324
rect 2150 3836 2214 3840
rect 2150 3780 2154 3836
rect 2154 3780 2210 3836
rect 2210 3780 2214 3836
rect 2150 3776 2214 3780
rect 2230 3836 2294 3840
rect 2230 3780 2234 3836
rect 2234 3780 2290 3836
rect 2290 3780 2294 3836
rect 2230 3776 2294 3780
rect 2310 3836 2374 3840
rect 2310 3780 2314 3836
rect 2314 3780 2370 3836
rect 2370 3780 2374 3836
rect 2310 3776 2374 3780
rect 2390 3836 2454 3840
rect 2390 3780 2394 3836
rect 2394 3780 2450 3836
rect 2450 3780 2454 3836
rect 2390 3776 2454 3780
rect 4414 3836 4478 3840
rect 4414 3780 4418 3836
rect 4418 3780 4474 3836
rect 4474 3780 4478 3836
rect 4414 3776 4478 3780
rect 4494 3836 4558 3840
rect 4494 3780 4498 3836
rect 4498 3780 4554 3836
rect 4554 3780 4558 3836
rect 4494 3776 4558 3780
rect 4574 3836 4638 3840
rect 4574 3780 4578 3836
rect 4578 3780 4634 3836
rect 4634 3780 4638 3836
rect 4574 3776 4638 3780
rect 4654 3836 4718 3840
rect 4654 3780 4658 3836
rect 4658 3780 4714 3836
rect 4714 3780 4718 3836
rect 4654 3776 4718 3780
rect 1018 3292 1082 3296
rect 1018 3236 1022 3292
rect 1022 3236 1078 3292
rect 1078 3236 1082 3292
rect 1018 3232 1082 3236
rect 1098 3292 1162 3296
rect 1098 3236 1102 3292
rect 1102 3236 1158 3292
rect 1158 3236 1162 3292
rect 1098 3232 1162 3236
rect 1178 3292 1242 3296
rect 1178 3236 1182 3292
rect 1182 3236 1238 3292
rect 1238 3236 1242 3292
rect 1178 3232 1242 3236
rect 1258 3292 1322 3296
rect 1258 3236 1262 3292
rect 1262 3236 1318 3292
rect 1318 3236 1322 3292
rect 1258 3232 1322 3236
rect 3282 3292 3346 3296
rect 3282 3236 3286 3292
rect 3286 3236 3342 3292
rect 3342 3236 3346 3292
rect 3282 3232 3346 3236
rect 3362 3292 3426 3296
rect 3362 3236 3366 3292
rect 3366 3236 3422 3292
rect 3422 3236 3426 3292
rect 3362 3232 3426 3236
rect 3442 3292 3506 3296
rect 3442 3236 3446 3292
rect 3446 3236 3502 3292
rect 3502 3236 3506 3292
rect 3442 3232 3506 3236
rect 3522 3292 3586 3296
rect 3522 3236 3526 3292
rect 3526 3236 3582 3292
rect 3582 3236 3586 3292
rect 3522 3232 3586 3236
rect 5546 3292 5610 3296
rect 5546 3236 5550 3292
rect 5550 3236 5606 3292
rect 5606 3236 5610 3292
rect 5546 3232 5610 3236
rect 5626 3292 5690 3296
rect 5626 3236 5630 3292
rect 5630 3236 5686 3292
rect 5686 3236 5690 3292
rect 5626 3232 5690 3236
rect 5706 3292 5770 3296
rect 5706 3236 5710 3292
rect 5710 3236 5766 3292
rect 5766 3236 5770 3292
rect 5706 3232 5770 3236
rect 5786 3292 5850 3296
rect 5786 3236 5790 3292
rect 5790 3236 5846 3292
rect 5846 3236 5850 3292
rect 5786 3232 5850 3236
rect 2150 2748 2214 2752
rect 2150 2692 2154 2748
rect 2154 2692 2210 2748
rect 2210 2692 2214 2748
rect 2150 2688 2214 2692
rect 2230 2748 2294 2752
rect 2230 2692 2234 2748
rect 2234 2692 2290 2748
rect 2290 2692 2294 2748
rect 2230 2688 2294 2692
rect 2310 2748 2374 2752
rect 2310 2692 2314 2748
rect 2314 2692 2370 2748
rect 2370 2692 2374 2748
rect 2310 2688 2374 2692
rect 2390 2748 2454 2752
rect 2390 2692 2394 2748
rect 2394 2692 2450 2748
rect 2450 2692 2454 2748
rect 2390 2688 2454 2692
rect 4414 2748 4478 2752
rect 4414 2692 4418 2748
rect 4418 2692 4474 2748
rect 4474 2692 4478 2748
rect 4414 2688 4478 2692
rect 4494 2748 4558 2752
rect 4494 2692 4498 2748
rect 4498 2692 4554 2748
rect 4554 2692 4558 2748
rect 4494 2688 4558 2692
rect 4574 2748 4638 2752
rect 4574 2692 4578 2748
rect 4578 2692 4634 2748
rect 4634 2692 4638 2748
rect 4574 2688 4638 2692
rect 4654 2748 4718 2752
rect 4654 2692 4658 2748
rect 4658 2692 4714 2748
rect 4714 2692 4718 2748
rect 4654 2688 4718 2692
rect 1018 2204 1082 2208
rect 1018 2148 1022 2204
rect 1022 2148 1078 2204
rect 1078 2148 1082 2204
rect 1018 2144 1082 2148
rect 1098 2204 1162 2208
rect 1098 2148 1102 2204
rect 1102 2148 1158 2204
rect 1158 2148 1162 2204
rect 1098 2144 1162 2148
rect 1178 2204 1242 2208
rect 1178 2148 1182 2204
rect 1182 2148 1238 2204
rect 1238 2148 1242 2204
rect 1178 2144 1242 2148
rect 1258 2204 1322 2208
rect 1258 2148 1262 2204
rect 1262 2148 1318 2204
rect 1318 2148 1322 2204
rect 1258 2144 1322 2148
rect 3282 2204 3346 2208
rect 3282 2148 3286 2204
rect 3286 2148 3342 2204
rect 3342 2148 3346 2204
rect 3282 2144 3346 2148
rect 3362 2204 3426 2208
rect 3362 2148 3366 2204
rect 3366 2148 3422 2204
rect 3422 2148 3426 2204
rect 3362 2144 3426 2148
rect 3442 2204 3506 2208
rect 3442 2148 3446 2204
rect 3446 2148 3502 2204
rect 3502 2148 3506 2204
rect 3442 2144 3506 2148
rect 3522 2204 3586 2208
rect 3522 2148 3526 2204
rect 3526 2148 3582 2204
rect 3582 2148 3586 2204
rect 3522 2144 3586 2148
rect 5546 2204 5610 2208
rect 5546 2148 5550 2204
rect 5550 2148 5606 2204
rect 5606 2148 5610 2204
rect 5546 2144 5610 2148
rect 5626 2204 5690 2208
rect 5626 2148 5630 2204
rect 5630 2148 5686 2204
rect 5686 2148 5690 2204
rect 5626 2144 5690 2148
rect 5706 2204 5770 2208
rect 5706 2148 5710 2204
rect 5710 2148 5766 2204
rect 5766 2148 5770 2204
rect 5706 2144 5770 2148
rect 5786 2204 5850 2208
rect 5786 2148 5790 2204
rect 5790 2148 5846 2204
rect 5846 2148 5850 2204
rect 5786 2144 5850 2148
<< metal4 >>
rect 1010 14176 1330 14736
rect 1010 14112 1018 14176
rect 1082 14112 1098 14176
rect 1162 14112 1178 14176
rect 1242 14112 1258 14176
rect 1322 14112 1330 14176
rect 1010 13088 1330 14112
rect 1010 13024 1018 13088
rect 1082 13024 1098 13088
rect 1162 13024 1178 13088
rect 1242 13024 1258 13088
rect 1322 13024 1330 13088
rect 1010 12000 1330 13024
rect 1010 11936 1018 12000
rect 1082 11936 1098 12000
rect 1162 11936 1178 12000
rect 1242 11936 1258 12000
rect 1322 11936 1330 12000
rect 1010 10912 1330 11936
rect 1010 10848 1018 10912
rect 1082 10848 1098 10912
rect 1162 10848 1178 10912
rect 1242 10848 1258 10912
rect 1322 10848 1330 10912
rect 1010 9824 1330 10848
rect 1010 9760 1018 9824
rect 1082 9760 1098 9824
rect 1162 9760 1178 9824
rect 1242 9760 1258 9824
rect 1322 9760 1330 9824
rect 1010 8736 1330 9760
rect 1010 8672 1018 8736
rect 1082 8672 1098 8736
rect 1162 8672 1178 8736
rect 1242 8672 1258 8736
rect 1322 8672 1330 8736
rect 1010 7648 1330 8672
rect 1010 7584 1018 7648
rect 1082 7584 1098 7648
rect 1162 7584 1178 7648
rect 1242 7584 1258 7648
rect 1322 7584 1330 7648
rect 1010 6560 1330 7584
rect 1010 6496 1018 6560
rect 1082 6496 1098 6560
rect 1162 6496 1178 6560
rect 1242 6496 1258 6560
rect 1322 6496 1330 6560
rect 1010 5472 1330 6496
rect 1010 5408 1018 5472
rect 1082 5408 1098 5472
rect 1162 5408 1178 5472
rect 1242 5408 1258 5472
rect 1322 5408 1330 5472
rect 1010 4384 1330 5408
rect 1010 4320 1018 4384
rect 1082 4320 1098 4384
rect 1162 4320 1178 4384
rect 1242 4320 1258 4384
rect 1322 4320 1330 4384
rect 1010 3296 1330 4320
rect 1010 3232 1018 3296
rect 1082 3232 1098 3296
rect 1162 3232 1178 3296
rect 1242 3232 1258 3296
rect 1322 3232 1330 3296
rect 1010 2208 1330 3232
rect 1010 2144 1018 2208
rect 1082 2144 1098 2208
rect 1162 2144 1178 2208
rect 1242 2144 1258 2208
rect 1322 2144 1330 2208
rect 1010 2128 1330 2144
rect 2142 14720 2462 14736
rect 2142 14656 2150 14720
rect 2214 14656 2230 14720
rect 2294 14656 2310 14720
rect 2374 14656 2390 14720
rect 2454 14656 2462 14720
rect 2142 13632 2462 14656
rect 2142 13568 2150 13632
rect 2214 13568 2230 13632
rect 2294 13568 2310 13632
rect 2374 13568 2390 13632
rect 2454 13568 2462 13632
rect 2142 12544 2462 13568
rect 2142 12480 2150 12544
rect 2214 12480 2230 12544
rect 2294 12480 2310 12544
rect 2374 12480 2390 12544
rect 2454 12480 2462 12544
rect 2142 11456 2462 12480
rect 2142 11392 2150 11456
rect 2214 11392 2230 11456
rect 2294 11392 2310 11456
rect 2374 11392 2390 11456
rect 2454 11392 2462 11456
rect 2142 10368 2462 11392
rect 2142 10304 2150 10368
rect 2214 10304 2230 10368
rect 2294 10304 2310 10368
rect 2374 10304 2390 10368
rect 2454 10304 2462 10368
rect 2142 9280 2462 10304
rect 2142 9216 2150 9280
rect 2214 9216 2230 9280
rect 2294 9216 2310 9280
rect 2374 9216 2390 9280
rect 2454 9216 2462 9280
rect 2142 8192 2462 9216
rect 2142 8128 2150 8192
rect 2214 8128 2230 8192
rect 2294 8128 2310 8192
rect 2374 8128 2390 8192
rect 2454 8128 2462 8192
rect 2142 7104 2462 8128
rect 2142 7040 2150 7104
rect 2214 7040 2230 7104
rect 2294 7040 2310 7104
rect 2374 7040 2390 7104
rect 2454 7040 2462 7104
rect 2142 6016 2462 7040
rect 2142 5952 2150 6016
rect 2214 5952 2230 6016
rect 2294 5952 2310 6016
rect 2374 5952 2390 6016
rect 2454 5952 2462 6016
rect 2142 4928 2462 5952
rect 2142 4864 2150 4928
rect 2214 4864 2230 4928
rect 2294 4864 2310 4928
rect 2374 4864 2390 4928
rect 2454 4864 2462 4928
rect 2142 3840 2462 4864
rect 2142 3776 2150 3840
rect 2214 3776 2230 3840
rect 2294 3776 2310 3840
rect 2374 3776 2390 3840
rect 2454 3776 2462 3840
rect 2142 2752 2462 3776
rect 2142 2688 2150 2752
rect 2214 2688 2230 2752
rect 2294 2688 2310 2752
rect 2374 2688 2390 2752
rect 2454 2688 2462 2752
rect 2142 2128 2462 2688
rect 3274 14176 3594 14736
rect 3274 14112 3282 14176
rect 3346 14112 3362 14176
rect 3426 14112 3442 14176
rect 3506 14112 3522 14176
rect 3586 14112 3594 14176
rect 3274 13088 3594 14112
rect 3274 13024 3282 13088
rect 3346 13024 3362 13088
rect 3426 13024 3442 13088
rect 3506 13024 3522 13088
rect 3586 13024 3594 13088
rect 3274 12000 3594 13024
rect 3274 11936 3282 12000
rect 3346 11936 3362 12000
rect 3426 11936 3442 12000
rect 3506 11936 3522 12000
rect 3586 11936 3594 12000
rect 3274 10912 3594 11936
rect 3274 10848 3282 10912
rect 3346 10848 3362 10912
rect 3426 10848 3442 10912
rect 3506 10848 3522 10912
rect 3586 10848 3594 10912
rect 3274 9824 3594 10848
rect 3274 9760 3282 9824
rect 3346 9760 3362 9824
rect 3426 9760 3442 9824
rect 3506 9760 3522 9824
rect 3586 9760 3594 9824
rect 3274 8736 3594 9760
rect 3274 8672 3282 8736
rect 3346 8672 3362 8736
rect 3426 8672 3442 8736
rect 3506 8672 3522 8736
rect 3586 8672 3594 8736
rect 3274 7648 3594 8672
rect 3274 7584 3282 7648
rect 3346 7584 3362 7648
rect 3426 7584 3442 7648
rect 3506 7584 3522 7648
rect 3586 7584 3594 7648
rect 3274 6560 3594 7584
rect 3274 6496 3282 6560
rect 3346 6496 3362 6560
rect 3426 6496 3442 6560
rect 3506 6496 3522 6560
rect 3586 6496 3594 6560
rect 3274 5472 3594 6496
rect 3274 5408 3282 5472
rect 3346 5408 3362 5472
rect 3426 5408 3442 5472
rect 3506 5408 3522 5472
rect 3586 5408 3594 5472
rect 3274 4384 3594 5408
rect 3274 4320 3282 4384
rect 3346 4320 3362 4384
rect 3426 4320 3442 4384
rect 3506 4320 3522 4384
rect 3586 4320 3594 4384
rect 3274 3296 3594 4320
rect 3274 3232 3282 3296
rect 3346 3232 3362 3296
rect 3426 3232 3442 3296
rect 3506 3232 3522 3296
rect 3586 3232 3594 3296
rect 3274 2208 3594 3232
rect 3274 2144 3282 2208
rect 3346 2144 3362 2208
rect 3426 2144 3442 2208
rect 3506 2144 3522 2208
rect 3586 2144 3594 2208
rect 3274 2128 3594 2144
rect 4406 14720 4726 14736
rect 4406 14656 4414 14720
rect 4478 14656 4494 14720
rect 4558 14656 4574 14720
rect 4638 14656 4654 14720
rect 4718 14656 4726 14720
rect 4406 13632 4726 14656
rect 4406 13568 4414 13632
rect 4478 13568 4494 13632
rect 4558 13568 4574 13632
rect 4638 13568 4654 13632
rect 4718 13568 4726 13632
rect 4406 12544 4726 13568
rect 4406 12480 4414 12544
rect 4478 12480 4494 12544
rect 4558 12480 4574 12544
rect 4638 12480 4654 12544
rect 4718 12480 4726 12544
rect 4406 11456 4726 12480
rect 4406 11392 4414 11456
rect 4478 11392 4494 11456
rect 4558 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4726 11456
rect 4406 10368 4726 11392
rect 4406 10304 4414 10368
rect 4478 10304 4494 10368
rect 4558 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4726 10368
rect 4406 9280 4726 10304
rect 4406 9216 4414 9280
rect 4478 9216 4494 9280
rect 4558 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4726 9280
rect 4406 8192 4726 9216
rect 4406 8128 4414 8192
rect 4478 8128 4494 8192
rect 4558 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4726 8192
rect 4406 7104 4726 8128
rect 4406 7040 4414 7104
rect 4478 7040 4494 7104
rect 4558 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4726 7104
rect 4406 6016 4726 7040
rect 4406 5952 4414 6016
rect 4478 5952 4494 6016
rect 4558 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4726 6016
rect 4406 4928 4726 5952
rect 4406 4864 4414 4928
rect 4478 4864 4494 4928
rect 4558 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4726 4928
rect 4406 3840 4726 4864
rect 4406 3776 4414 3840
rect 4478 3776 4494 3840
rect 4558 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4726 3840
rect 4406 2752 4726 3776
rect 4406 2688 4414 2752
rect 4478 2688 4494 2752
rect 4558 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4726 2752
rect 4406 2128 4726 2688
rect 5538 14176 5858 14736
rect 5538 14112 5546 14176
rect 5610 14112 5626 14176
rect 5690 14112 5706 14176
rect 5770 14112 5786 14176
rect 5850 14112 5858 14176
rect 5538 13088 5858 14112
rect 5538 13024 5546 13088
rect 5610 13024 5626 13088
rect 5690 13024 5706 13088
rect 5770 13024 5786 13088
rect 5850 13024 5858 13088
rect 5538 12000 5858 13024
rect 5538 11936 5546 12000
rect 5610 11936 5626 12000
rect 5690 11936 5706 12000
rect 5770 11936 5786 12000
rect 5850 11936 5858 12000
rect 5538 10912 5858 11936
rect 5538 10848 5546 10912
rect 5610 10848 5626 10912
rect 5690 10848 5706 10912
rect 5770 10848 5786 10912
rect 5850 10848 5858 10912
rect 5538 9824 5858 10848
rect 5538 9760 5546 9824
rect 5610 9760 5626 9824
rect 5690 9760 5706 9824
rect 5770 9760 5786 9824
rect 5850 9760 5858 9824
rect 5538 8736 5858 9760
rect 5538 8672 5546 8736
rect 5610 8672 5626 8736
rect 5690 8672 5706 8736
rect 5770 8672 5786 8736
rect 5850 8672 5858 8736
rect 5538 7648 5858 8672
rect 5538 7584 5546 7648
rect 5610 7584 5626 7648
rect 5690 7584 5706 7648
rect 5770 7584 5786 7648
rect 5850 7584 5858 7648
rect 5538 6560 5858 7584
rect 5538 6496 5546 6560
rect 5610 6496 5626 6560
rect 5690 6496 5706 6560
rect 5770 6496 5786 6560
rect 5850 6496 5858 6560
rect 5538 5472 5858 6496
rect 5538 5408 5546 5472
rect 5610 5408 5626 5472
rect 5690 5408 5706 5472
rect 5770 5408 5786 5472
rect 5850 5408 5858 5472
rect 5538 4384 5858 5408
rect 5538 4320 5546 4384
rect 5610 4320 5626 4384
rect 5690 4320 5706 4384
rect 5770 4320 5786 4384
rect 5850 4320 5858 4384
rect 5538 3296 5858 4320
rect 5538 3232 5546 3296
rect 5610 3232 5626 3296
rect 5690 3232 5706 3296
rect 5770 3232 5786 3296
rect 5850 3232 5858 3296
rect 5538 2208 5858 3232
rect 5538 2144 5546 2208
rect 5610 2144 5626 2208
rect 5690 2144 5706 2208
rect 5770 2144 5786 2208
rect 5850 2144 5858 2208
rect 5538 2128 5858 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 38 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 38 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 314 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 1418 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 314 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 1418 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2890 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2522 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 2982 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 2522 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 4086 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 3626 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1605641404
transform 1 0 5742 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1605641404
transform 1 0 5650 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5190 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1605641404
transform 1 0 5834 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4730 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5466 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1605641404
transform 1 0 5742 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 6754 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 6754 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6386 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 38 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 314 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 1418 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1605641404
transform 1 0 2890 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 2522 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 2982 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 4086 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 5190 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 6754 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1605641404
transform 1 0 6294 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 38 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 314 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1605641404
transform 1 0 1418 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1602 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_33
timestamp 1605641404
transform 1 0 3074 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_45
timestamp 1605641404
transform 1 0 4178 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1605641404
transform 1 0 5650 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1605641404
transform 1 0 5282 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1605641404
transform 1 0 5742 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 6754 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 38 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 314 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 1418 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 2890 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 2522 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 2982 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4546 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1605641404
transform 1 0 4086 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_48
timestamp 1605641404
transform 1 0 4454 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp 1605641404
transform 1 0 5742 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 6754 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 38 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 314 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 1418 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 2522 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 3626 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 5650 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 4730 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 5466 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1605641404
transform 1 0 5742 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 6754 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 38 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 38 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 314 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 1418 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 314 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 1418 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 2890 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 2522 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 2982 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_27
timestamp 1605641404
transform 1 0 2522 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_33
timestamp 1605641404
transform 1 0 3074 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3166 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_44
timestamp 1605641404
transform 1 0 4086 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1605641404
transform 1 0 3994 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5098 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 5650 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_52
timestamp 1605641404
transform 1 0 4822 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1605641404
transform 1 0 5374 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_55
timestamp 1605641404
transform 1 0 5098 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1605641404
transform 1 0 5742 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 6754 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 6754 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 38 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 314 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 1418 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 2890 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 2522 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 2982 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1605641404
transform 1 0 4086 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1605641404
transform 1 0 5190 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 6754 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1605641404
transform 1 0 6294 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 38 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 314 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 1418 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1605641404
transform 1 0 2522 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1605641404
transform 1 0 3626 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 5650 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1605641404
transform 1 0 4730 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 5466 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1605641404
transform 1 0 5742 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 6754 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 38 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 314 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1605641404
transform 1 0 1418 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 2890 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1605641404
transform 1 0 2522 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1605641404
transform 1 0 2982 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 4546 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_10_44
timestamp 1605641404
transform 1 0 4086 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1605641404
transform 1 0 4454 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_62
timestamp 1605641404
transform 1 0 5742 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 6754 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 38 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 314 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1605641404
transform 1 0 1418 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1605641404
transform 1 0 2522 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1605641404
transform 1 0 3626 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 5650 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1605641404
transform 1 0 4730 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 5466 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1605641404
transform 1 0 5742 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 6754 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 38 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 314 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 1418 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 2890 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 2522 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 2982 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1605641404
transform 1 0 4086 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5374 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1605641404
transform 1 0 5190 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_62
timestamp 1605641404
transform 1 0 5742 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 6754 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 38 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 38 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 314 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 1418 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 314 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 1418 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 2890 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1605641404
transform 1 0 2522 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 2522 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1605641404
transform 1 0 2982 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1605641404
transform 1 0 3626 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1605641404
transform 1 0 4086 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 5650 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1605641404
transform 1 0 4730 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 5466 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1605641404
transform 1 0 5742 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1605641404
transform 1 0 5190 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 6754 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 6754 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1605641404
transform 1 0 6294 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 38 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 314 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 1418 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1605641404
transform 1 0 2522 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1605641404
transform 1 0 3626 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 5650 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1605641404
transform 1 0 4730 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 5466 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1605641404
transform 1 0 5742 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 6754 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 38 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 314 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 1418 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 2890 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 2522 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1605641404
transform 1 0 2982 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1605641404
transform 1 0 4086 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1605641404
transform 1 0 5190 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 6754 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1605641404
transform 1 0 6294 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 38 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 314 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 1418 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1605641404
transform 1 0 2522 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1605641404
transform 1 0 3626 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 5650 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1605641404
transform 1 0 4730 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 5466 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1605641404
transform 1 0 5742 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 6754 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 38 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 314 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 1418 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 2890 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 2522 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1605641404
transform 1 0 2982 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1605641404
transform 1 0 4086 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1605641404
transform 1 0 5190 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 6754 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1605641404
transform 1 0 6294 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 38 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 38 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 314 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 1418 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 314 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 1418 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 2890 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 2522 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 2522 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 2982 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 3626 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 4086 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 5650 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 4730 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 5466 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1605641404
transform 1 0 5742 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 5190 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 6754 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 6754 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1605641404
transform 1 0 6294 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 38 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 314 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 1418 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1605641404
transform 1 0 2522 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1605641404
transform 1 0 3626 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 5650 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1605641404
transform 1 0 4730 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 5466 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1605641404
transform 1 0 5742 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 6754 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 38 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 314 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 1418 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 2890 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 2522 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 2982 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 4086 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 5742 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1605641404
transform 1 0 5190 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_63
timestamp 1605641404
transform 1 0 5834 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 6754 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1605641404
transform 1 0 6386 0 -1 14688
box -38 -48 130 592
<< labels >>
rlabel metal2 s 1160 16520 1216 17000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 2264 0 2320 480 6 ccff_head
port 1 nsew default input
rlabel metal2 s 4564 0 4620 480 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 7454 14696 7934 14816 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 3 nsew default tristate
rlabel metal2 s 6772 0 6828 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 4 nsew default input
rlabel metal2 s 5668 16520 5724 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 5 nsew default tristate
rlabel metal2 s 56 0 112 480 6 prog_clk
port 6 nsew default input
rlabel metal3 s 7454 6264 7934 6384 6 right_width_0_height_0__pin_0_
port 7 nsew default input
rlabel metal3 s 7454 2048 7934 2168 6 right_width_0_height_0__pin_1_lower
port 8 nsew default tristate
rlabel metal3 s 7454 10480 7934 10600 6 right_width_0_height_0__pin_1_upper
port 9 nsew default tristate
rlabel metal4 s 1010 2128 1330 14736 6 VPWR
port 10 nsew default input
rlabel metal4 s 2142 2128 2462 14736 6 VGND
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 7934 17000
<< end >>
