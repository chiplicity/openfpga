magic
tech sky130A
magscale 1 2
timestamp 1608134292
<< obsli1 >>
rect 1104 2159 15824 17425
<< obsm1 >>
rect 198 1912 16822 17456
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3882 19200 3938 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5170 19200 5226 20000
rect 5538 19200 5594 20000
rect 5998 19200 6054 20000
rect 6366 19200 6422 20000
rect 6826 19200 6882 20000
rect 7194 19200 7250 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8482 19200 8538 20000
rect 8850 19200 8906 20000
rect 9310 19200 9366 20000
rect 9678 19200 9734 20000
rect 10138 19200 10194 20000
rect 10506 19200 10562 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12162 19200 12218 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13450 19200 13506 20000
rect 13818 19200 13874 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 15106 19200 15162 20000
rect 15474 19200 15530 20000
rect 15934 19200 15990 20000
rect 16302 19200 16358 20000
rect 16762 19200 16818 20000
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6550 0 6606 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16762 0 16818 800
<< obsm2 >>
rect 314 19144 514 19200
rect 682 19144 974 19200
rect 1142 19144 1342 19200
rect 1510 19144 1802 19200
rect 1970 19144 2170 19200
rect 2338 19144 2630 19200
rect 2798 19144 2998 19200
rect 3166 19144 3458 19200
rect 3626 19144 3826 19200
rect 3994 19144 4286 19200
rect 4454 19144 4654 19200
rect 4822 19144 5114 19200
rect 5282 19144 5482 19200
rect 5650 19144 5942 19200
rect 6110 19144 6310 19200
rect 6478 19144 6770 19200
rect 6938 19144 7138 19200
rect 7306 19144 7598 19200
rect 7766 19144 7966 19200
rect 8134 19144 8426 19200
rect 8594 19144 8794 19200
rect 8962 19144 9254 19200
rect 9422 19144 9622 19200
rect 9790 19144 10082 19200
rect 10250 19144 10450 19200
rect 10618 19144 10910 19200
rect 11078 19144 11278 19200
rect 11446 19144 11738 19200
rect 11906 19144 12106 19200
rect 12274 19144 12566 19200
rect 12734 19144 12934 19200
rect 13102 19144 13394 19200
rect 13562 19144 13762 19200
rect 13930 19144 14222 19200
rect 14390 19144 14590 19200
rect 14758 19144 15050 19200
rect 15218 19144 15418 19200
rect 15586 19144 15878 19200
rect 16046 19144 16246 19200
rect 16414 19144 16706 19200
rect 204 856 16816 19144
rect 314 800 514 856
rect 682 800 974 856
rect 1142 800 1342 856
rect 1510 800 1802 856
rect 1970 800 2262 856
rect 2430 800 2630 856
rect 2798 800 3090 856
rect 3258 800 3550 856
rect 3718 800 3918 856
rect 4086 800 4378 856
rect 4546 800 4746 856
rect 4914 800 5206 856
rect 5374 800 5666 856
rect 5834 800 6034 856
rect 6202 800 6494 856
rect 6662 800 6954 856
rect 7122 800 7322 856
rect 7490 800 7782 856
rect 7950 800 8150 856
rect 8318 800 8610 856
rect 8778 800 9070 856
rect 9238 800 9438 856
rect 9606 800 9898 856
rect 10066 800 10358 856
rect 10526 800 10726 856
rect 10894 800 11186 856
rect 11354 800 11554 856
rect 11722 800 12014 856
rect 12182 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13302 856
rect 13470 800 13762 856
rect 13930 800 14130 856
rect 14298 800 14590 856
rect 14758 800 14958 856
rect 15126 800 15418 856
rect 15586 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16706 856
<< metal3 >>
rect 0 18232 800 18352
rect 16200 17416 17000 17536
rect 0 14968 800 15088
rect 16200 12384 17000 12504
rect 0 11568 800 11688
rect 0 8304 800 8424
rect 16200 7352 17000 7472
rect 0 4904 800 5024
rect 16200 2456 17000 2576
rect 0 1640 800 1760
<< obsm3 >>
rect 880 18152 16200 18325
rect 800 17616 16200 18152
rect 800 17336 16120 17616
rect 800 15168 16200 17336
rect 880 14888 16200 15168
rect 800 12584 16200 14888
rect 800 12304 16120 12584
rect 800 11768 16200 12304
rect 880 11488 16200 11768
rect 800 8504 16200 11488
rect 880 8224 16200 8504
rect 800 7552 16200 8224
rect 800 7272 16120 7552
rect 800 5104 16200 7272
rect 880 4824 16200 5104
rect 800 2656 16200 4824
rect 800 2376 16120 2656
rect 800 1840 16200 2376
rect 880 1560 16200 1840
rect 800 851 16200 1560
<< metal4 >>
rect 3409 2128 3729 17456
rect 5875 2128 6195 17456
<< obsm4 >>
rect 6275 2128 13590 17456
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 1 nsew default input
rlabel metal3 s 0 18232 800 18352 6 ccff_head
port 2 nsew default input
rlabel metal3 s 16200 12384 17000 12504 6 ccff_tail
port 3 nsew default output
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[0]
port 4 nsew default input
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_in[10]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 800 6 chany_bottom_in[11]
port 6 nsew default input
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_in[12]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_in[13]
port 8 nsew default input
rlabel metal2 s 14646 0 14702 800 6 chany_bottom_in[14]
port 9 nsew default input
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_in[15]
port 10 nsew default input
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_in[16]
port 11 nsew default input
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_in[17]
port 12 nsew default input
rlabel metal2 s 16302 0 16358 800 6 chany_bottom_in[18]
port 13 nsew default input
rlabel metal2 s 16762 0 16818 800 6 chany_bottom_in[19]
port 14 nsew default input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[1]
port 15 nsew default input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[2]
port 16 nsew default input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[3]
port 17 nsew default input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[4]
port 18 nsew default input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[5]
port 19 nsew default input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[6]
port 20 nsew default input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[7]
port 21 nsew default input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[8]
port 22 nsew default input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_in[9]
port 23 nsew default input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 24 nsew default output
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_out[10]
port 25 nsew default output
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[11]
port 26 nsew default output
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_out[12]
port 27 nsew default output
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_out[13]
port 28 nsew default output
rlabel metal2 s 6090 0 6146 800 6 chany_bottom_out[14]
port 29 nsew default output
rlabel metal2 s 6550 0 6606 800 6 chany_bottom_out[15]
port 30 nsew default output
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[16]
port 31 nsew default output
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_out[17]
port 32 nsew default output
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_out[18]
port 33 nsew default output
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_out[19]
port 34 nsew default output
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 35 nsew default output
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 36 nsew default output
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[3]
port 37 nsew default output
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 38 nsew default output
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[5]
port 39 nsew default output
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[6]
port 40 nsew default output
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[7]
port 41 nsew default output
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[8]
port 42 nsew default output
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[9]
port 43 nsew default output
rlabel metal2 s 8850 19200 8906 20000 6 chany_top_in[0]
port 44 nsew default input
rlabel metal2 s 12990 19200 13046 20000 6 chany_top_in[10]
port 45 nsew default input
rlabel metal2 s 13450 19200 13506 20000 6 chany_top_in[11]
port 46 nsew default input
rlabel metal2 s 13818 19200 13874 20000 6 chany_top_in[12]
port 47 nsew default input
rlabel metal2 s 14278 19200 14334 20000 6 chany_top_in[13]
port 48 nsew default input
rlabel metal2 s 14646 19200 14702 20000 6 chany_top_in[14]
port 49 nsew default input
rlabel metal2 s 15106 19200 15162 20000 6 chany_top_in[15]
port 50 nsew default input
rlabel metal2 s 15474 19200 15530 20000 6 chany_top_in[16]
port 51 nsew default input
rlabel metal2 s 15934 19200 15990 20000 6 chany_top_in[17]
port 52 nsew default input
rlabel metal2 s 16302 19200 16358 20000 6 chany_top_in[18]
port 53 nsew default input
rlabel metal2 s 16762 19200 16818 20000 6 chany_top_in[19]
port 54 nsew default input
rlabel metal2 s 9310 19200 9366 20000 6 chany_top_in[1]
port 55 nsew default input
rlabel metal2 s 9678 19200 9734 20000 6 chany_top_in[2]
port 56 nsew default input
rlabel metal2 s 10138 19200 10194 20000 6 chany_top_in[3]
port 57 nsew default input
rlabel metal2 s 10506 19200 10562 20000 6 chany_top_in[4]
port 58 nsew default input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[5]
port 59 nsew default input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[6]
port 60 nsew default input
rlabel metal2 s 11794 19200 11850 20000 6 chany_top_in[7]
port 61 nsew default input
rlabel metal2 s 12162 19200 12218 20000 6 chany_top_in[8]
port 62 nsew default input
rlabel metal2 s 12622 19200 12678 20000 6 chany_top_in[9]
port 63 nsew default input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 64 nsew default output
rlabel metal2 s 4710 19200 4766 20000 6 chany_top_out[10]
port 65 nsew default output
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[11]
port 66 nsew default output
rlabel metal2 s 5538 19200 5594 20000 6 chany_top_out[12]
port 67 nsew default output
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[13]
port 68 nsew default output
rlabel metal2 s 6366 19200 6422 20000 6 chany_top_out[14]
port 69 nsew default output
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_out[15]
port 70 nsew default output
rlabel metal2 s 7194 19200 7250 20000 6 chany_top_out[16]
port 71 nsew default output
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[17]
port 72 nsew default output
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[18]
port 73 nsew default output
rlabel metal2 s 8482 19200 8538 20000 6 chany_top_out[19]
port 74 nsew default output
rlabel metal2 s 1030 19200 1086 20000 6 chany_top_out[1]
port 75 nsew default output
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 76 nsew default output
rlabel metal2 s 1858 19200 1914 20000 6 chany_top_out[3]
port 77 nsew default output
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 78 nsew default output
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[5]
port 79 nsew default output
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 80 nsew default output
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[7]
port 81 nsew default output
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[8]
port 82 nsew default output
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[9]
port 83 nsew default output
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 84 nsew default output
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 85 nsew default input
rlabel metal3 s 0 14968 800 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 86 nsew default output
rlabel metal3 s 0 4904 800 5024 6 left_grid_pin_0_
port 87 nsew default output
rlabel metal3 s 16200 7352 17000 7472 6 prog_clk_0_E_in
port 88 nsew default input
rlabel metal3 s 0 1640 800 1760 6 right_width_0_height_0__pin_0_
port 89 nsew default input
rlabel metal3 s 16200 2456 17000 2576 6 right_width_0_height_0__pin_1_lower
port 90 nsew default output
rlabel metal3 s 16200 17416 17000 17536 6 right_width_0_height_0__pin_1_upper
port 91 nsew default output
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 92 nsew power input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 93 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17000 20000
string LEFview TRUE
<< end >>
