VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_0__1_
  CLASS BLOCK ;
  FOREIGN cby_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 26.560 80.000 27.160 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 44.920 80.000 45.520 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 63.280 80.000 63.880 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 80.960 80.000 81.560 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 99.320 80.000 99.920 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 117.680 80.000 118.280 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 136.040 80.000 136.640 ;
    END
  END address[6]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 197.600 2.210 200.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 197.600 6.350 200.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 197.600 10.950 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 197.600 15.550 200.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 197.600 19.690 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 197.600 24.290 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 197.600 28.890 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 197.600 33.030 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 197.600 37.630 200.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 197.600 42.230 200.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 197.600 46.370 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 197.600 50.970 200.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 197.600 55.570 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 197.600 59.710 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 197.600 64.310 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 197.600 68.910 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 197.600 73.050 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 197.600 77.650 200.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 153.720 80.000 154.320 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 8.880 80.000 9.480 ;
    END
  END enable
  PIN left_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END left_grid_pin_0_
  PIN left_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END left_grid_pin_10_
  PIN left_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 2.400 162.480 ;
    END
  END left_grid_pin_12_
  PIN left_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 2.400 187.640 ;
    END
  END left_grid_pin_14_
  PIN left_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END left_grid_pin_2_
  PIN left_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END left_grid_pin_4_
  PIN left_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.400 87.680 ;
    END
  END left_grid_pin_6_
  PIN left_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END left_grid_pin_8_
  PIN right_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 172.080 80.000 172.680 ;
    END
  END right_grid_pin_3_
  PIN right_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 190.440 80.000 191.040 ;
    END
  END right_grid_pin_7_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 5.520 2.760 74.060 187.920 ;
      LAYER met2 ;
        RECT 2.490 197.320 5.790 197.610 ;
        RECT 6.630 197.320 10.390 197.610 ;
        RECT 11.230 197.320 14.990 197.610 ;
        RECT 15.830 197.320 19.130 197.610 ;
        RECT 19.970 197.320 23.730 197.610 ;
        RECT 24.570 197.320 28.330 197.610 ;
        RECT 29.170 197.320 32.470 197.610 ;
        RECT 33.310 197.320 37.070 197.610 ;
        RECT 37.910 197.320 41.670 197.610 ;
        RECT 42.510 197.320 45.810 197.610 ;
        RECT 46.650 197.320 50.410 197.610 ;
        RECT 51.250 197.320 55.010 197.610 ;
        RECT 55.850 197.320 59.150 197.610 ;
        RECT 59.990 197.320 63.750 197.610 ;
        RECT 64.590 197.320 68.350 197.610 ;
        RECT 69.190 197.320 72.490 197.610 ;
        RECT 73.330 197.320 77.090 197.610 ;
        RECT 1.930 2.680 77.650 197.320 ;
        RECT 2.490 2.400 5.790 2.680 ;
        RECT 6.630 2.400 10.390 2.680 ;
        RECT 11.230 2.400 14.990 2.680 ;
        RECT 15.830 2.400 19.130 2.680 ;
        RECT 19.970 2.400 23.730 2.680 ;
        RECT 24.570 2.400 28.330 2.680 ;
        RECT 29.170 2.400 32.470 2.680 ;
        RECT 33.310 2.400 37.070 2.680 ;
        RECT 37.910 2.400 41.670 2.680 ;
        RECT 42.510 2.400 45.810 2.680 ;
        RECT 46.650 2.400 50.410 2.680 ;
        RECT 51.250 2.400 55.010 2.680 ;
        RECT 55.850 2.400 59.150 2.680 ;
        RECT 59.990 2.400 63.750 2.680 ;
        RECT 64.590 2.400 68.350 2.680 ;
        RECT 69.190 2.400 72.490 2.680 ;
        RECT 73.330 2.400 77.090 2.680 ;
      LAYER met3 ;
        RECT 1.905 190.040 77.200 190.905 ;
        RECT 1.905 188.040 77.675 190.040 ;
        RECT 2.800 186.640 77.675 188.040 ;
        RECT 1.905 173.080 77.675 186.640 ;
        RECT 1.905 171.680 77.200 173.080 ;
        RECT 1.905 162.880 77.675 171.680 ;
        RECT 2.800 161.480 77.675 162.880 ;
        RECT 1.905 154.720 77.675 161.480 ;
        RECT 1.905 153.320 77.200 154.720 ;
        RECT 1.905 137.720 77.675 153.320 ;
        RECT 2.800 137.040 77.675 137.720 ;
        RECT 2.800 136.320 77.200 137.040 ;
        RECT 1.905 135.640 77.200 136.320 ;
        RECT 1.905 118.680 77.675 135.640 ;
        RECT 1.905 117.280 77.200 118.680 ;
        RECT 1.905 113.240 77.675 117.280 ;
        RECT 2.800 111.840 77.675 113.240 ;
        RECT 1.905 100.320 77.675 111.840 ;
        RECT 1.905 98.920 77.200 100.320 ;
        RECT 1.905 88.080 77.675 98.920 ;
        RECT 2.800 86.680 77.675 88.080 ;
        RECT 1.905 81.960 77.675 86.680 ;
        RECT 1.905 80.560 77.200 81.960 ;
        RECT 1.905 64.280 77.675 80.560 ;
        RECT 1.905 62.920 77.200 64.280 ;
        RECT 2.800 62.880 77.200 62.920 ;
        RECT 2.800 61.520 77.675 62.880 ;
        RECT 1.905 45.920 77.675 61.520 ;
        RECT 1.905 44.520 77.200 45.920 ;
        RECT 1.905 37.760 77.675 44.520 ;
        RECT 2.800 36.360 77.675 37.760 ;
        RECT 1.905 27.560 77.675 36.360 ;
        RECT 1.905 26.160 77.200 27.560 ;
        RECT 1.905 13.280 77.675 26.160 ;
        RECT 2.800 11.880 77.675 13.280 ;
        RECT 1.905 9.880 77.675 11.880 ;
        RECT 1.905 9.015 77.200 9.880 ;
      LAYER met4 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_0__1_
END LIBRARY

