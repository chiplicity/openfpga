magic
tech EFS8A
magscale 1 2
timestamp 1604337330
<< locali >>
rect 7941 24599 7975 24701
rect 3985 15895 4019 16133
<< viali >>
rect 2421 25449 2455 25483
rect 1961 25381 1995 25415
rect 8677 25381 8711 25415
rect 9597 25381 9631 25415
rect 10333 25381 10367 25415
rect 1777 25313 1811 25347
rect 8769 25313 8803 25347
rect 2053 25245 2087 25279
rect 8585 25245 8619 25279
rect 10241 25245 10275 25279
rect 10425 25245 10459 25279
rect 12633 25245 12667 25279
rect 1501 25177 1535 25211
rect 2881 25177 2915 25211
rect 8217 25177 8251 25211
rect 3157 25109 3191 25143
rect 9229 25109 9263 25143
rect 9873 25109 9907 25143
rect 2237 24905 2271 24939
rect 10241 24905 10275 24939
rect 9873 24837 9907 24871
rect 3433 24769 3467 24803
rect 10793 24769 10827 24803
rect 12265 24769 12299 24803
rect 13553 24769 13587 24803
rect 7757 24701 7791 24735
rect 7941 24701 7975 24735
rect 8125 24701 8159 24735
rect 8659 24701 8693 24735
rect 11897 24701 11931 24735
rect 12615 24701 12649 24735
rect 14105 24701 14139 24735
rect 14841 24701 14875 24735
rect 15393 24701 15427 24735
rect 15945 24701 15979 24735
rect 2789 24633 2823 24667
rect 3065 24633 3099 24667
rect 7481 24633 7515 24667
rect 8953 24633 8987 24667
rect 9229 24633 9263 24667
rect 10517 24633 10551 24667
rect 10701 24633 10735 24667
rect 12909 24633 12943 24667
rect 13185 24633 13219 24667
rect 14381 24633 14415 24667
rect 1593 24565 1627 24599
rect 2503 24565 2537 24599
rect 2973 24565 3007 24599
rect 3893 24565 3927 24599
rect 5457 24565 5491 24599
rect 7941 24565 7975 24599
rect 9137 24565 9171 24599
rect 11161 24565 11195 24599
rect 13093 24565 13127 24599
rect 15577 24565 15611 24599
rect 1685 24361 1719 24395
rect 8217 24361 8251 24395
rect 8585 24361 8619 24395
rect 9413 24361 9447 24395
rect 10149 24361 10183 24395
rect 10609 24361 10643 24395
rect 12707 24361 12741 24395
rect 16773 24361 16807 24395
rect 24317 24361 24351 24395
rect 2973 24293 3007 24327
rect 11621 24293 11655 24327
rect 13185 24293 13219 24327
rect 21916 24293 21950 24327
rect 2495 24225 2529 24259
rect 5825 24225 5859 24259
rect 6092 24225 6126 24259
rect 13001 24225 13035 24259
rect 15301 24225 15335 24259
rect 15577 24225 15611 24259
rect 16589 24225 16623 24259
rect 24133 24225 24167 24259
rect 2881 24157 2915 24191
rect 3065 24157 3099 24191
rect 4629 24157 4663 24191
rect 11529 24157 11563 24191
rect 11713 24157 11747 24191
rect 13277 24157 13311 24191
rect 21649 24157 21683 24191
rect 3801 24089 3835 24123
rect 11161 24089 11195 24123
rect 12081 24089 12115 24123
rect 23029 24089 23063 24123
rect 2329 24021 2363 24055
rect 3433 24021 3467 24055
rect 4261 24021 4295 24055
rect 5273 24021 5307 24055
rect 7205 24021 7239 24055
rect 9137 24021 9171 24055
rect 12541 24021 12575 24055
rect 13645 24021 13679 24055
rect 23949 24021 23983 24055
rect 2053 23817 2087 23851
rect 3893 23817 3927 23851
rect 10609 23817 10643 23851
rect 11253 23817 11287 23851
rect 11897 23817 11931 23851
rect 14473 23817 14507 23851
rect 16589 23817 16623 23851
rect 21741 23817 21775 23851
rect 24133 23817 24167 23851
rect 25237 23817 25271 23851
rect 5273 23749 5307 23783
rect 6929 23749 6963 23783
rect 17049 23749 17083 23783
rect 1409 23681 1443 23715
rect 5825 23681 5859 23715
rect 7389 23681 7423 23715
rect 8585 23681 8619 23715
rect 11529 23681 11563 23715
rect 22017 23681 22051 23715
rect 2513 23613 2547 23647
rect 5089 23613 5123 23647
rect 5549 23613 5583 23647
rect 7481 23613 7515 23647
rect 7849 23613 7883 23647
rect 9137 23613 9171 23647
rect 9229 23613 9263 23647
rect 13093 23613 13127 23647
rect 15577 23613 15611 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 23949 23613 23983 23647
rect 25053 23613 25087 23647
rect 25605 23613 25639 23647
rect 2780 23545 2814 23579
rect 6193 23545 6227 23579
rect 9474 23545 9508 23579
rect 13360 23545 13394 23579
rect 15853 23545 15887 23579
rect 24501 23545 24535 23579
rect 2329 23477 2363 23511
rect 4721 23477 4755 23511
rect 5733 23477 5767 23511
rect 6653 23477 6687 23511
rect 7389 23477 7423 23511
rect 8217 23477 8251 23511
rect 13001 23477 13035 23511
rect 15301 23477 15335 23511
rect 3709 23273 3743 23307
rect 6101 23273 6135 23307
rect 11069 23273 11103 23307
rect 12081 23273 12115 23307
rect 16773 23273 16807 23307
rect 17877 23273 17911 23307
rect 19073 23273 19107 23307
rect 1676 23205 1710 23239
rect 6377 23205 6411 23239
rect 9956 23205 9990 23239
rect 15577 23205 15611 23239
rect 22661 23205 22695 23239
rect 23949 23205 23983 23239
rect 4077 23137 4111 23171
rect 4344 23137 4378 23171
rect 6817 23137 6851 23171
rect 9689 23137 9723 23171
rect 12440 23137 12474 23171
rect 15301 23137 15335 23171
rect 16589 23137 16623 23171
rect 17693 23137 17727 23171
rect 18889 23137 18923 23171
rect 22385 23137 22419 23171
rect 23673 23137 23707 23171
rect 1409 23069 1443 23103
rect 6561 23069 6595 23103
rect 12173 23069 12207 23103
rect 16037 23069 16071 23103
rect 2789 22933 2823 22967
rect 3433 22933 3467 22967
rect 5457 22933 5491 22967
rect 7941 22933 7975 22967
rect 9321 22933 9355 22967
rect 13553 22933 13587 22967
rect 3341 22729 3375 22763
rect 3617 22729 3651 22763
rect 4537 22729 4571 22763
rect 5273 22729 5307 22763
rect 6561 22729 6595 22763
rect 6929 22729 6963 22763
rect 8861 22729 8895 22763
rect 9229 22729 9263 22763
rect 13369 22729 13403 22763
rect 15853 22729 15887 22763
rect 16957 22729 16991 22763
rect 18245 22729 18279 22763
rect 19349 22729 19383 22763
rect 2053 22661 2087 22695
rect 7849 22661 7883 22695
rect 2513 22593 2547 22627
rect 3065 22593 3099 22627
rect 4169 22593 4203 22627
rect 5089 22593 5123 22627
rect 5825 22593 5859 22627
rect 9321 22593 9355 22627
rect 22569 22593 22603 22627
rect 5549 22525 5583 22559
rect 7205 22525 7239 22559
rect 7481 22525 7515 22559
rect 8217 22525 8251 22559
rect 9588 22525 9622 22559
rect 11253 22525 11287 22559
rect 13921 22525 13955 22559
rect 14177 22525 14211 22559
rect 16405 22525 16439 22559
rect 18061 22525 18095 22559
rect 18613 22525 18647 22559
rect 19165 22525 19199 22559
rect 19717 22525 19751 22559
rect 22293 22525 22327 22559
rect 23029 22525 23063 22559
rect 2605 22457 2639 22491
rect 3893 22457 3927 22491
rect 4077 22457 4111 22491
rect 6285 22457 6319 22491
rect 7389 22457 7423 22491
rect 12265 22457 12299 22491
rect 13829 22457 13863 22491
rect 17693 22457 17727 22491
rect 1593 22389 1627 22423
rect 2513 22389 2547 22423
rect 5733 22389 5767 22423
rect 10701 22389 10735 22423
rect 12725 22389 12759 22423
rect 12909 22389 12943 22423
rect 15301 22389 15335 22423
rect 16221 22389 16255 22423
rect 16589 22389 16623 22423
rect 18981 22389 19015 22423
rect 22109 22389 22143 22423
rect 23857 22389 23891 22423
rect 1409 22185 1443 22219
rect 2329 22185 2363 22219
rect 2973 22185 3007 22219
rect 4353 22185 4387 22219
rect 7389 22185 7423 22219
rect 9413 22185 9447 22219
rect 10241 22185 10275 22219
rect 5825 22117 5859 22151
rect 7205 22117 7239 22151
rect 8401 22117 8435 22151
rect 12541 22117 12575 22151
rect 14105 22117 14139 22151
rect 15761 22117 15795 22151
rect 3065 22049 3099 22083
rect 4813 22049 4847 22083
rect 5917 22049 5951 22083
rect 6285 22049 6319 22083
rect 7481 22049 7515 22083
rect 12633 22049 12667 22083
rect 13461 22049 13495 22083
rect 14197 22049 14231 22083
rect 15485 22049 15519 22083
rect 16773 22049 16807 22083
rect 17049 22049 17083 22083
rect 18061 22049 18095 22083
rect 18337 22049 18371 22083
rect 19349 22049 19383 22083
rect 2973 21981 3007 22015
rect 5825 21981 5859 22015
rect 10149 21981 10183 22015
rect 10333 21981 10367 22015
rect 12449 21981 12483 22015
rect 14013 21981 14047 22015
rect 2513 21913 2547 21947
rect 3801 21913 3835 21947
rect 5365 21913 5399 21947
rect 6929 21913 6963 21947
rect 9781 21913 9815 21947
rect 12081 21913 12115 21947
rect 13093 21913 13127 21947
rect 13645 21913 13679 21947
rect 19533 21913 19567 21947
rect 1869 21845 1903 21879
rect 3433 21845 3467 21879
rect 5181 21845 5215 21879
rect 6745 21845 6779 21879
rect 7849 21845 7883 21879
rect 8953 21845 8987 21879
rect 10701 21845 10735 21879
rect 14657 21845 14691 21879
rect 2145 21641 2179 21675
rect 3985 21641 4019 21675
rect 4905 21641 4939 21675
rect 6101 21641 6135 21675
rect 6653 21641 6687 21675
rect 7849 21641 7883 21675
rect 9505 21641 9539 21675
rect 11713 21641 11747 21675
rect 12541 21641 12575 21675
rect 15485 21641 15519 21675
rect 19533 21641 19567 21675
rect 20637 21641 20671 21675
rect 4629 21573 4663 21607
rect 5181 21573 5215 21607
rect 6929 21573 6963 21607
rect 8493 21573 8527 21607
rect 10057 21573 10091 21607
rect 11345 21573 11379 21607
rect 14105 21573 14139 21607
rect 19901 21573 19935 21607
rect 5549 21505 5583 21539
rect 7481 21505 7515 21539
rect 9045 21505 9079 21539
rect 10609 21505 10643 21539
rect 13093 21505 13127 21539
rect 14657 21505 14691 21539
rect 16221 21505 16255 21539
rect 16681 21505 16715 21539
rect 18337 21505 18371 21539
rect 2605 21437 2639 21471
rect 5733 21437 5767 21471
rect 7205 21437 7239 21471
rect 12817 21437 12851 21471
rect 16405 21437 16439 21471
rect 17141 21437 17175 21471
rect 18061 21437 18095 21471
rect 18797 21437 18831 21471
rect 19349 21437 19383 21471
rect 20453 21437 20487 21471
rect 21005 21437 21039 21471
rect 2421 21369 2455 21403
rect 2872 21369 2906 21403
rect 5641 21369 5675 21403
rect 7389 21369 7423 21403
rect 8309 21369 8343 21403
rect 8769 21369 8803 21403
rect 10333 21369 10367 21403
rect 10517 21369 10551 21403
rect 13001 21369 13035 21403
rect 14381 21369 14415 21403
rect 1593 21301 1627 21335
rect 8953 21301 8987 21335
rect 9781 21301 9815 21335
rect 11989 21301 12023 21335
rect 13553 21301 13587 21335
rect 14565 21301 14599 21335
rect 15117 21301 15151 21335
rect 17785 21301 17819 21335
rect 19257 21301 19291 21335
rect 2881 21097 2915 21131
rect 4629 21097 4663 21131
rect 5181 21097 5215 21131
rect 5549 21097 5583 21131
rect 7113 21097 7147 21131
rect 7665 21097 7699 21131
rect 8493 21097 8527 21131
rect 9413 21097 9447 21131
rect 9965 21097 9999 21131
rect 10333 21097 10367 21131
rect 12541 21097 12575 21131
rect 12909 21097 12943 21131
rect 13645 21097 13679 21131
rect 15025 21097 15059 21131
rect 15945 21097 15979 21131
rect 21097 21097 21131 21131
rect 1768 21029 1802 21063
rect 4445 21029 4479 21063
rect 5978 21029 6012 21063
rect 10762 21029 10796 21063
rect 13461 21029 13495 21063
rect 17509 21029 17543 21063
rect 18797 21029 18831 21063
rect 3525 20961 3559 20995
rect 3893 20961 3927 20995
rect 4721 20961 4755 20995
rect 10517 20961 10551 20995
rect 15761 20961 15795 20995
rect 16865 20961 16899 20995
rect 17601 20961 17635 20995
rect 18521 20961 18555 20995
rect 20913 20961 20947 20995
rect 1501 20893 1535 20927
rect 5733 20893 5767 20927
rect 13737 20893 13771 20927
rect 16037 20893 16071 20927
rect 17417 20893 17451 20927
rect 4169 20825 4203 20859
rect 15485 20825 15519 20859
rect 8953 20757 8987 20791
rect 11897 20757 11931 20791
rect 13185 20757 13219 20791
rect 14105 20757 14139 20791
rect 14565 20757 14599 20791
rect 17049 20757 17083 20791
rect 18153 20757 18187 20791
rect 1685 20553 1719 20587
rect 1961 20553 1995 20587
rect 3801 20553 3835 20587
rect 5641 20553 5675 20587
rect 10701 20553 10735 20587
rect 11253 20553 11287 20587
rect 11897 20553 11931 20587
rect 14381 20553 14415 20587
rect 16497 20553 16531 20587
rect 17509 20553 17543 20587
rect 19073 20553 19107 20587
rect 3433 20485 3467 20519
rect 12173 20485 12207 20519
rect 18153 20485 18187 20519
rect 2513 20417 2547 20451
rect 9229 20417 9263 20451
rect 9321 20417 9355 20451
rect 18705 20417 18739 20451
rect 19809 20417 19843 20451
rect 21097 20417 21131 20451
rect 21649 20417 21683 20451
rect 2237 20349 2271 20383
rect 2881 20349 2915 20383
rect 4169 20349 4203 20383
rect 4261 20349 4295 20383
rect 6837 20349 6871 20383
rect 7104 20349 7138 20383
rect 12449 20349 12483 20383
rect 15025 20349 15059 20383
rect 15117 20349 15151 20383
rect 19625 20349 19659 20383
rect 20361 20349 20395 20383
rect 20913 20349 20947 20383
rect 2421 20281 2455 20315
rect 4506 20281 4540 20315
rect 6285 20281 6319 20315
rect 6653 20281 6687 20315
rect 9566 20281 9600 20315
rect 12694 20281 12728 20315
rect 15362 20281 15396 20315
rect 18429 20281 18463 20315
rect 8217 20213 8251 20247
rect 13829 20213 13863 20247
rect 17049 20213 17083 20247
rect 17785 20213 17819 20247
rect 18613 20213 18647 20247
rect 20729 20213 20763 20247
rect 2605 20009 2639 20043
rect 3157 20009 3191 20043
rect 3525 20009 3559 20043
rect 3801 20009 3835 20043
rect 4251 20009 4285 20043
rect 6285 20009 6319 20043
rect 6929 20009 6963 20043
rect 8033 20009 8067 20043
rect 9413 20009 9447 20043
rect 10701 20009 10735 20043
rect 12541 20009 12575 20043
rect 14105 20009 14139 20043
rect 15025 20009 15059 20043
rect 17601 20009 17635 20043
rect 18521 20009 18555 20043
rect 21281 20009 21315 20043
rect 22477 20009 22511 20043
rect 2697 19941 2731 19975
rect 4537 19941 4571 19975
rect 4721 19941 4755 19975
rect 5549 19941 5583 19975
rect 7205 19941 7239 19975
rect 11713 19941 11747 19975
rect 12992 19941 13026 19975
rect 15945 19941 15979 19975
rect 16466 19941 16500 19975
rect 18153 19941 18187 19975
rect 19349 19941 19383 19975
rect 2421 19873 2455 19907
rect 6101 19873 6135 19907
rect 8493 19873 8527 19907
rect 11529 19873 11563 19907
rect 19073 19873 19107 19907
rect 21097 19873 21131 19907
rect 22293 19873 22327 19907
rect 4813 19805 4847 19839
rect 6377 19805 6411 19839
rect 7941 19805 7975 19839
rect 8125 19805 8159 19839
rect 10149 19805 10183 19839
rect 11805 19805 11839 19839
rect 12725 19805 12759 19839
rect 16221 19805 16255 19839
rect 2145 19737 2179 19771
rect 5825 19737 5859 19771
rect 7573 19737 7607 19771
rect 11253 19737 11287 19771
rect 1685 19669 1719 19703
rect 5181 19669 5215 19703
rect 14657 19669 14691 19703
rect 15485 19669 15519 19703
rect 4077 19465 4111 19499
rect 6009 19465 6043 19499
rect 7573 19465 7607 19499
rect 9597 19465 9631 19499
rect 10517 19465 10551 19499
rect 11713 19465 11747 19499
rect 15393 19465 15427 19499
rect 21373 19465 21407 19499
rect 5549 19397 5583 19431
rect 6653 19397 6687 19431
rect 2053 19329 2087 19363
rect 5089 19329 5123 19363
rect 12817 19329 12851 19363
rect 16957 19329 16991 19363
rect 2320 19261 2354 19295
rect 4611 19261 4645 19295
rect 8217 19261 8251 19295
rect 10149 19261 10183 19295
rect 11069 19261 11103 19295
rect 11345 19261 11379 19295
rect 13001 19261 13035 19295
rect 13553 19261 13587 19295
rect 13921 19261 13955 19295
rect 14013 19261 14047 19295
rect 16589 19261 16623 19295
rect 18061 19261 18095 19295
rect 18317 19261 18351 19295
rect 19993 19261 20027 19295
rect 20637 19261 20671 19295
rect 20913 19261 20947 19295
rect 21925 19261 21959 19295
rect 22477 19261 22511 19295
rect 5181 19193 5215 19227
rect 6837 19193 6871 19227
rect 8462 19193 8496 19227
rect 11253 19193 11287 19227
rect 14258 19193 14292 19227
rect 16313 19193 16347 19227
rect 17877 19193 17911 19227
rect 1869 19125 1903 19159
rect 3433 19125 3467 19159
rect 4353 19125 4387 19159
rect 5089 19125 5123 19159
rect 8125 19125 8159 19159
rect 10783 19125 10817 19159
rect 12173 19125 12207 19159
rect 19441 19125 19475 19159
rect 20453 19125 20487 19159
rect 22109 19125 22143 19159
rect 22845 19125 22879 19159
rect 2605 18921 2639 18955
rect 5733 18921 5767 18955
rect 8309 18921 8343 18955
rect 10793 18921 10827 18955
rect 11621 18921 11655 18955
rect 19165 18921 19199 18955
rect 22937 18921 22971 18955
rect 2421 18853 2455 18887
rect 4620 18853 4654 18887
rect 7389 18853 7423 18887
rect 10241 18853 10275 18887
rect 11253 18853 11287 18887
rect 12357 18853 12391 18887
rect 13277 18853 13311 18887
rect 13921 18853 13955 18887
rect 15853 18853 15887 18887
rect 18052 18853 18086 18887
rect 21189 18853 21223 18887
rect 1685 18785 1719 18819
rect 4353 18785 4387 18819
rect 7205 18785 7239 18819
rect 8585 18785 8619 18819
rect 10057 18785 10091 18819
rect 12173 18785 12207 18819
rect 13737 18785 13771 18819
rect 15669 18785 15703 18819
rect 17785 18785 17819 18819
rect 20913 18785 20947 18819
rect 22753 18785 22787 18819
rect 2697 18717 2731 18751
rect 7481 18717 7515 18751
rect 10333 18717 10367 18751
rect 12449 18717 12483 18751
rect 14013 18717 14047 18751
rect 14381 18717 14415 18751
rect 15945 18717 15979 18751
rect 2145 18649 2179 18683
rect 6929 18649 6963 18683
rect 9781 18649 9815 18683
rect 11897 18649 11931 18683
rect 15393 18649 15427 18683
rect 16681 18649 16715 18683
rect 3157 18581 3191 18615
rect 3433 18581 3467 18615
rect 3801 18581 3835 18615
rect 6285 18581 6319 18615
rect 6745 18581 6779 18615
rect 7941 18581 7975 18615
rect 9413 18581 9447 18615
rect 13461 18581 13495 18615
rect 16313 18581 16347 18615
rect 4537 18377 4571 18411
rect 5549 18377 5583 18411
rect 6285 18377 6319 18411
rect 9045 18377 9079 18411
rect 12265 18377 12299 18411
rect 13185 18377 13219 18411
rect 13553 18377 13587 18411
rect 15025 18377 15059 18411
rect 15945 18377 15979 18411
rect 16221 18377 16255 18411
rect 17785 18377 17819 18411
rect 18337 18377 18371 18411
rect 20913 18377 20947 18411
rect 1501 18309 1535 18343
rect 2053 18241 2087 18275
rect 2513 18241 2547 18275
rect 5641 18241 5675 18275
rect 12633 18241 12667 18275
rect 13645 18241 13679 18275
rect 21557 18241 21591 18275
rect 3065 18173 3099 18207
rect 3157 18173 3191 18207
rect 6837 18173 6871 18207
rect 9505 18173 9539 18207
rect 21281 18173 21315 18207
rect 22017 18173 22051 18207
rect 1777 18105 1811 18139
rect 3424 18105 3458 18139
rect 7082 18105 7116 18139
rect 9772 18105 9806 18139
rect 13912 18105 13946 18139
rect 16497 18105 16531 18139
rect 16681 18105 16715 18139
rect 16773 18105 16807 18139
rect 17141 18105 17175 18139
rect 1961 18037 1995 18071
rect 5089 18037 5123 18071
rect 6561 18037 6595 18071
rect 8217 18037 8251 18071
rect 9413 18037 9447 18071
rect 10885 18037 10919 18071
rect 11437 18037 11471 18071
rect 11805 18037 11839 18071
rect 15577 18037 15611 18071
rect 22753 18037 22787 18071
rect 3341 17833 3375 17867
rect 4813 17833 4847 17867
rect 5273 17833 5307 17867
rect 6745 17833 6779 17867
rect 7389 17833 7423 17867
rect 7665 17833 7699 17867
rect 8401 17833 8435 17867
rect 9505 17833 9539 17867
rect 11069 17833 11103 17867
rect 11897 17833 11931 17867
rect 15117 17833 15151 17867
rect 16681 17833 16715 17867
rect 4353 17765 4387 17799
rect 5610 17765 5644 17799
rect 15546 17765 15580 17799
rect 22017 17765 22051 17799
rect 1409 17697 1443 17731
rect 1676 17697 1710 17731
rect 3709 17697 3743 17731
rect 4077 17697 4111 17731
rect 8493 17697 8527 17731
rect 9689 17697 9723 17731
rect 9956 17697 9990 17731
rect 12429 17697 12463 17731
rect 15301 17697 15335 17731
rect 21741 17697 21775 17731
rect 5365 17629 5399 17663
rect 8309 17629 8343 17663
rect 12173 17629 12207 17663
rect 17785 17629 17819 17663
rect 2789 17561 2823 17595
rect 7941 17561 7975 17595
rect 8861 17561 8895 17595
rect 13553 17493 13587 17527
rect 14105 17493 14139 17527
rect 18337 17493 18371 17527
rect 3249 17289 3283 17323
rect 5733 17289 5767 17323
rect 6469 17289 6503 17323
rect 7021 17289 7055 17323
rect 11161 17289 11195 17323
rect 11529 17289 11563 17323
rect 14657 17289 14691 17323
rect 15025 17289 15059 17323
rect 15393 17289 15427 17323
rect 17785 17289 17819 17323
rect 21741 17289 21775 17323
rect 1869 17221 1903 17255
rect 4445 17221 4479 17255
rect 10149 17221 10183 17255
rect 18153 17221 18187 17255
rect 2421 17153 2455 17187
rect 3341 17153 3375 17187
rect 10701 17153 10735 17187
rect 15485 17153 15519 17187
rect 18521 17153 18555 17187
rect 1685 17085 1719 17119
rect 2881 17085 2915 17119
rect 4997 17085 5031 17119
rect 7389 17085 7423 17119
rect 7573 17085 7607 17119
rect 9505 17085 9539 17119
rect 11805 17085 11839 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 12716 17085 12750 17119
rect 15752 17085 15786 17119
rect 2145 17017 2179 17051
rect 2329 17017 2363 17051
rect 4721 17017 4755 17051
rect 4905 17017 4939 17051
rect 6101 17017 6135 17051
rect 7818 17017 7852 17051
rect 10425 17017 10459 17051
rect 10609 17017 10643 17051
rect 18705 17017 18739 17051
rect 3893 16949 3927 16983
rect 4261 16949 4295 16983
rect 5365 16949 5399 16983
rect 8953 16949 8987 16983
rect 9873 16949 9907 16983
rect 13829 16949 13863 16983
rect 16865 16949 16899 16983
rect 17417 16949 17451 16983
rect 18613 16949 18647 16983
rect 2881 16745 2915 16779
rect 3801 16745 3835 16779
rect 7205 16745 7239 16779
rect 7573 16745 7607 16779
rect 8023 16745 8057 16779
rect 10057 16745 10091 16779
rect 10875 16745 10909 16779
rect 12541 16745 12575 16779
rect 14013 16745 14047 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 17969 16745 18003 16779
rect 4353 16677 4387 16711
rect 8493 16677 8527 16711
rect 11345 16677 11379 16711
rect 11437 16677 11471 16711
rect 12878 16677 12912 16711
rect 1768 16609 1802 16643
rect 3433 16609 3467 16643
rect 5264 16609 5298 16643
rect 8585 16609 8619 16643
rect 9505 16609 9539 16643
rect 10425 16609 10459 16643
rect 11161 16609 11195 16643
rect 12633 16609 12667 16643
rect 16589 16609 16623 16643
rect 16856 16609 16890 16643
rect 1501 16541 1535 16575
rect 4997 16541 5031 16575
rect 8401 16541 8435 16575
rect 4721 16405 4755 16439
rect 6377 16405 6411 16439
rect 2237 16201 2271 16235
rect 7757 16201 7791 16235
rect 8401 16201 8435 16235
rect 8677 16201 8711 16235
rect 9597 16201 9631 16235
rect 11621 16201 11655 16235
rect 12265 16201 12299 16235
rect 13001 16201 13035 16235
rect 16037 16201 16071 16235
rect 16957 16201 16991 16235
rect 2789 16133 2823 16167
rect 3985 16133 4019 16167
rect 6193 16133 6227 16167
rect 3801 16065 3835 16099
rect 1409 15997 1443 16031
rect 1685 15929 1719 15963
rect 2605 15929 2639 15963
rect 3065 15929 3099 15963
rect 3341 15929 3375 15963
rect 9413 16065 9447 16099
rect 10057 16065 10091 16099
rect 10885 16065 10919 16099
rect 11069 16065 11103 16099
rect 13093 16065 13127 16099
rect 15485 16065 15519 16099
rect 16589 16065 16623 16099
rect 17325 16065 17359 16099
rect 4261 15997 4295 16031
rect 4528 15997 4562 16031
rect 4169 15929 4203 15963
rect 6561 15929 6595 15963
rect 10149 15929 10183 15963
rect 13338 15929 13372 15963
rect 16313 15929 16347 15963
rect 16497 15929 16531 15963
rect 3249 15861 3283 15895
rect 3985 15861 4019 15895
rect 5641 15861 5675 15895
rect 6837 15861 6871 15895
rect 7849 15861 7883 15895
rect 10057 15861 10091 15895
rect 14473 15861 14507 15895
rect 15761 15861 15795 15895
rect 3249 15657 3283 15691
rect 5549 15657 5583 15691
rect 8125 15657 8159 15691
rect 11253 15657 11287 15691
rect 12633 15657 12667 15691
rect 13185 15657 13219 15691
rect 16037 15657 16071 15691
rect 2697 15589 2731 15623
rect 4629 15589 4663 15623
rect 5908 15589 5942 15623
rect 10241 15589 10275 15623
rect 10793 15589 10827 15623
rect 1685 15521 1719 15555
rect 5181 15521 5215 15555
rect 5641 15521 5675 15555
rect 9137 15521 9171 15555
rect 10333 15521 10367 15555
rect 2053 15453 2087 15487
rect 2697 15453 2731 15487
rect 2789 15453 2823 15487
rect 4629 15453 4663 15487
rect 4721 15453 4755 15487
rect 10149 15453 10183 15487
rect 7021 15385 7055 15419
rect 9781 15385 9815 15419
rect 2237 15317 2271 15351
rect 3893 15317 3927 15351
rect 4169 15317 4203 15351
rect 9505 15317 9539 15351
rect 4169 15113 4203 15147
rect 5273 15113 5307 15147
rect 6561 15113 6595 15147
rect 8677 15113 8711 15147
rect 9689 15045 9723 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 4721 14977 4755 15011
rect 5825 14977 5859 15011
rect 2412 14909 2446 14943
rect 5089 14909 5123 14943
rect 7297 14909 7331 14943
rect 9781 14909 9815 14943
rect 10048 14909 10082 14943
rect 5549 14841 5583 14875
rect 5733 14841 5767 14875
rect 7542 14841 7576 14875
rect 3525 14773 3559 14807
rect 6285 14773 6319 14807
rect 7113 14773 7147 14807
rect 9229 14773 9263 14807
rect 11161 14773 11195 14807
rect 2789 14569 2823 14603
rect 3341 14569 3375 14603
rect 3709 14569 3743 14603
rect 4629 14569 4663 14603
rect 5733 14569 5767 14603
rect 7021 14569 7055 14603
rect 9137 14569 9171 14603
rect 9505 14569 9539 14603
rect 4445 14501 4479 14535
rect 6469 14501 6503 14535
rect 7849 14501 7883 14535
rect 8033 14501 8067 14535
rect 1409 14433 1443 14467
rect 1676 14433 1710 14467
rect 5273 14433 5307 14467
rect 6285 14433 6319 14467
rect 10221 14433 10255 14467
rect 4721 14365 4755 14399
rect 6561 14365 6595 14399
rect 8125 14365 8159 14399
rect 9965 14365 9999 14399
rect 4169 14297 4203 14331
rect 7573 14297 7607 14331
rect 8493 14297 8527 14331
rect 6009 14229 6043 14263
rect 7389 14229 7423 14263
rect 11345 14229 11379 14263
rect 4629 14025 4663 14059
rect 5641 14025 5675 14059
rect 6377 14025 6411 14059
rect 9045 14025 9079 14059
rect 9689 14025 9723 14059
rect 1501 13957 1535 13991
rect 3065 13957 3099 13991
rect 3985 13957 4019 13991
rect 7205 13957 7239 13991
rect 10333 13957 10367 13991
rect 2053 13889 2087 13923
rect 3617 13889 3651 13923
rect 5181 13889 5215 13923
rect 7573 13889 7607 13923
rect 2513 13821 2547 13855
rect 6009 13821 6043 13855
rect 7665 13821 7699 13855
rect 7932 13821 7966 13855
rect 10149 13821 10183 13855
rect 10701 13821 10735 13855
rect 1777 13753 1811 13787
rect 3341 13753 3375 13787
rect 3525 13753 3559 13787
rect 4905 13753 4939 13787
rect 1961 13685 1995 13719
rect 2881 13685 2915 13719
rect 4445 13685 4479 13719
rect 5089 13685 5123 13719
rect 10057 13685 10091 13719
rect 11253 13685 11287 13719
rect 2513 13481 2547 13515
rect 3525 13481 3559 13515
rect 3893 13481 3927 13515
rect 6009 13481 6043 13515
rect 6837 13481 6871 13515
rect 8585 13481 8619 13515
rect 11069 13481 11103 13515
rect 1961 13413 1995 13447
rect 4261 13413 4295 13447
rect 4896 13413 4930 13447
rect 7665 13413 7699 13447
rect 8861 13413 8895 13447
rect 1777 13345 1811 13379
rect 2973 13345 3007 13379
rect 7481 13345 7515 13379
rect 9956 13345 9990 13379
rect 2053 13277 2087 13311
rect 4629 13277 4663 13311
rect 7757 13277 7791 13311
rect 9689 13277 9723 13311
rect 1501 13209 1535 13243
rect 7205 13209 7239 13243
rect 2881 13141 2915 13175
rect 8125 13141 8159 13175
rect 2421 12937 2455 12971
rect 3985 12937 4019 12971
rect 5273 12937 5307 12971
rect 6193 12937 6227 12971
rect 10609 12937 10643 12971
rect 9689 12869 9723 12903
rect 11345 12869 11379 12903
rect 3433 12801 3467 12835
rect 4445 12801 4479 12835
rect 2973 12733 3007 12767
rect 5457 12733 5491 12767
rect 6837 12733 6871 12767
rect 11161 12733 11195 12767
rect 11713 12733 11747 12767
rect 2697 12665 2731 12699
rect 4537 12665 4571 12699
rect 5733 12665 5767 12699
rect 7082 12665 7116 12699
rect 9965 12665 9999 12699
rect 10241 12665 10275 12699
rect 10977 12665 11011 12699
rect 1685 12597 1719 12631
rect 2145 12597 2179 12631
rect 2881 12597 2915 12631
rect 3801 12597 3835 12631
rect 4445 12597 4479 12631
rect 4997 12597 5031 12631
rect 6561 12597 6595 12631
rect 8217 12597 8251 12631
rect 9045 12597 9079 12631
rect 9505 12597 9539 12631
rect 10149 12597 10183 12631
rect 1869 12393 1903 12427
rect 2329 12393 2363 12427
rect 3433 12393 3467 12427
rect 3893 12393 3927 12427
rect 4721 12393 4755 12427
rect 6653 12393 6687 12427
rect 7297 12393 7331 12427
rect 8585 12393 8619 12427
rect 11437 12393 11471 12427
rect 2973 12325 3007 12359
rect 5540 12325 5574 12359
rect 4077 12257 4111 12291
rect 5273 12257 5307 12291
rect 8677 12257 8711 12291
rect 10313 12257 10347 12291
rect 1409 12189 1443 12223
rect 2973 12189 3007 12223
rect 3065 12189 3099 12223
rect 8493 12189 8527 12223
rect 10057 12189 10091 12223
rect 2513 12053 2547 12087
rect 4261 12053 4295 12087
rect 5181 12053 5215 12087
rect 7849 12053 7883 12087
rect 8125 12053 8159 12087
rect 9965 12053 9999 12087
rect 1685 11849 1719 11883
rect 4813 11849 4847 11883
rect 6193 11849 6227 11883
rect 7297 11849 7331 11883
rect 4169 11781 4203 11815
rect 6469 11781 6503 11815
rect 11345 11713 11379 11747
rect 2145 11645 2179 11679
rect 2237 11645 2271 11679
rect 5089 11645 5123 11679
rect 7757 11645 7791 11679
rect 10241 11645 10275 11679
rect 10793 11645 10827 11679
rect 2504 11577 2538 11611
rect 5365 11577 5399 11611
rect 8002 11577 8036 11611
rect 3617 11509 3651 11543
rect 4629 11509 4663 11543
rect 5273 11509 5307 11543
rect 5825 11509 5859 11543
rect 7573 11509 7607 11543
rect 9137 11509 9171 11543
rect 9781 11509 9815 11543
rect 10057 11509 10091 11543
rect 10425 11509 10459 11543
rect 2513 11305 2547 11339
rect 3709 11305 3743 11339
rect 6561 11305 6595 11339
rect 7941 11305 7975 11339
rect 8493 11305 8527 11339
rect 8861 11305 8895 11339
rect 11621 11305 11655 11339
rect 12909 11305 12943 11339
rect 1777 11237 1811 11271
rect 4629 11237 4663 11271
rect 2329 11169 2363 11203
rect 2605 11169 2639 11203
rect 3065 11169 3099 11203
rect 5641 11169 5675 11203
rect 6193 11169 6227 11203
rect 8033 11169 8067 11203
rect 10508 11169 10542 11203
rect 12725 11169 12759 11203
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 7941 11101 7975 11135
rect 10241 11101 10275 11135
rect 2053 11033 2087 11067
rect 3341 11033 3375 11067
rect 4169 11033 4203 11067
rect 5273 11033 5307 11067
rect 5825 11033 5859 11067
rect 7021 10965 7055 10999
rect 7481 10965 7515 10999
rect 1685 10761 1719 10795
rect 4169 10761 4203 10795
rect 6653 10761 6687 10795
rect 8953 10761 8987 10795
rect 11805 10761 11839 10795
rect 12909 10761 12943 10795
rect 5273 10693 5307 10727
rect 8401 10693 8435 10727
rect 5733 10625 5767 10659
rect 2145 10557 2179 10591
rect 2412 10557 2446 10591
rect 7021 10557 7055 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 5089 10489 5123 10523
rect 5733 10489 5767 10523
rect 5825 10489 5859 10523
rect 6285 10489 6319 10523
rect 7288 10489 7322 10523
rect 9750 10489 9784 10523
rect 11437 10489 11471 10523
rect 12449 10489 12483 10523
rect 1961 10421 1995 10455
rect 3525 10421 3559 10455
rect 4537 10421 4571 10455
rect 10885 10421 10919 10455
rect 1685 10217 1719 10251
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 4353 10217 4387 10251
rect 5457 10217 5491 10251
rect 7021 10217 7055 10251
rect 9873 10217 9907 10251
rect 11621 10217 11655 10251
rect 2329 10149 2363 10183
rect 2881 10149 2915 10183
rect 7665 10149 7699 10183
rect 7481 10081 7515 10115
rect 10508 10081 10542 10115
rect 2329 10013 2363 10047
rect 2421 10013 2455 10047
rect 4979 10013 5013 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 7757 10013 7791 10047
rect 10241 10013 10275 10047
rect 1869 9877 1903 9911
rect 4813 9877 4847 9911
rect 6009 9877 6043 9911
rect 7205 9877 7239 9911
rect 8217 9877 8251 9911
rect 8585 9877 8619 9911
rect 3157 9673 3191 9707
rect 5273 9673 5307 9707
rect 1777 9605 1811 9639
rect 5549 9605 5583 9639
rect 6285 9605 6319 9639
rect 8585 9605 8619 9639
rect 10333 9605 10367 9639
rect 2789 9537 2823 9571
rect 5733 9537 5767 9571
rect 6653 9537 6687 9571
rect 8953 9537 8987 9571
rect 9137 9537 9171 9571
rect 10885 9537 10919 9571
rect 11253 9537 11287 9571
rect 2053 9469 2087 9503
rect 2329 9469 2363 9503
rect 3249 9469 3283 9503
rect 3516 9469 3550 9503
rect 8033 9469 8067 9503
rect 10149 9469 10183 9503
rect 2237 9401 2271 9435
rect 7297 9401 7331 9435
rect 7481 9401 7515 9435
rect 7573 9401 7607 9435
rect 9045 9401 9079 9435
rect 9781 9401 9815 9435
rect 10609 9401 10643 9435
rect 10793 9401 10827 9435
rect 4629 9333 4663 9367
rect 7011 9333 7045 9367
rect 8401 9333 8435 9367
rect 12449 9333 12483 9367
rect 2145 9129 2179 9163
rect 2513 9129 2547 9163
rect 3341 9129 3375 9163
rect 6653 9129 6687 9163
rect 8125 9129 8159 9163
rect 8493 9129 8527 9163
rect 10241 9129 10275 9163
rect 11069 9129 11103 9163
rect 11805 9129 11839 9163
rect 3617 9061 3651 9095
rect 7481 9061 7515 9095
rect 7665 9061 7699 9095
rect 7757 9061 7791 9095
rect 11897 9061 11931 9095
rect 1409 8993 1443 9027
rect 2697 8993 2731 9027
rect 4629 8993 4663 9027
rect 4896 8993 4930 9027
rect 7021 8993 7055 9027
rect 10333 8993 10367 9027
rect 1685 8925 1719 8959
rect 10241 8925 10275 8959
rect 11805 8925 11839 8959
rect 2881 8789 2915 8823
rect 4537 8789 4571 8823
rect 6009 8789 6043 8823
rect 7205 8789 7239 8823
rect 9505 8789 9539 8823
rect 9781 8789 9815 8823
rect 10701 8789 10735 8823
rect 11345 8789 11379 8823
rect 1961 8585 1995 8619
rect 2329 8585 2363 8619
rect 4721 8585 4755 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9781 8585 9815 8619
rect 11253 8585 11287 8619
rect 11805 8585 11839 8619
rect 1593 8517 1627 8551
rect 3709 8517 3743 8551
rect 6929 8517 6963 8551
rect 7941 8517 7975 8551
rect 9413 8517 9447 8551
rect 12173 8517 12207 8551
rect 4077 8449 4111 8483
rect 4997 8449 5031 8483
rect 7297 8449 7331 8483
rect 1409 8381 1443 8415
rect 2513 8381 2547 8415
rect 3525 8381 3559 8415
rect 4261 8381 4295 8415
rect 5825 8381 5859 8415
rect 6653 8381 6687 8415
rect 8401 8381 8435 8415
rect 8953 8381 8987 8415
rect 9873 8381 9907 8415
rect 5549 8313 5583 8347
rect 5733 8313 5767 8347
rect 6285 8313 6319 8347
rect 7481 8313 7515 8347
rect 10118 8313 10152 8347
rect 2697 8245 2731 8279
rect 3157 8245 3191 8279
rect 4169 8245 4203 8279
rect 5255 8245 5289 8279
rect 7389 8245 7423 8279
rect 2421 8041 2455 8075
rect 3157 8041 3191 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 5917 8041 5951 8075
rect 6929 8041 6963 8075
rect 11069 8041 11103 8075
rect 11621 8041 11655 8075
rect 2881 7973 2915 8007
rect 7757 7973 7791 8007
rect 9137 7973 9171 8007
rect 9956 7973 9990 8007
rect 1685 7905 1719 7939
rect 4537 7905 4571 7939
rect 4804 7905 4838 7939
rect 7573 7905 7607 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 1869 7837 1903 7871
rect 7849 7837 7883 7871
rect 6561 7769 6595 7803
rect 7297 7769 7331 7803
rect 8585 7701 8619 7735
rect 2513 7497 2547 7531
rect 2881 7497 2915 7531
rect 3801 7497 3835 7531
rect 4077 7497 4111 7531
rect 6653 7497 6687 7531
rect 7849 7497 7883 7531
rect 9965 7497 9999 7531
rect 10885 7497 10919 7531
rect 6929 7429 6963 7463
rect 3157 7361 3191 7395
rect 4261 7361 4295 7395
rect 8401 7361 8435 7395
rect 1685 7293 1719 7327
rect 2973 7293 3007 7327
rect 4517 7293 4551 7327
rect 6285 7293 6319 7327
rect 7481 7293 7515 7327
rect 8585 7293 8619 7327
rect 1961 7225 1995 7259
rect 7205 7225 7239 7259
rect 7389 7225 7423 7259
rect 8830 7225 8864 7259
rect 5641 7157 5675 7191
rect 10609 7157 10643 7191
rect 2513 6953 2547 6987
rect 3525 6953 3559 6987
rect 5089 6953 5123 6987
rect 6929 6953 6963 6987
rect 8493 6953 8527 6987
rect 4629 6885 4663 6919
rect 7380 6885 7414 6919
rect 10241 6885 10275 6919
rect 1685 6817 1719 6851
rect 1961 6817 1995 6851
rect 2973 6817 3007 6851
rect 4445 6817 4479 6851
rect 4721 6817 4755 6851
rect 5641 6817 5675 6851
rect 6561 6817 6595 6851
rect 10057 6817 10091 6851
rect 10333 6817 10367 6851
rect 7113 6749 7147 6783
rect 3893 6681 3927 6715
rect 5825 6681 5859 6715
rect 2881 6613 2915 6647
rect 4169 6613 4203 6647
rect 5549 6613 5583 6647
rect 9781 6613 9815 6647
rect 3709 6409 3743 6443
rect 4169 6409 4203 6443
rect 8217 6409 8251 6443
rect 9873 6409 9907 6443
rect 10517 6409 10551 6443
rect 2789 6341 2823 6375
rect 10241 6341 10275 6375
rect 3249 6273 3283 6307
rect 4261 6273 4295 6307
rect 9321 6273 9355 6307
rect 1409 6205 1443 6239
rect 2053 6205 2087 6239
rect 2605 6205 2639 6239
rect 3341 6205 3375 6239
rect 4528 6205 4562 6239
rect 6561 6205 6595 6239
rect 6837 6205 6871 6239
rect 7082 6137 7116 6171
rect 1593 6069 1627 6103
rect 3249 6069 3283 6103
rect 5641 6069 5675 6103
rect 6193 6069 6227 6103
rect 1685 5865 1719 5899
rect 3157 5865 3191 5899
rect 3801 5865 3835 5899
rect 5641 5865 5675 5899
rect 6837 5865 6871 5899
rect 7021 5865 7055 5899
rect 7573 5865 7607 5899
rect 4721 5797 4755 5831
rect 1777 5729 1811 5763
rect 3525 5729 3559 5763
rect 4813 5729 4847 5763
rect 1961 5661 1995 5695
rect 4629 5661 4663 5695
rect 2789 5593 2823 5627
rect 4261 5593 4295 5627
rect 2513 5321 2547 5355
rect 3985 5321 4019 5355
rect 4721 5321 4755 5355
rect 1961 5185 1995 5219
rect 1685 5117 1719 5151
rect 2973 5117 3007 5151
rect 3525 5117 3559 5151
rect 4077 5117 4111 5151
rect 3157 4981 3191 5015
rect 4261 4981 4295 5015
rect 4997 4981 5031 5015
rect 4261 4777 4295 4811
rect 1409 4641 1443 4675
rect 2513 4641 2547 4675
rect 2789 4573 2823 4607
rect 1593 4437 1627 4471
rect 2053 4437 2087 4471
rect 1685 4233 1719 4267
rect 3617 4233 3651 4267
rect 3249 4097 3283 4131
rect 2145 4029 2179 4063
rect 3433 4029 3467 4063
rect 3985 4029 4019 4063
rect 2421 3961 2455 3995
rect 2973 3961 3007 3995
rect 1685 3689 1719 3723
rect 1777 3553 1811 3587
rect 1961 3485 1995 3519
rect 2237 3145 2271 3179
rect 2881 3145 2915 3179
rect 3249 3145 3283 3179
rect 1409 2941 1443 2975
rect 2697 2941 2731 2975
rect 1685 2873 1719 2907
rect 1961 2601 1995 2635
rect 4629 2533 4663 2567
rect 1409 2465 1443 2499
rect 2513 2465 2547 2499
rect 3065 2465 3099 2499
rect 4077 2465 4111 2499
rect 1593 2261 1627 2295
rect 2697 2261 2731 2295
rect 4261 2261 4295 2295
<< metal1 >>
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 7282 26568 7288 26580
rect 4120 26540 7288 26568
rect 4120 26528 4126 26540
rect 7282 26528 7288 26540
rect 7340 26528 7346 26580
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2038 25440 2044 25492
rect 2096 25480 2102 25492
rect 2409 25483 2467 25489
rect 2409 25480 2421 25483
rect 2096 25452 2421 25480
rect 2096 25440 2102 25452
rect 2409 25449 2421 25452
rect 2455 25480 2467 25483
rect 2682 25480 2688 25492
rect 2455 25452 2688 25480
rect 2455 25449 2467 25452
rect 2409 25443 2467 25449
rect 2682 25440 2688 25452
rect 2740 25440 2746 25492
rect 1578 25372 1584 25424
rect 1636 25412 1642 25424
rect 1949 25415 2007 25421
rect 1949 25412 1961 25415
rect 1636 25384 1961 25412
rect 1636 25372 1642 25384
rect 1949 25381 1961 25384
rect 1995 25381 2007 25415
rect 1949 25375 2007 25381
rect 8202 25372 8208 25424
rect 8260 25412 8266 25424
rect 8665 25415 8723 25421
rect 8665 25412 8677 25415
rect 8260 25384 8677 25412
rect 8260 25372 8266 25384
rect 8665 25381 8677 25384
rect 8711 25381 8723 25415
rect 8665 25375 8723 25381
rect 9585 25415 9643 25421
rect 9585 25381 9597 25415
rect 9631 25412 9643 25415
rect 10226 25412 10232 25424
rect 9631 25384 10232 25412
rect 9631 25381 9643 25384
rect 9585 25375 9643 25381
rect 10226 25372 10232 25384
rect 10284 25412 10290 25424
rect 10321 25415 10379 25421
rect 10321 25412 10333 25415
rect 10284 25384 10333 25412
rect 10284 25372 10290 25384
rect 10321 25381 10333 25384
rect 10367 25381 10379 25415
rect 10321 25375 10379 25381
rect 1762 25344 1768 25356
rect 1723 25316 1768 25344
rect 1762 25304 1768 25316
rect 1820 25304 1826 25356
rect 8294 25304 8300 25356
rect 8352 25344 8358 25356
rect 8757 25347 8815 25353
rect 8757 25344 8769 25347
rect 8352 25316 8769 25344
rect 8352 25304 8358 25316
rect 8757 25313 8769 25316
rect 8803 25344 8815 25347
rect 10134 25344 10140 25356
rect 8803 25316 10140 25344
rect 8803 25313 8815 25316
rect 8757 25307 8815 25313
rect 10134 25304 10140 25316
rect 10192 25304 10198 25356
rect 2041 25279 2099 25285
rect 2041 25245 2053 25279
rect 2087 25276 2099 25279
rect 3418 25276 3424 25288
rect 2087 25248 3424 25276
rect 2087 25245 2099 25248
rect 2041 25239 2099 25245
rect 3418 25236 3424 25248
rect 3476 25236 3482 25288
rect 8570 25276 8576 25288
rect 8531 25248 8576 25276
rect 8570 25236 8576 25248
rect 8628 25236 8634 25288
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25245 10287 25279
rect 10410 25276 10416 25288
rect 10371 25248 10416 25276
rect 10229 25239 10287 25245
rect 1489 25211 1547 25217
rect 1489 25177 1501 25211
rect 1535 25208 1547 25211
rect 2774 25208 2780 25220
rect 1535 25180 2780 25208
rect 1535 25177 1547 25180
rect 1489 25171 1547 25177
rect 2774 25168 2780 25180
rect 2832 25168 2838 25220
rect 2869 25211 2927 25217
rect 2869 25177 2881 25211
rect 2915 25208 2927 25211
rect 3050 25208 3056 25220
rect 2915 25180 3056 25208
rect 2915 25177 2927 25180
rect 2869 25171 2927 25177
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 8205 25211 8263 25217
rect 8205 25177 8217 25211
rect 8251 25208 8263 25211
rect 9398 25208 9404 25220
rect 8251 25180 9404 25208
rect 8251 25177 8263 25180
rect 8205 25171 8263 25177
rect 9398 25168 9404 25180
rect 9456 25208 9462 25220
rect 10244 25208 10272 25239
rect 10410 25236 10416 25248
rect 10468 25236 10474 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 12802 25276 12808 25288
rect 12667 25248 12808 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 9456 25180 10272 25208
rect 9456 25168 9462 25180
rect 23658 25168 23664 25220
rect 23716 25208 23722 25220
rect 24302 25208 24308 25220
rect 23716 25180 24308 25208
rect 23716 25168 23722 25180
rect 24302 25168 24308 25180
rect 24360 25168 24366 25220
rect 3142 25140 3148 25152
rect 3103 25112 3148 25140
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 9217 25143 9275 25149
rect 9217 25109 9229 25143
rect 9263 25140 9275 25143
rect 9306 25140 9312 25152
rect 9263 25112 9312 25140
rect 9263 25109 9275 25112
rect 9217 25103 9275 25109
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 9861 25143 9919 25149
rect 9861 25109 9873 25143
rect 9907 25140 9919 25143
rect 15286 25140 15292 25152
rect 9907 25112 15292 25140
rect 9907 25109 9919 25112
rect 9861 25103 9919 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 842 24896 848 24948
rect 900 24936 906 24948
rect 2225 24939 2283 24945
rect 2225 24936 2237 24939
rect 900 24908 2237 24936
rect 900 24896 906 24908
rect 2225 24905 2237 24908
rect 2271 24905 2283 24939
rect 2225 24899 2283 24905
rect 2240 24732 2268 24899
rect 2774 24896 2780 24948
rect 2832 24936 2838 24948
rect 3878 24936 3884 24948
rect 2832 24908 3884 24936
rect 2832 24896 2838 24908
rect 3878 24896 3884 24908
rect 3936 24896 3942 24948
rect 10226 24936 10232 24948
rect 10187 24908 10232 24936
rect 10226 24896 10232 24908
rect 10284 24896 10290 24948
rect 2682 24828 2688 24880
rect 2740 24828 2746 24880
rect 9674 24828 9680 24880
rect 9732 24868 9738 24880
rect 9861 24871 9919 24877
rect 9861 24868 9873 24871
rect 9732 24840 9873 24868
rect 9732 24828 9738 24840
rect 9861 24837 9873 24840
rect 9907 24868 9919 24871
rect 10410 24868 10416 24880
rect 9907 24840 10416 24868
rect 9907 24837 9919 24840
rect 9861 24831 9919 24837
rect 10410 24828 10416 24840
rect 10468 24868 10474 24880
rect 10962 24868 10968 24880
rect 10468 24840 10968 24868
rect 10468 24828 10474 24840
rect 10962 24828 10968 24840
rect 11020 24828 11026 24880
rect 12986 24868 12992 24880
rect 12820 24840 12992 24868
rect 2700 24800 2728 24828
rect 3418 24800 3424 24812
rect 2700 24772 2820 24800
rect 3379 24772 3424 24800
rect 2240 24704 2728 24732
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2491 24599 2549 24605
rect 2491 24565 2503 24599
rect 2537 24596 2549 24599
rect 2590 24596 2596 24608
rect 2537 24568 2596 24596
rect 2537 24565 2549 24568
rect 2491 24559 2549 24565
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 2700 24596 2728 24704
rect 2792 24676 2820 24772
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 5994 24760 6000 24812
rect 6052 24800 6058 24812
rect 6546 24800 6552 24812
rect 6052 24772 6552 24800
rect 6052 24760 6058 24772
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 10192 24772 10793 24800
rect 10192 24760 10198 24772
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12820 24800 12848 24840
rect 12986 24828 12992 24840
rect 13044 24828 13050 24880
rect 12299 24772 12848 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 12952 24772 13553 24800
rect 12952 24760 12958 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 6086 24732 6092 24744
rect 3712 24704 6092 24732
rect 2774 24624 2780 24676
rect 2832 24664 2838 24676
rect 3050 24664 3056 24676
rect 2832 24636 2877 24664
rect 3011 24636 3056 24664
rect 2832 24624 2838 24636
rect 3050 24624 3056 24636
rect 3108 24624 3114 24676
rect 2961 24599 3019 24605
rect 2961 24596 2973 24599
rect 2700 24568 2973 24596
rect 2961 24565 2973 24568
rect 3007 24596 3019 24599
rect 3712 24596 3740 24704
rect 6086 24692 6092 24704
rect 6144 24732 6150 24744
rect 7745 24735 7803 24741
rect 7745 24732 7757 24735
rect 6144 24704 7757 24732
rect 6144 24692 6150 24704
rect 7745 24701 7757 24704
rect 7791 24732 7803 24735
rect 7929 24735 7987 24741
rect 7929 24732 7941 24735
rect 7791 24704 7941 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 7929 24701 7941 24704
rect 7975 24701 7987 24735
rect 8110 24732 8116 24744
rect 8071 24704 8116 24732
rect 7929 24695 7987 24701
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 8647 24735 8705 24741
rect 8647 24701 8659 24735
rect 8693 24732 8705 24735
rect 11885 24735 11943 24741
rect 8693 24704 10732 24732
rect 8693 24701 8705 24704
rect 8647 24695 8705 24701
rect 10704 24676 10732 24704
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 12434 24732 12440 24744
rect 11931 24704 12440 24732
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 12434 24692 12440 24704
rect 12492 24692 12498 24744
rect 12603 24735 12661 24741
rect 12603 24701 12615 24735
rect 12649 24732 12661 24735
rect 14093 24735 14151 24741
rect 14093 24732 14105 24735
rect 12649 24704 14105 24732
rect 12649 24701 12661 24704
rect 12603 24695 12661 24701
rect 14093 24701 14105 24704
rect 14139 24732 14151 24735
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 14139 24704 14841 24732
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14829 24701 14841 24704
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24732 15439 24735
rect 15562 24732 15568 24744
rect 15427 24704 15568 24732
rect 15427 24701 15439 24704
rect 15381 24695 15439 24701
rect 15562 24692 15568 24704
rect 15620 24732 15626 24744
rect 15933 24735 15991 24741
rect 15933 24732 15945 24735
rect 15620 24704 15945 24732
rect 15620 24692 15626 24704
rect 15933 24701 15945 24704
rect 15979 24701 15991 24735
rect 15933 24695 15991 24701
rect 7469 24667 7527 24673
rect 7469 24633 7481 24667
rect 7515 24664 7527 24667
rect 8294 24664 8300 24676
rect 7515 24636 8300 24664
rect 7515 24633 7527 24636
rect 7469 24627 7527 24633
rect 8294 24624 8300 24636
rect 8352 24624 8358 24676
rect 8938 24664 8944 24676
rect 8899 24636 8944 24664
rect 8938 24624 8944 24636
rect 8996 24624 9002 24676
rect 9217 24667 9275 24673
rect 9217 24633 9229 24667
rect 9263 24664 9275 24667
rect 9306 24664 9312 24676
rect 9263 24636 9312 24664
rect 9263 24633 9275 24636
rect 9217 24627 9275 24633
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 10042 24624 10048 24676
rect 10100 24664 10106 24676
rect 10505 24667 10563 24673
rect 10505 24664 10517 24667
rect 10100 24636 10517 24664
rect 10100 24624 10106 24636
rect 10505 24633 10517 24636
rect 10551 24633 10563 24667
rect 10686 24664 10692 24676
rect 10599 24636 10692 24664
rect 10505 24627 10563 24633
rect 3878 24596 3884 24608
rect 3007 24568 3740 24596
rect 3839 24568 3884 24596
rect 3007 24565 3019 24568
rect 2961 24559 3019 24565
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 5445 24599 5503 24605
rect 5445 24565 5457 24599
rect 5491 24596 5503 24599
rect 5534 24596 5540 24608
rect 5491 24568 5540 24596
rect 5491 24565 5503 24568
rect 5445 24559 5503 24565
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 7929 24599 7987 24605
rect 7929 24565 7941 24599
rect 7975 24596 7987 24599
rect 9122 24596 9128 24608
rect 7975 24568 9128 24596
rect 7975 24565 7987 24568
rect 7929 24559 7987 24565
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 10520 24596 10548 24627
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 12894 24664 12900 24676
rect 12855 24636 12900 24664
rect 12894 24624 12900 24636
rect 12952 24624 12958 24676
rect 12986 24624 12992 24676
rect 13044 24664 13050 24676
rect 13173 24667 13231 24673
rect 13173 24664 13185 24667
rect 13044 24636 13185 24664
rect 13044 24624 13050 24636
rect 13173 24633 13185 24636
rect 13219 24664 13231 24667
rect 13354 24664 13360 24676
rect 13219 24636 13360 24664
rect 13219 24633 13231 24636
rect 13173 24627 13231 24633
rect 13354 24624 13360 24636
rect 13412 24624 13418 24676
rect 14366 24664 14372 24676
rect 14327 24636 14372 24664
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 16482 24664 16488 24676
rect 15580 24636 16488 24664
rect 11149 24599 11207 24605
rect 11149 24596 11161 24599
rect 10520 24568 11161 24596
rect 11149 24565 11161 24568
rect 11195 24565 11207 24599
rect 11149 24559 11207 24565
rect 13081 24599 13139 24605
rect 13081 24565 13093 24599
rect 13127 24596 13139 24599
rect 13262 24596 13268 24608
rect 13127 24568 13268 24596
rect 13127 24565 13139 24568
rect 13081 24559 13139 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 15580 24605 15608 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 15565 24599 15623 24605
rect 15565 24565 15577 24599
rect 15611 24565 15623 24599
rect 15565 24559 15623 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1673 24395 1731 24401
rect 1673 24361 1685 24395
rect 1719 24392 1731 24395
rect 1762 24392 1768 24404
rect 1719 24364 1768 24392
rect 1719 24361 1731 24364
rect 1673 24355 1731 24361
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 7558 24352 7564 24404
rect 7616 24392 7622 24404
rect 8018 24392 8024 24404
rect 7616 24364 8024 24392
rect 7616 24352 7622 24364
rect 8018 24352 8024 24364
rect 8076 24352 8082 24404
rect 8205 24395 8263 24401
rect 8205 24361 8217 24395
rect 8251 24392 8263 24395
rect 8570 24392 8576 24404
rect 8251 24364 8576 24392
rect 8251 24361 8263 24364
rect 8205 24355 8263 24361
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 9398 24392 9404 24404
rect 9359 24364 9404 24392
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 10134 24392 10140 24404
rect 10095 24364 10140 24392
rect 10134 24352 10140 24364
rect 10192 24352 10198 24404
rect 10597 24395 10655 24401
rect 10597 24361 10609 24395
rect 10643 24392 10655 24395
rect 10686 24392 10692 24404
rect 10643 24364 10692 24392
rect 10643 24361 10655 24364
rect 10597 24355 10655 24361
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 12695 24395 12753 24401
rect 12695 24392 12707 24395
rect 12492 24364 12707 24392
rect 12492 24352 12498 24364
rect 12695 24361 12707 24364
rect 12741 24392 12753 24395
rect 13262 24392 13268 24404
rect 12741 24364 13268 24392
rect 12741 24361 12753 24364
rect 12695 24355 12753 24361
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 16761 24395 16819 24401
rect 16761 24361 16773 24395
rect 16807 24392 16819 24395
rect 17034 24392 17040 24404
rect 16807 24364 17040 24392
rect 16807 24361 16819 24364
rect 16761 24355 16819 24361
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 24305 24395 24363 24401
rect 24305 24361 24317 24395
rect 24351 24392 24363 24395
rect 25406 24392 25412 24404
rect 24351 24364 25412 24392
rect 24351 24361 24363 24364
rect 24305 24355 24363 24361
rect 25406 24352 25412 24364
rect 25464 24352 25470 24404
rect 2866 24284 2872 24336
rect 2924 24324 2930 24336
rect 2961 24327 3019 24333
rect 2961 24324 2973 24327
rect 2924 24296 2973 24324
rect 2924 24284 2930 24296
rect 2961 24293 2973 24296
rect 3007 24293 3019 24327
rect 6178 24324 6184 24336
rect 2961 24287 3019 24293
rect 5828 24296 6184 24324
rect 2498 24265 2504 24268
rect 2483 24259 2504 24265
rect 2483 24225 2495 24259
rect 2483 24219 2504 24225
rect 2498 24216 2504 24219
rect 2556 24216 2562 24268
rect 5828 24265 5856 24296
rect 6178 24284 6184 24296
rect 6236 24284 6242 24336
rect 11606 24324 11612 24336
rect 11567 24296 11612 24324
rect 11606 24284 11612 24296
rect 11664 24284 11670 24336
rect 21910 24333 21916 24336
rect 13173 24327 13231 24333
rect 13173 24324 13185 24327
rect 12084 24296 13185 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24225 5871 24259
rect 5813 24219 5871 24225
rect 6080 24259 6138 24265
rect 6080 24225 6092 24259
rect 6126 24256 6138 24259
rect 6638 24256 6644 24268
rect 6126 24228 6644 24256
rect 6126 24225 6138 24228
rect 6080 24219 6138 24225
rect 6638 24216 6644 24228
rect 6696 24216 6702 24268
rect 2774 24148 2780 24200
rect 2832 24188 2838 24200
rect 2869 24191 2927 24197
rect 2869 24188 2881 24191
rect 2832 24160 2881 24188
rect 2832 24148 2838 24160
rect 2869 24157 2881 24160
rect 2915 24157 2927 24191
rect 3050 24188 3056 24200
rect 2963 24160 3056 24188
rect 2869 24151 2927 24157
rect 3050 24148 3056 24160
rect 3108 24188 3114 24200
rect 3418 24188 3424 24200
rect 3108 24160 3424 24188
rect 3108 24148 3114 24160
rect 3418 24148 3424 24160
rect 3476 24148 3482 24200
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 4304 24160 4629 24188
rect 4304 24148 4310 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 11514 24188 11520 24200
rect 11475 24160 11520 24188
rect 4617 24151 4675 24157
rect 11514 24148 11520 24160
rect 11572 24148 11578 24200
rect 11698 24188 11704 24200
rect 11659 24160 11704 24188
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 2406 24080 2412 24132
rect 2464 24120 2470 24132
rect 3789 24123 3847 24129
rect 3789 24120 3801 24123
rect 2464 24092 3801 24120
rect 2464 24080 2470 24092
rect 3789 24089 3801 24092
rect 3835 24089 3847 24123
rect 3789 24083 3847 24089
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7742 24120 7748 24132
rect 6972 24092 7748 24120
rect 6972 24080 6978 24092
rect 7742 24080 7748 24092
rect 7800 24080 7806 24132
rect 12084 24129 12112 24296
rect 13173 24293 13185 24296
rect 13219 24293 13231 24327
rect 21904 24324 21916 24333
rect 21871 24296 21916 24324
rect 13173 24287 13231 24293
rect 21904 24287 21916 24296
rect 21910 24284 21916 24287
rect 21968 24284 21974 24336
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 12989 24259 13047 24265
rect 12989 24256 13001 24259
rect 12492 24228 13001 24256
rect 12492 24216 12498 24228
rect 12989 24225 13001 24228
rect 13035 24225 13047 24259
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 12989 24219 13047 24225
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 15565 24259 15623 24265
rect 15565 24225 15577 24259
rect 15611 24256 15623 24259
rect 16574 24256 16580 24268
rect 15611 24228 16580 24256
rect 15611 24225 15623 24228
rect 15565 24219 15623 24225
rect 16574 24216 16580 24228
rect 16632 24216 16638 24268
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24121 24259 24179 24265
rect 24121 24256 24133 24259
rect 24084 24228 24133 24256
rect 24084 24216 24090 24228
rect 24121 24225 24133 24228
rect 24167 24225 24179 24259
rect 24121 24219 24179 24225
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24157 13323 24191
rect 21634 24188 21640 24200
rect 21595 24160 21640 24188
rect 13265 24151 13323 24157
rect 11149 24123 11207 24129
rect 11149 24089 11161 24123
rect 11195 24120 11207 24123
rect 12069 24123 12127 24129
rect 12069 24120 12081 24123
rect 11195 24092 12081 24120
rect 11195 24089 11207 24092
rect 11149 24083 11207 24089
rect 12069 24089 12081 24092
rect 12115 24089 12127 24123
rect 12069 24083 12127 24089
rect 2314 24052 2320 24064
rect 2227 24024 2320 24052
rect 2314 24012 2320 24024
rect 2372 24052 2378 24064
rect 2774 24052 2780 24064
rect 2372 24024 2780 24052
rect 2372 24012 2378 24024
rect 2774 24012 2780 24024
rect 2832 24012 2838 24064
rect 3418 24052 3424 24064
rect 3379 24024 3424 24052
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 4249 24055 4307 24061
rect 4249 24052 4261 24055
rect 4212 24024 4261 24052
rect 4212 24012 4218 24024
rect 4249 24021 4261 24024
rect 4295 24021 4307 24055
rect 4249 24015 4307 24021
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5350 24052 5356 24064
rect 5307 24024 5356 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5350 24012 5356 24024
rect 5408 24052 5414 24064
rect 7193 24055 7251 24061
rect 7193 24052 7205 24055
rect 5408 24024 7205 24052
rect 5408 24012 5414 24024
rect 7193 24021 7205 24024
rect 7239 24021 7251 24055
rect 7193 24015 7251 24021
rect 8938 24012 8944 24064
rect 8996 24052 9002 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 8996 24024 9137 24052
rect 8996 24012 9002 24024
rect 9125 24021 9137 24024
rect 9171 24052 9183 24055
rect 9858 24052 9864 24064
rect 9171 24024 9864 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 9858 24012 9864 24024
rect 9916 24012 9922 24064
rect 12529 24055 12587 24061
rect 12529 24021 12541 24055
rect 12575 24052 12587 24055
rect 13280 24052 13308 24151
rect 21634 24148 21640 24160
rect 21692 24148 21698 24200
rect 23014 24120 23020 24132
rect 22975 24092 23020 24120
rect 23014 24080 23020 24092
rect 23072 24080 23078 24132
rect 13446 24052 13452 24064
rect 12575 24024 13452 24052
rect 12575 24021 12587 24024
rect 12529 24015 12587 24021
rect 13446 24012 13452 24024
rect 13504 24052 13510 24064
rect 13633 24055 13691 24061
rect 13633 24052 13645 24055
rect 13504 24024 13645 24052
rect 13504 24012 13510 24024
rect 13633 24021 13645 24024
rect 13679 24021 13691 24055
rect 23934 24052 23940 24064
rect 23895 24024 23940 24052
rect 13633 24015 13691 24021
rect 23934 24012 23940 24024
rect 23992 24012 23998 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2041 23851 2099 23857
rect 2041 23817 2053 23851
rect 2087 23848 2099 23851
rect 2866 23848 2872 23860
rect 2087 23820 2872 23848
rect 2087 23817 2099 23820
rect 2041 23811 2099 23817
rect 2866 23808 2872 23820
rect 2924 23848 2930 23860
rect 2924 23820 3464 23848
rect 2924 23808 2930 23820
rect 3436 23780 3464 23820
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 3881 23851 3939 23857
rect 3881 23848 3893 23851
rect 3568 23820 3893 23848
rect 3568 23808 3574 23820
rect 3881 23817 3893 23820
rect 3927 23817 3939 23851
rect 8846 23848 8852 23860
rect 3881 23811 3939 23817
rect 5184 23820 8852 23848
rect 5184 23780 5212 23820
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10597 23851 10655 23857
rect 10597 23848 10609 23851
rect 10192 23820 10609 23848
rect 10192 23808 10198 23820
rect 10597 23817 10609 23820
rect 10643 23817 10655 23851
rect 10597 23811 10655 23817
rect 11241 23851 11299 23857
rect 11241 23817 11253 23851
rect 11287 23848 11299 23851
rect 11606 23848 11612 23860
rect 11287 23820 11612 23848
rect 11287 23817 11299 23820
rect 11241 23811 11299 23817
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 11698 23808 11704 23860
rect 11756 23848 11762 23860
rect 11885 23851 11943 23857
rect 11885 23848 11897 23851
rect 11756 23820 11897 23848
rect 11756 23808 11762 23820
rect 11885 23817 11897 23820
rect 11931 23817 11943 23851
rect 11885 23811 11943 23817
rect 13354 23808 13360 23860
rect 13412 23848 13418 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 13412 23820 14473 23848
rect 13412 23808 13418 23820
rect 14461 23817 14473 23820
rect 14507 23817 14519 23851
rect 16574 23848 16580 23860
rect 16535 23820 16580 23848
rect 14461 23811 14519 23817
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 21729 23851 21787 23857
rect 21729 23817 21741 23851
rect 21775 23848 21787 23851
rect 21910 23848 21916 23860
rect 21775 23820 21916 23848
rect 21775 23817 21787 23820
rect 21729 23811 21787 23817
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 24118 23848 24124 23860
rect 24079 23820 24124 23848
rect 24118 23808 24124 23820
rect 24176 23808 24182 23860
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 26510 23848 26516 23860
rect 25271 23820 26516 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 26510 23808 26516 23820
rect 26568 23808 26574 23860
rect 3436 23752 5212 23780
rect 5261 23783 5319 23789
rect 5261 23749 5273 23783
rect 5307 23780 5319 23783
rect 5442 23780 5448 23792
rect 5307 23752 5448 23780
rect 5307 23749 5319 23752
rect 5261 23743 5319 23749
rect 5442 23740 5448 23752
rect 5500 23740 5506 23792
rect 6822 23740 6828 23792
rect 6880 23780 6886 23792
rect 6917 23783 6975 23789
rect 6917 23780 6929 23783
rect 6880 23752 6929 23780
rect 6880 23740 6886 23752
rect 6917 23749 6929 23752
rect 6963 23749 6975 23783
rect 6917 23743 6975 23749
rect 15930 23740 15936 23792
rect 15988 23780 15994 23792
rect 17037 23783 17095 23789
rect 17037 23780 17049 23783
rect 15988 23752 17049 23780
rect 15988 23740 15994 23752
rect 17037 23749 17049 23752
rect 17083 23749 17095 23783
rect 17037 23743 17095 23749
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 1762 23712 1768 23724
rect 1443 23684 1768 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 5350 23672 5356 23724
rect 5408 23712 5414 23724
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 5408 23684 5825 23712
rect 5408 23672 5414 23684
rect 5813 23681 5825 23684
rect 5859 23712 5871 23715
rect 6270 23712 6276 23724
rect 5859 23684 6276 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6270 23672 6276 23684
rect 6328 23672 6334 23724
rect 7374 23712 7380 23724
rect 7287 23684 7380 23712
rect 7374 23672 7380 23684
rect 7432 23712 7438 23724
rect 8573 23715 8631 23721
rect 8573 23712 8585 23715
rect 7432 23684 8585 23712
rect 7432 23672 7438 23684
rect 8573 23681 8585 23684
rect 8619 23681 8631 23715
rect 11514 23712 11520 23724
rect 11475 23684 11520 23712
rect 8573 23675 8631 23681
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 22002 23712 22008 23724
rect 21963 23684 22008 23712
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2332 23616 2513 23644
rect 1670 23468 1676 23520
rect 1728 23508 1734 23520
rect 2332 23517 2360 23616
rect 2501 23613 2513 23616
rect 2547 23644 2559 23647
rect 3970 23644 3976 23656
rect 2547 23616 3976 23644
rect 2547 23613 2559 23616
rect 2501 23607 2559 23613
rect 3970 23604 3976 23616
rect 4028 23604 4034 23656
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23644 5135 23647
rect 5534 23644 5540 23656
rect 5123 23616 5540 23644
rect 5123 23613 5135 23616
rect 5077 23607 5135 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 6288 23644 6316 23672
rect 7469 23647 7527 23653
rect 7469 23644 7481 23647
rect 6288 23616 7481 23644
rect 7469 23613 7481 23616
rect 7515 23644 7527 23647
rect 7837 23647 7895 23653
rect 7837 23644 7849 23647
rect 7515 23616 7849 23644
rect 7515 23613 7527 23616
rect 7469 23607 7527 23613
rect 7837 23613 7849 23616
rect 7883 23613 7895 23647
rect 7837 23607 7895 23613
rect 9125 23647 9183 23653
rect 9125 23613 9137 23647
rect 9171 23644 9183 23647
rect 9214 23644 9220 23656
rect 9171 23616 9220 23644
rect 9171 23613 9183 23616
rect 9125 23607 9183 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 13081 23647 13139 23653
rect 13081 23644 13093 23647
rect 13004 23616 13093 23644
rect 2768 23579 2826 23585
rect 2768 23545 2780 23579
rect 2814 23576 2826 23579
rect 3418 23576 3424 23588
rect 2814 23548 3424 23576
rect 2814 23545 2826 23548
rect 2768 23539 2826 23545
rect 3418 23536 3424 23548
rect 3476 23536 3482 23588
rect 3988 23576 4016 23604
rect 6178 23576 6184 23588
rect 3988 23548 6184 23576
rect 6178 23536 6184 23548
rect 6236 23536 6242 23588
rect 9306 23536 9312 23588
rect 9364 23576 9370 23588
rect 9462 23579 9520 23585
rect 9462 23576 9474 23579
rect 9364 23548 9474 23576
rect 9364 23536 9370 23548
rect 9462 23545 9474 23548
rect 9508 23545 9520 23579
rect 9462 23539 9520 23545
rect 13004 23520 13032 23616
rect 13081 23613 13093 23616
rect 13127 23613 13139 23647
rect 13081 23607 13139 23613
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23644 15623 23647
rect 16022 23644 16028 23656
rect 15611 23616 16028 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 16022 23604 16028 23616
rect 16080 23604 16086 23656
rect 16850 23644 16856 23656
rect 16811 23616 16856 23644
rect 16850 23604 16856 23616
rect 16908 23644 16914 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16908 23616 17417 23644
rect 16908 23604 16914 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23934 23644 23940 23656
rect 23532 23616 23940 23644
rect 23532 23604 23538 23616
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 25041 23647 25099 23653
rect 25041 23644 25053 23647
rect 24912 23616 25053 23644
rect 24912 23604 24918 23616
rect 25041 23613 25053 23616
rect 25087 23644 25099 23647
rect 25593 23647 25651 23653
rect 25593 23644 25605 23647
rect 25087 23616 25605 23644
rect 25087 23613 25099 23616
rect 25041 23607 25099 23613
rect 25593 23613 25605 23616
rect 25639 23613 25651 23647
rect 25593 23607 25651 23613
rect 13348 23579 13406 23585
rect 13348 23545 13360 23579
rect 13394 23576 13406 23579
rect 13446 23576 13452 23588
rect 13394 23548 13452 23576
rect 13394 23545 13406 23548
rect 13348 23539 13406 23545
rect 13446 23536 13452 23548
rect 13504 23536 13510 23588
rect 15841 23579 15899 23585
rect 15841 23545 15853 23579
rect 15887 23576 15899 23579
rect 16482 23576 16488 23588
rect 15887 23548 16488 23576
rect 15887 23545 15899 23548
rect 15841 23539 15899 23545
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 23566 23536 23572 23588
rect 23624 23576 23630 23588
rect 24026 23576 24032 23588
rect 23624 23548 24032 23576
rect 23624 23536 23630 23548
rect 24026 23536 24032 23548
rect 24084 23576 24090 23588
rect 24489 23579 24547 23585
rect 24489 23576 24501 23579
rect 24084 23548 24501 23576
rect 24084 23536 24090 23548
rect 24489 23545 24501 23548
rect 24535 23545 24547 23579
rect 24489 23539 24547 23545
rect 2317 23511 2375 23517
rect 2317 23508 2329 23511
rect 1728 23480 2329 23508
rect 1728 23468 1734 23480
rect 2317 23477 2329 23480
rect 2363 23477 2375 23511
rect 2317 23471 2375 23477
rect 4709 23511 4767 23517
rect 4709 23477 4721 23511
rect 4755 23508 4767 23511
rect 5350 23508 5356 23520
rect 4755 23480 5356 23508
rect 4755 23477 4767 23480
rect 4709 23471 4767 23477
rect 5350 23468 5356 23480
rect 5408 23508 5414 23520
rect 5721 23511 5779 23517
rect 5721 23508 5733 23511
rect 5408 23480 5733 23508
rect 5408 23468 5414 23480
rect 5721 23477 5733 23480
rect 5767 23477 5779 23511
rect 6638 23508 6644 23520
rect 6599 23480 6644 23508
rect 5721 23471 5779 23477
rect 6638 23468 6644 23480
rect 6696 23468 6702 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7377 23511 7435 23517
rect 7377 23508 7389 23511
rect 6972 23480 7389 23508
rect 6972 23468 6978 23480
rect 7377 23477 7389 23480
rect 7423 23508 7435 23511
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 7423 23480 8217 23508
rect 7423 23477 7435 23480
rect 7377 23471 7435 23477
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8205 23471 8263 23477
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 12710 23508 12716 23520
rect 11756 23480 12716 23508
rect 11756 23468 11762 23480
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 12986 23508 12992 23520
rect 12947 23480 12992 23508
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 15286 23508 15292 23520
rect 15247 23480 15292 23508
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2406 23264 2412 23316
rect 2464 23304 2470 23316
rect 2590 23304 2596 23316
rect 2464 23276 2596 23304
rect 2464 23264 2470 23276
rect 2590 23264 2596 23276
rect 2648 23304 2654 23316
rect 3697 23307 3755 23313
rect 3697 23304 3709 23307
rect 2648 23276 3709 23304
rect 2648 23264 2654 23276
rect 3697 23273 3709 23276
rect 3743 23273 3755 23307
rect 3697 23267 3755 23273
rect 5994 23264 6000 23316
rect 6052 23304 6058 23316
rect 6089 23307 6147 23313
rect 6089 23304 6101 23307
rect 6052 23276 6101 23304
rect 6052 23264 6058 23276
rect 6089 23273 6101 23276
rect 6135 23304 6147 23307
rect 6822 23304 6828 23316
rect 6135 23276 6828 23304
rect 6135 23273 6147 23276
rect 6089 23267 6147 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12069 23307 12127 23313
rect 12069 23273 12081 23307
rect 12115 23304 12127 23307
rect 12342 23304 12348 23316
rect 12115 23276 12348 23304
rect 12115 23273 12127 23276
rect 12069 23267 12127 23273
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 16761 23307 16819 23313
rect 16761 23273 16773 23307
rect 16807 23304 16819 23307
rect 17586 23304 17592 23316
rect 16807 23276 17592 23304
rect 16807 23273 16819 23276
rect 16761 23267 16819 23273
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 17862 23304 17868 23316
rect 17823 23276 17868 23304
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 19058 23304 19064 23316
rect 19019 23276 19064 23304
rect 19058 23264 19064 23276
rect 19116 23264 19122 23316
rect 1664 23239 1722 23245
rect 1664 23205 1676 23239
rect 1710 23236 1722 23239
rect 3050 23236 3056 23248
rect 1710 23208 3056 23236
rect 1710 23205 1722 23208
rect 1664 23199 1722 23205
rect 3050 23196 3056 23208
rect 3108 23236 3114 23248
rect 3510 23236 3516 23248
rect 3108 23208 3516 23236
rect 3108 23196 3114 23208
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 6270 23196 6276 23248
rect 6328 23236 6334 23248
rect 6365 23239 6423 23245
rect 6365 23236 6377 23239
rect 6328 23208 6377 23236
rect 6328 23196 6334 23208
rect 6365 23205 6377 23208
rect 6411 23205 6423 23239
rect 6365 23199 6423 23205
rect 9944 23239 10002 23245
rect 9944 23205 9956 23239
rect 9990 23236 10002 23239
rect 10134 23236 10140 23248
rect 9990 23208 10140 23236
rect 9990 23205 10002 23208
rect 9944 23199 10002 23205
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 4028 23140 4077 23168
rect 4028 23128 4034 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 4065 23131 4123 23137
rect 4332 23171 4390 23177
rect 4332 23137 4344 23171
rect 4378 23168 4390 23171
rect 5074 23168 5080 23180
rect 4378 23140 5080 23168
rect 4378 23137 4390 23140
rect 4332 23131 4390 23137
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 6380 23168 6408 23199
rect 10134 23196 10140 23208
rect 10192 23196 10198 23248
rect 15562 23236 15568 23248
rect 15523 23208 15568 23236
rect 15562 23196 15568 23208
rect 15620 23196 15626 23248
rect 22649 23239 22707 23245
rect 22649 23205 22661 23239
rect 22695 23236 22707 23239
rect 23474 23236 23480 23248
rect 22695 23208 23480 23236
rect 22695 23205 22707 23208
rect 22649 23199 22707 23205
rect 23474 23196 23480 23208
rect 23532 23196 23538 23248
rect 23937 23239 23995 23245
rect 23937 23205 23949 23239
rect 23983 23236 23995 23239
rect 24762 23236 24768 23248
rect 23983 23208 24768 23236
rect 23983 23205 23995 23208
rect 23937 23199 23995 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 6805 23171 6863 23177
rect 6805 23168 6817 23171
rect 6380 23140 6817 23168
rect 6805 23137 6817 23140
rect 6851 23137 6863 23171
rect 6805 23131 6863 23137
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9272 23140 9689 23168
rect 9272 23128 9278 23140
rect 9677 23137 9689 23140
rect 9723 23168 9735 23171
rect 10962 23168 10968 23180
rect 9723 23140 10968 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 10962 23128 10968 23140
rect 11020 23128 11026 23180
rect 12428 23171 12486 23177
rect 12428 23137 12440 23171
rect 12474 23168 12486 23171
rect 12710 23168 12716 23180
rect 12474 23140 12716 23168
rect 12474 23137 12486 23140
rect 12428 23131 12486 23137
rect 12710 23128 12716 23140
rect 12768 23128 12774 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15378 23168 15384 23180
rect 15335 23140 15384 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 17678 23168 17684 23180
rect 17639 23140 17684 23168
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 18782 23128 18788 23180
rect 18840 23168 18846 23180
rect 18877 23171 18935 23177
rect 18877 23168 18889 23171
rect 18840 23140 18889 23168
rect 18840 23128 18846 23140
rect 18877 23137 18889 23140
rect 18923 23137 18935 23171
rect 18877 23131 18935 23137
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22152 23140 22385 23168
rect 22152 23128 22158 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22373 23131 22431 23137
rect 23661 23171 23719 23177
rect 23661 23137 23673 23171
rect 23707 23168 23719 23171
rect 23750 23168 23756 23180
rect 23707 23140 23756 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23069 1455 23103
rect 1397 23063 1455 23069
rect 1412 22964 1440 23063
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6549 23103 6607 23109
rect 6549 23100 6561 23103
rect 6236 23072 6561 23100
rect 6236 23060 6242 23072
rect 6549 23069 6561 23072
rect 6595 23069 6607 23103
rect 12158 23100 12164 23112
rect 12119 23072 12164 23100
rect 6549 23063 6607 23069
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 16022 23100 16028 23112
rect 15983 23072 16028 23100
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 1578 22964 1584 22976
rect 1412 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 2774 22924 2780 22976
rect 2832 22964 2838 22976
rect 3418 22964 3424 22976
rect 2832 22936 2877 22964
rect 3331 22936 3424 22964
rect 2832 22924 2838 22936
rect 3418 22924 3424 22936
rect 3476 22964 3482 22976
rect 5445 22967 5503 22973
rect 5445 22964 5457 22967
rect 3476 22936 5457 22964
rect 3476 22924 3482 22936
rect 5445 22933 5457 22936
rect 5491 22933 5503 22967
rect 7926 22964 7932 22976
rect 7887 22936 7932 22964
rect 5445 22927 5503 22933
rect 7926 22924 7932 22936
rect 7984 22924 7990 22976
rect 9306 22964 9312 22976
rect 9267 22936 9312 22964
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 13446 22924 13452 22976
rect 13504 22964 13510 22976
rect 13541 22967 13599 22973
rect 13541 22964 13553 22967
rect 13504 22936 13553 22964
rect 13504 22924 13510 22936
rect 13541 22933 13553 22936
rect 13587 22933 13599 22967
rect 13541 22927 13599 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3329 22763 3387 22769
rect 3329 22760 3341 22763
rect 2832 22732 3341 22760
rect 2832 22720 2838 22732
rect 3329 22729 3341 22732
rect 3375 22729 3387 22763
rect 3602 22760 3608 22772
rect 3563 22732 3608 22760
rect 3329 22723 3387 22729
rect 2041 22695 2099 22701
rect 2041 22661 2053 22695
rect 2087 22692 2099 22695
rect 2087 22664 3280 22692
rect 2087 22661 2099 22664
rect 2041 22655 2099 22661
rect 2498 22624 2504 22636
rect 2459 22596 2504 22624
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 3050 22624 3056 22636
rect 2608 22596 3056 22624
rect 2608 22500 2636 22596
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3252 22556 3280 22664
rect 3344 22624 3372 22723
rect 3602 22720 3608 22732
rect 3660 22720 3666 22772
rect 3970 22720 3976 22772
rect 4028 22760 4034 22772
rect 4525 22763 4583 22769
rect 4525 22760 4537 22763
rect 4028 22732 4537 22760
rect 4028 22720 4034 22732
rect 4525 22729 4537 22732
rect 4571 22729 4583 22763
rect 4525 22723 4583 22729
rect 5166 22720 5172 22772
rect 5224 22760 5230 22772
rect 5261 22763 5319 22769
rect 5261 22760 5273 22763
rect 5224 22732 5273 22760
rect 5224 22720 5230 22732
rect 5261 22729 5273 22732
rect 5307 22729 5319 22763
rect 5261 22723 5319 22729
rect 6178 22720 6184 22772
rect 6236 22760 6242 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6236 22732 6561 22760
rect 6236 22720 6242 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 6549 22723 6607 22729
rect 6917 22763 6975 22769
rect 6917 22729 6929 22763
rect 6963 22760 6975 22763
rect 7374 22760 7380 22772
rect 6963 22732 7380 22760
rect 6963 22729 6975 22732
rect 6917 22723 6975 22729
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 8849 22763 8907 22769
rect 8849 22729 8861 22763
rect 8895 22760 8907 22763
rect 9214 22760 9220 22772
rect 8895 22732 9220 22760
rect 8895 22729 8907 22732
rect 8849 22723 8907 22729
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 13354 22760 13360 22772
rect 13315 22732 13360 22760
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 15378 22720 15384 22772
rect 15436 22760 15442 22772
rect 15841 22763 15899 22769
rect 15841 22760 15853 22763
rect 15436 22732 15853 22760
rect 15436 22720 15442 22732
rect 15841 22729 15853 22732
rect 15887 22729 15899 22763
rect 15841 22723 15899 22729
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16945 22763 17003 22769
rect 16945 22760 16957 22763
rect 16632 22732 16957 22760
rect 16632 22720 16638 22732
rect 16945 22729 16957 22732
rect 16991 22729 17003 22763
rect 16945 22723 17003 22729
rect 18233 22763 18291 22769
rect 18233 22729 18245 22763
rect 18279 22760 18291 22763
rect 18690 22760 18696 22772
rect 18279 22732 18696 22760
rect 18279 22729 18291 22732
rect 18233 22723 18291 22729
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 19518 22760 19524 22772
rect 19383 22732 19524 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 19518 22720 19524 22732
rect 19576 22720 19582 22772
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 7837 22695 7895 22701
rect 7837 22692 7849 22695
rect 7156 22664 7849 22692
rect 7156 22652 7162 22664
rect 7837 22661 7849 22664
rect 7883 22692 7895 22695
rect 8202 22692 8208 22704
rect 7883 22664 8208 22692
rect 7883 22661 7895 22664
rect 7837 22655 7895 22661
rect 8202 22652 8208 22664
rect 8260 22652 8266 22704
rect 4157 22627 4215 22633
rect 4157 22624 4169 22627
rect 3344 22596 4169 22624
rect 4157 22593 4169 22596
rect 4203 22593 4215 22627
rect 5074 22624 5080 22636
rect 4987 22596 5080 22624
rect 4157 22587 4215 22593
rect 5074 22584 5080 22596
rect 5132 22624 5138 22636
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5132 22596 5825 22624
rect 5132 22584 5138 22596
rect 5813 22593 5825 22596
rect 5859 22624 5871 22627
rect 7926 22624 7932 22636
rect 5859 22596 7932 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 7926 22584 7932 22596
rect 7984 22584 7990 22636
rect 9232 22624 9260 22720
rect 9309 22627 9367 22633
rect 9309 22624 9321 22627
rect 9232 22596 9321 22624
rect 9309 22593 9321 22596
rect 9355 22593 9367 22627
rect 13372 22624 13400 22720
rect 22557 22627 22615 22633
rect 13372 22596 14044 22624
rect 9309 22587 9367 22593
rect 5534 22556 5540 22568
rect 3252 22528 4108 22556
rect 5495 22528 5540 22556
rect 4080 22500 4108 22528
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 7098 22516 7104 22568
rect 7156 22556 7162 22568
rect 7193 22559 7251 22565
rect 7193 22556 7205 22559
rect 7156 22528 7205 22556
rect 7156 22516 7162 22528
rect 7193 22525 7205 22528
rect 7239 22525 7251 22559
rect 7466 22556 7472 22568
rect 7427 22528 7472 22556
rect 7193 22519 7251 22525
rect 7466 22516 7472 22528
rect 7524 22556 7530 22568
rect 9582 22565 9588 22568
rect 8205 22559 8263 22565
rect 8205 22556 8217 22559
rect 7524 22528 8217 22556
rect 7524 22516 7530 22528
rect 8205 22525 8217 22528
rect 8251 22525 8263 22559
rect 9576 22556 9588 22565
rect 9543 22528 9588 22556
rect 8205 22519 8263 22525
rect 9576 22519 9588 22528
rect 2590 22488 2596 22500
rect 2551 22460 2596 22488
rect 2590 22448 2596 22460
rect 2648 22448 2654 22500
rect 3878 22488 3884 22500
rect 3839 22460 3884 22488
rect 3878 22448 3884 22460
rect 3936 22448 3942 22500
rect 4062 22488 4068 22500
rect 4023 22460 4068 22488
rect 4062 22448 4068 22460
rect 4120 22448 4126 22500
rect 6270 22488 6276 22500
rect 6183 22460 6276 22488
rect 6270 22448 6276 22460
rect 6328 22488 6334 22500
rect 7374 22488 7380 22500
rect 6328 22460 7380 22488
rect 6328 22448 6334 22460
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 2406 22380 2412 22432
rect 2464 22420 2470 22432
rect 2501 22423 2559 22429
rect 2501 22420 2513 22423
rect 2464 22392 2513 22420
rect 2464 22380 2470 22392
rect 2501 22389 2513 22392
rect 2547 22389 2559 22423
rect 2501 22383 2559 22389
rect 5721 22423 5779 22429
rect 5721 22389 5733 22423
rect 5767 22420 5779 22423
rect 5994 22420 6000 22432
rect 5767 22392 6000 22420
rect 5767 22389 5779 22392
rect 5721 22383 5779 22389
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 8220 22420 8248 22519
rect 9582 22516 9588 22519
rect 9640 22516 9646 22568
rect 10134 22516 10140 22568
rect 10192 22556 10198 22568
rect 11241 22559 11299 22565
rect 11241 22556 11253 22559
rect 10192 22528 11253 22556
rect 10192 22516 10198 22528
rect 11241 22525 11253 22528
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 13909 22559 13967 22565
rect 13909 22525 13921 22559
rect 13955 22525 13967 22559
rect 14016 22556 14044 22596
rect 22557 22593 22569 22627
rect 22603 22624 22615 22627
rect 23566 22624 23572 22636
rect 22603 22596 23572 22624
rect 22603 22593 22615 22596
rect 22557 22587 22615 22593
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 14165 22559 14223 22565
rect 14165 22556 14177 22559
rect 14016 22528 14177 22556
rect 13909 22519 13967 22525
rect 14165 22525 14177 22528
rect 14211 22525 14223 22559
rect 16393 22559 16451 22565
rect 16393 22556 16405 22559
rect 14165 22519 14223 22525
rect 16224 22528 16405 22556
rect 10962 22448 10968 22500
rect 11020 22488 11026 22500
rect 12158 22488 12164 22500
rect 11020 22460 12164 22488
rect 11020 22448 11026 22460
rect 12158 22448 12164 22460
rect 12216 22488 12222 22500
rect 12253 22491 12311 22497
rect 12253 22488 12265 22491
rect 12216 22460 12265 22488
rect 12216 22448 12222 22460
rect 12253 22457 12265 22460
rect 12299 22488 12311 22491
rect 12986 22488 12992 22500
rect 12299 22460 12992 22488
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 12986 22448 12992 22460
rect 13044 22488 13050 22500
rect 13817 22491 13875 22497
rect 13817 22488 13829 22491
rect 13044 22460 13829 22488
rect 13044 22448 13050 22460
rect 13817 22457 13829 22460
rect 13863 22488 13875 22491
rect 13924 22488 13952 22519
rect 13863 22460 13952 22488
rect 13863 22457 13875 22460
rect 13817 22451 13875 22457
rect 16224 22432 16252 22528
rect 16393 22525 16405 22528
rect 16439 22525 16451 22559
rect 16393 22519 16451 22525
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18049 22559 18107 22565
rect 18049 22556 18061 22559
rect 17920 22528 18061 22556
rect 17920 22516 17926 22528
rect 18049 22525 18061 22528
rect 18095 22556 18107 22559
rect 18601 22559 18659 22565
rect 18601 22556 18613 22559
rect 18095 22528 18613 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 18601 22525 18613 22528
rect 18647 22525 18659 22559
rect 19150 22556 19156 22568
rect 19063 22528 19156 22556
rect 18601 22519 18659 22525
rect 19150 22516 19156 22528
rect 19208 22556 19214 22568
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 19208 22528 19717 22556
rect 19208 22516 19214 22528
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 22278 22556 22284 22568
rect 22239 22528 22284 22556
rect 19705 22519 19763 22525
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 23017 22559 23075 22565
rect 23017 22556 23029 22559
rect 22336 22528 23029 22556
rect 22336 22516 22342 22528
rect 23017 22525 23029 22528
rect 23063 22525 23075 22559
rect 23017 22519 23075 22525
rect 16666 22448 16672 22500
rect 16724 22488 16730 22500
rect 17678 22488 17684 22500
rect 16724 22460 17684 22488
rect 16724 22448 16730 22460
rect 17678 22448 17684 22460
rect 17736 22448 17742 22500
rect 10689 22423 10747 22429
rect 10689 22420 10701 22423
rect 8220 22392 10701 22420
rect 10689 22389 10701 22392
rect 10735 22389 10747 22423
rect 12710 22420 12716 22432
rect 12671 22392 12716 22420
rect 10689 22383 10747 22389
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 12897 22423 12955 22429
rect 12897 22389 12909 22423
rect 12943 22420 12955 22423
rect 13262 22420 13268 22432
rect 12943 22392 13268 22420
rect 12943 22389 12955 22392
rect 12897 22383 12955 22389
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 13538 22380 13544 22432
rect 13596 22420 13602 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 13596 22392 15301 22420
rect 13596 22380 13602 22392
rect 15289 22389 15301 22392
rect 15335 22389 15347 22423
rect 16206 22420 16212 22432
rect 16167 22392 16212 22420
rect 15289 22383 15347 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 16577 22423 16635 22429
rect 16577 22389 16589 22423
rect 16623 22420 16635 22423
rect 17770 22420 17776 22432
rect 16623 22392 17776 22420
rect 16623 22389 16635 22392
rect 16577 22383 16635 22389
rect 17770 22380 17776 22392
rect 17828 22380 17834 22432
rect 18782 22380 18788 22432
rect 18840 22420 18846 22432
rect 18969 22423 19027 22429
rect 18969 22420 18981 22423
rect 18840 22392 18981 22420
rect 18840 22380 18846 22392
rect 18969 22389 18981 22392
rect 19015 22389 19027 22423
rect 22094 22420 22100 22432
rect 22055 22392 22100 22420
rect 18969 22383 19027 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 23842 22420 23848 22432
rect 23803 22392 23848 22420
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1397 22219 1455 22225
rect 1397 22185 1409 22219
rect 1443 22216 1455 22219
rect 2130 22216 2136 22228
rect 1443 22188 2136 22216
rect 1443 22185 1455 22188
rect 1397 22179 1455 22185
rect 2130 22176 2136 22188
rect 2188 22176 2194 22228
rect 2317 22219 2375 22225
rect 2317 22185 2329 22219
rect 2363 22216 2375 22219
rect 2590 22216 2596 22228
rect 2363 22188 2596 22216
rect 2363 22185 2375 22188
rect 2317 22179 2375 22185
rect 2590 22176 2596 22188
rect 2648 22176 2654 22228
rect 2961 22219 3019 22225
rect 2961 22185 2973 22219
rect 3007 22216 3019 22219
rect 3142 22216 3148 22228
rect 3007 22188 3148 22216
rect 3007 22185 3019 22188
rect 2961 22179 3019 22185
rect 3142 22176 3148 22188
rect 3200 22216 3206 22228
rect 3970 22216 3976 22228
rect 3200 22188 3976 22216
rect 3200 22176 3206 22188
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 4341 22219 4399 22225
rect 4341 22185 4353 22219
rect 4387 22216 4399 22219
rect 5074 22216 5080 22228
rect 4387 22188 5080 22216
rect 4387 22185 4399 22188
rect 4341 22179 4399 22185
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 5460 22188 6776 22216
rect 1486 22108 1492 22160
rect 1544 22148 1550 22160
rect 5460 22148 5488 22188
rect 1544 22120 5488 22148
rect 1544 22108 1550 22120
rect 5534 22108 5540 22160
rect 5592 22148 5598 22160
rect 5813 22151 5871 22157
rect 5813 22148 5825 22151
rect 5592 22120 5825 22148
rect 5592 22108 5598 22120
rect 5813 22117 5825 22120
rect 5859 22117 5871 22151
rect 6748 22148 6776 22188
rect 6822 22176 6828 22228
rect 6880 22216 6886 22228
rect 7377 22219 7435 22225
rect 7377 22216 7389 22219
rect 6880 22188 7389 22216
rect 6880 22176 6886 22188
rect 7377 22185 7389 22188
rect 7423 22216 7435 22219
rect 7650 22216 7656 22228
rect 7423 22188 7656 22216
rect 7423 22185 7435 22188
rect 7377 22179 7435 22185
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 9401 22219 9459 22225
rect 9401 22185 9413 22219
rect 9447 22216 9459 22219
rect 9582 22216 9588 22228
rect 9447 22188 9588 22216
rect 9447 22185 9459 22188
rect 9401 22179 9459 22185
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 10229 22219 10287 22225
rect 10229 22185 10241 22219
rect 10275 22216 10287 22219
rect 14550 22216 14556 22228
rect 10275 22188 14556 22216
rect 10275 22185 10287 22188
rect 10229 22179 10287 22185
rect 7190 22148 7196 22160
rect 6748 22120 7196 22148
rect 5813 22111 5871 22117
rect 7190 22108 7196 22120
rect 7248 22108 7254 22160
rect 8389 22151 8447 22157
rect 8389 22148 8401 22151
rect 8312 22120 8401 22148
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 3053 22083 3111 22089
rect 3053 22080 3065 22083
rect 2188 22052 3065 22080
rect 2188 22040 2194 22052
rect 3053 22049 3065 22052
rect 3099 22049 3111 22083
rect 3053 22043 3111 22049
rect 4801 22083 4859 22089
rect 4801 22049 4813 22083
rect 4847 22080 4859 22083
rect 5442 22080 5448 22092
rect 4847 22052 5448 22080
rect 4847 22049 4859 22052
rect 4801 22043 4859 22049
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 5905 22083 5963 22089
rect 5905 22080 5917 22083
rect 5644 22052 5917 22080
rect 2682 22012 2688 22024
rect 1872 21984 2688 22012
rect 1872 21888 1900 21984
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 22012 3019 22015
rect 4246 22012 4252 22024
rect 3007 21984 4252 22012
rect 3007 21981 3019 21984
rect 2961 21975 3019 21981
rect 2498 21944 2504 21956
rect 2459 21916 2504 21944
rect 2498 21904 2504 21916
rect 2556 21904 2562 21956
rect 2590 21904 2596 21956
rect 2648 21944 2654 21956
rect 2976 21944 3004 21975
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 4614 21972 4620 22024
rect 4672 22012 4678 22024
rect 5644 22012 5672 22052
rect 5905 22049 5917 22052
rect 5951 22080 5963 22083
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 5951 22052 6285 22080
rect 5951 22049 5963 22052
rect 5905 22043 5963 22049
rect 6273 22049 6285 22052
rect 6319 22080 6331 22083
rect 6638 22080 6644 22092
rect 6319 22052 6644 22080
rect 6319 22049 6331 22052
rect 6273 22043 6331 22049
rect 6638 22040 6644 22052
rect 6696 22080 6702 22092
rect 7466 22080 7472 22092
rect 6696 22052 7472 22080
rect 6696 22040 6702 22052
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 8312 22080 8340 22120
rect 8389 22117 8401 22120
rect 8435 22117 8447 22151
rect 8389 22111 8447 22117
rect 8846 22108 8852 22160
rect 8904 22148 8910 22160
rect 9490 22148 9496 22160
rect 8904 22120 9496 22148
rect 8904 22108 8910 22120
rect 9490 22108 9496 22120
rect 9548 22148 9554 22160
rect 10244 22148 10272 22179
rect 14550 22176 14556 22188
rect 14608 22176 14614 22228
rect 12529 22151 12587 22157
rect 12529 22148 12541 22151
rect 9548 22120 10272 22148
rect 12360 22120 12541 22148
rect 9548 22108 9554 22120
rect 7616 22052 8340 22080
rect 7616 22040 7622 22052
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9364 22052 10364 22080
rect 9364 22040 9370 22052
rect 4672 21984 5672 22012
rect 4672 21972 4678 21984
rect 5718 21972 5724 22024
rect 5776 22012 5782 22024
rect 5813 22015 5871 22021
rect 5813 22012 5825 22015
rect 5776 21984 5825 22012
rect 5776 21972 5782 21984
rect 5813 21981 5825 21984
rect 5859 21981 5871 22015
rect 10134 22012 10140 22024
rect 10095 21984 10140 22012
rect 5813 21975 5871 21981
rect 2648 21916 3004 21944
rect 2648 21904 2654 21916
rect 3142 21904 3148 21956
rect 3200 21944 3206 21956
rect 3789 21947 3847 21953
rect 3789 21944 3801 21947
rect 3200 21916 3801 21944
rect 3200 21904 3206 21916
rect 3789 21913 3801 21916
rect 3835 21913 3847 21947
rect 5350 21944 5356 21956
rect 5311 21916 5356 21944
rect 3789 21907 3847 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 5828 21944 5856 21975
rect 10134 21972 10140 21984
rect 10192 21972 10198 22024
rect 10336 22021 10364 22052
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 12360 22080 12388 22120
rect 12529 22117 12541 22120
rect 12575 22117 12587 22151
rect 12529 22111 12587 22117
rect 13998 22108 14004 22160
rect 14056 22148 14062 22160
rect 14093 22151 14151 22157
rect 14093 22148 14105 22151
rect 14056 22120 14105 22148
rect 14056 22108 14062 22120
rect 14093 22117 14105 22120
rect 14139 22117 14151 22151
rect 14093 22111 14151 22117
rect 15749 22151 15807 22157
rect 15749 22117 15761 22151
rect 15795 22148 15807 22151
rect 16206 22148 16212 22160
rect 15795 22120 16212 22148
rect 15795 22117 15807 22120
rect 15749 22111 15807 22117
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 11940 22052 12388 22080
rect 12621 22083 12679 22089
rect 11940 22040 11946 22052
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 12710 22080 12716 22092
rect 12667 22052 12716 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 12710 22040 12716 22052
rect 12768 22080 12774 22092
rect 13449 22083 13507 22089
rect 13449 22080 13461 22083
rect 12768 22052 13461 22080
rect 12768 22040 12774 22052
rect 13449 22049 13461 22052
rect 13495 22080 13507 22083
rect 13722 22080 13728 22092
rect 13495 22052 13728 22080
rect 13495 22049 13507 22052
rect 13449 22043 13507 22049
rect 13722 22040 13728 22052
rect 13780 22080 13786 22092
rect 14185 22083 14243 22089
rect 14185 22080 14197 22083
rect 13780 22052 14197 22080
rect 13780 22040 13786 22052
rect 14185 22049 14197 22052
rect 14231 22049 14243 22083
rect 15470 22080 15476 22092
rect 15431 22052 15476 22080
rect 14185 22043 14243 22049
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 16761 22083 16819 22089
rect 16761 22049 16773 22083
rect 16807 22049 16819 22083
rect 16761 22043 16819 22049
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22080 17095 22083
rect 17862 22080 17868 22092
rect 17083 22052 17868 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10367 21984 11652 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 6086 21944 6092 21956
rect 5828 21916 6092 21944
rect 6086 21904 6092 21916
rect 6144 21904 6150 21956
rect 6914 21944 6920 21956
rect 6875 21916 6920 21944
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 9769 21947 9827 21953
rect 9769 21913 9781 21947
rect 9815 21944 9827 21947
rect 10042 21944 10048 21956
rect 9815 21916 10048 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 10042 21904 10048 21916
rect 10100 21904 10106 21956
rect 1854 21876 1860 21888
rect 1815 21848 1860 21876
rect 1854 21836 1860 21848
rect 1912 21836 1918 21888
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 2924 21848 3433 21876
rect 2924 21836 2930 21848
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 3421 21839 3479 21845
rect 4430 21836 4436 21888
rect 4488 21876 4494 21888
rect 4982 21876 4988 21888
rect 4488 21848 4988 21876
rect 4488 21836 4494 21848
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 5166 21876 5172 21888
rect 5127 21848 5172 21876
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 6730 21876 6736 21888
rect 6691 21848 6736 21876
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 7432 21848 7849 21876
rect 7432 21836 7438 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 8938 21876 8944 21888
rect 8899 21848 8944 21876
rect 7837 21839 7895 21845
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 10686 21876 10692 21888
rect 10647 21848 10692 21876
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 11624 21876 11652 21984
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 12434 22012 12440 22024
rect 11756 21984 12440 22012
rect 11756 21972 11762 21984
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 12492 21984 12585 22012
rect 12492 21972 12498 21984
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 14001 22015 14059 22021
rect 14001 22012 14013 22015
rect 13412 21984 14013 22012
rect 13412 21972 13418 21984
rect 14001 21981 14013 21984
rect 14047 21981 14059 22015
rect 16776 22012 16804 22043
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18049 22083 18107 22089
rect 18049 22049 18061 22083
rect 18095 22049 18107 22083
rect 18049 22043 18107 22049
rect 18325 22083 18383 22089
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 19334 22080 19340 22092
rect 18371 22052 19340 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 17126 22012 17132 22024
rect 16776 21984 17132 22012
rect 14001 21975 14059 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 17770 21972 17776 22024
rect 17828 22012 17834 22024
rect 18064 22012 18092 22043
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 17828 21984 18092 22012
rect 17828 21972 17834 21984
rect 12069 21947 12127 21953
rect 12069 21913 12081 21947
rect 12115 21944 12127 21947
rect 12342 21944 12348 21956
rect 12115 21916 12348 21944
rect 12115 21913 12127 21916
rect 12069 21907 12127 21913
rect 12342 21904 12348 21916
rect 12400 21904 12406 21956
rect 12986 21904 12992 21956
rect 13044 21944 13050 21956
rect 13081 21947 13139 21953
rect 13081 21944 13093 21947
rect 13044 21916 13093 21944
rect 13044 21904 13050 21916
rect 13081 21913 13093 21916
rect 13127 21944 13139 21947
rect 13633 21947 13691 21953
rect 13633 21944 13645 21947
rect 13127 21916 13645 21944
rect 13127 21913 13139 21916
rect 13081 21907 13139 21913
rect 13633 21913 13645 21916
rect 13679 21913 13691 21947
rect 13633 21907 13691 21913
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 20346 21944 20352 21956
rect 19567 21916 20352 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 13538 21876 13544 21888
rect 11624 21848 13544 21876
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 14642 21876 14648 21888
rect 14603 21848 14648 21876
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2130 21672 2136 21684
rect 2091 21644 2136 21672
rect 2130 21632 2136 21644
rect 2188 21672 2194 21684
rect 3786 21672 3792 21684
rect 2188 21644 3792 21672
rect 2188 21632 2194 21644
rect 3786 21632 3792 21644
rect 3844 21672 3850 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3844 21644 3985 21672
rect 3844 21632 3850 21644
rect 3973 21641 3985 21644
rect 4019 21641 4031 21675
rect 3973 21635 4031 21641
rect 4522 21632 4528 21684
rect 4580 21672 4586 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 4580 21644 4905 21672
rect 4580 21632 4586 21644
rect 4893 21641 4905 21644
rect 4939 21641 4951 21675
rect 4893 21635 4951 21641
rect 4614 21604 4620 21616
rect 4575 21576 4620 21604
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 4908 21536 4936 21635
rect 4982 21632 4988 21684
rect 5040 21672 5046 21684
rect 6086 21672 6092 21684
rect 5040 21644 5571 21672
rect 6047 21644 6092 21672
rect 5040 21632 5046 21644
rect 5169 21607 5227 21613
rect 5169 21573 5181 21607
rect 5215 21604 5227 21607
rect 5442 21604 5448 21616
rect 5215 21576 5448 21604
rect 5215 21573 5227 21576
rect 5169 21567 5227 21573
rect 5442 21564 5448 21576
rect 5500 21564 5506 21616
rect 5543 21604 5571 21644
rect 6086 21632 6092 21644
rect 6144 21632 6150 21684
rect 6641 21675 6699 21681
rect 6641 21641 6653 21675
rect 6687 21672 6699 21675
rect 6822 21672 6828 21684
rect 6687 21644 6828 21672
rect 6687 21641 6699 21644
rect 6641 21635 6699 21641
rect 6656 21604 6684 21635
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 7190 21632 7196 21684
rect 7248 21672 7254 21684
rect 7650 21672 7656 21684
rect 7248 21644 7656 21672
rect 7248 21632 7254 21644
rect 7650 21632 7656 21644
rect 7708 21672 7714 21684
rect 7837 21675 7895 21681
rect 7837 21672 7849 21675
rect 7708 21644 7849 21672
rect 7708 21632 7714 21644
rect 7837 21641 7849 21644
rect 7883 21641 7895 21675
rect 9490 21672 9496 21684
rect 9451 21644 9496 21672
rect 7837 21635 7895 21641
rect 9490 21632 9496 21644
rect 9548 21632 9554 21684
rect 11698 21672 11704 21684
rect 11659 21644 11704 21672
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 12529 21675 12587 21681
rect 12529 21641 12541 21675
rect 12575 21672 12587 21675
rect 12894 21672 12900 21684
rect 12575 21644 12900 21672
rect 12575 21641 12587 21644
rect 12529 21635 12587 21641
rect 12894 21632 12900 21644
rect 12952 21632 12958 21684
rect 15470 21672 15476 21684
rect 15431 21644 15476 21672
rect 15470 21632 15476 21644
rect 15528 21632 15534 21684
rect 19521 21675 19579 21681
rect 19521 21641 19533 21675
rect 19567 21672 19579 21675
rect 19978 21672 19984 21684
rect 19567 21644 19984 21672
rect 19567 21641 19579 21644
rect 19521 21635 19579 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 20622 21672 20628 21684
rect 20583 21644 20628 21672
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 6914 21604 6920 21616
rect 5543 21576 6684 21604
rect 6875 21576 6920 21604
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 8478 21604 8484 21616
rect 8439 21576 8484 21604
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 10045 21607 10103 21613
rect 10045 21573 10057 21607
rect 10091 21604 10103 21607
rect 10134 21604 10140 21616
rect 10091 21576 10140 21604
rect 10091 21573 10103 21576
rect 10045 21567 10103 21573
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 11333 21607 11391 21613
rect 11333 21573 11345 21607
rect 11379 21604 11391 21607
rect 12710 21604 12716 21616
rect 11379 21576 12716 21604
rect 11379 21573 11391 21576
rect 11333 21567 11391 21573
rect 12710 21564 12716 21576
rect 12768 21564 12774 21616
rect 14093 21607 14151 21613
rect 14093 21573 14105 21607
rect 14139 21604 14151 21607
rect 15010 21604 15016 21616
rect 14139 21576 15016 21604
rect 14139 21573 14151 21576
rect 14093 21567 14151 21573
rect 15010 21564 15016 21576
rect 15068 21564 15074 21616
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 19889 21607 19947 21613
rect 19889 21604 19901 21607
rect 19392 21576 19901 21604
rect 19392 21564 19398 21576
rect 19889 21573 19901 21576
rect 19935 21573 19947 21607
rect 19889 21567 19947 21573
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 4908 21508 5549 21536
rect 5537 21505 5549 21508
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 7098 21536 7104 21548
rect 6788 21508 7104 21536
rect 6788 21496 6794 21508
rect 7098 21496 7104 21508
rect 7156 21536 7162 21548
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 7156 21508 7481 21536
rect 7156 21496 7162 21508
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8996 21508 9045 21536
rect 8996 21496 9002 21508
rect 9033 21505 9045 21508
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21536 10655 21539
rect 10686 21536 10692 21548
rect 10643 21508 10692 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 12894 21496 12900 21548
rect 12952 21536 12958 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12952 21508 13093 21536
rect 12952 21496 12958 21508
rect 13081 21505 13093 21508
rect 13127 21536 13139 21539
rect 13446 21536 13452 21548
rect 13127 21508 13452 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 14642 21536 14648 21548
rect 14603 21508 14648 21536
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 16206 21536 16212 21548
rect 16167 21508 16212 21536
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16666 21536 16672 21548
rect 16627 21508 16672 21536
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 18325 21539 18383 21545
rect 18325 21505 18337 21539
rect 18371 21536 18383 21539
rect 19150 21536 19156 21548
rect 18371 21508 19156 21536
rect 18371 21505 18383 21508
rect 18325 21499 18383 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 2593 21471 2651 21477
rect 2593 21437 2605 21471
rect 2639 21437 2651 21471
rect 2593 21431 2651 21437
rect 1486 21360 1492 21412
rect 1544 21400 1550 21412
rect 2409 21403 2467 21409
rect 2409 21400 2421 21403
rect 1544 21372 2421 21400
rect 1544 21360 1550 21372
rect 2409 21369 2421 21372
rect 2455 21400 2467 21403
rect 2608 21400 2636 21431
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5718 21468 5724 21480
rect 5224 21440 5724 21468
rect 5224 21428 5230 21440
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 7558 21468 7564 21480
rect 7239 21440 7564 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 9858 21428 9864 21480
rect 9916 21468 9922 21480
rect 12802 21468 12808 21480
rect 9916 21440 10548 21468
rect 12763 21440 12808 21468
rect 9916 21428 9922 21440
rect 2866 21409 2872 21412
rect 2860 21400 2872 21409
rect 2455 21372 2636 21400
rect 2827 21372 2872 21400
rect 2455 21369 2467 21372
rect 2409 21363 2467 21369
rect 2860 21363 2872 21372
rect 2866 21360 2872 21363
rect 2924 21360 2930 21412
rect 5258 21360 5264 21412
rect 5316 21400 5322 21412
rect 5629 21403 5687 21409
rect 5629 21400 5641 21403
rect 5316 21372 5641 21400
rect 5316 21360 5322 21372
rect 5629 21369 5641 21372
rect 5675 21400 5687 21403
rect 5994 21400 6000 21412
rect 5675 21372 6000 21400
rect 5675 21369 5687 21372
rect 5629 21363 5687 21369
rect 5994 21360 6000 21372
rect 6052 21360 6058 21412
rect 7374 21400 7380 21412
rect 7335 21372 7380 21400
rect 7374 21360 7380 21372
rect 7432 21360 7438 21412
rect 8297 21403 8355 21409
rect 8297 21369 8309 21403
rect 8343 21400 8355 21403
rect 8478 21400 8484 21412
rect 8343 21372 8484 21400
rect 8343 21369 8355 21372
rect 8297 21363 8355 21369
rect 8478 21360 8484 21372
rect 8536 21400 8542 21412
rect 10520 21409 10548 21440
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 16224 21468 16252 21496
rect 16393 21471 16451 21477
rect 16393 21468 16405 21471
rect 14056 21440 15148 21468
rect 16224 21440 16405 21468
rect 14056 21428 14062 21440
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 8536 21372 8769 21400
rect 8536 21360 8542 21372
rect 8757 21369 8769 21372
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 10321 21403 10379 21409
rect 10321 21369 10333 21403
rect 10367 21369 10379 21403
rect 10321 21363 10379 21369
rect 10505 21403 10563 21409
rect 10505 21369 10517 21403
rect 10551 21369 10563 21403
rect 12986 21400 12992 21412
rect 12947 21372 12992 21400
rect 10505 21363 10563 21369
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 8846 21292 8852 21344
rect 8904 21332 8910 21344
rect 8941 21335 8999 21341
rect 8941 21332 8953 21335
rect 8904 21304 8953 21332
rect 8904 21292 8910 21304
rect 8941 21301 8953 21304
rect 8987 21301 8999 21335
rect 9766 21332 9772 21344
rect 9727 21304 9772 21332
rect 8941 21295 8999 21301
rect 9766 21292 9772 21304
rect 9824 21332 9830 21344
rect 10336 21332 10364 21363
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 14369 21403 14427 21409
rect 14369 21400 14381 21403
rect 14148 21372 14381 21400
rect 14148 21360 14154 21372
rect 14369 21369 14381 21372
rect 14415 21369 14427 21403
rect 14369 21363 14427 21369
rect 15120 21344 15148 21440
rect 16393 21437 16405 21440
rect 16439 21437 16451 21471
rect 17126 21468 17132 21480
rect 17087 21440 17132 21468
rect 16393 21431 16451 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 18046 21468 18052 21480
rect 18007 21440 18052 21468
rect 18046 21428 18052 21440
rect 18104 21468 18110 21480
rect 18785 21471 18843 21477
rect 18785 21468 18797 21471
rect 18104 21440 18797 21468
rect 18104 21428 18110 21440
rect 18785 21437 18797 21440
rect 18831 21437 18843 21471
rect 18785 21431 18843 21437
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21437 19395 21471
rect 20438 21468 20444 21480
rect 20399 21440 20444 21468
rect 19337 21431 19395 21437
rect 19352 21344 19380 21431
rect 20438 21428 20444 21440
rect 20496 21468 20502 21480
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20496 21440 21005 21468
rect 20496 21428 20502 21440
rect 20993 21437 21005 21440
rect 21039 21437 21051 21471
rect 20993 21431 21051 21437
rect 9824 21304 10364 21332
rect 9824 21292 9830 21304
rect 11698 21292 11704 21344
rect 11756 21332 11762 21344
rect 11882 21332 11888 21344
rect 11756 21304 11888 21332
rect 11756 21292 11762 21304
rect 11882 21292 11888 21304
rect 11940 21332 11946 21344
rect 11977 21335 12035 21341
rect 11977 21332 11989 21335
rect 11940 21304 11989 21332
rect 11940 21292 11946 21304
rect 11977 21301 11989 21304
rect 12023 21301 12035 21335
rect 11977 21295 12035 21301
rect 13354 21292 13360 21344
rect 13412 21332 13418 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 13412 21304 13553 21332
rect 13412 21292 13418 21304
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 14550 21332 14556 21344
rect 14511 21304 14556 21332
rect 13541 21295 13599 21301
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 15102 21332 15108 21344
rect 15063 21304 15108 21332
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 17770 21332 17776 21344
rect 17731 21304 17776 21332
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 19245 21335 19303 21341
rect 19245 21301 19257 21335
rect 19291 21332 19303 21335
rect 19334 21332 19340 21344
rect 19291 21304 19340 21332
rect 19291 21301 19303 21304
rect 19245 21295 19303 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2866 21128 2872 21140
rect 2779 21100 2872 21128
rect 2866 21088 2872 21100
rect 2924 21128 2930 21140
rect 4617 21131 4675 21137
rect 2924 21100 3556 21128
rect 2924 21088 2930 21100
rect 1756 21063 1814 21069
rect 1756 21029 1768 21063
rect 1802 21060 1814 21063
rect 1854 21060 1860 21072
rect 1802 21032 1860 21060
rect 1802 21029 1814 21032
rect 1756 21023 1814 21029
rect 1854 21020 1860 21032
rect 1912 21020 1918 21072
rect 3528 21001 3556 21100
rect 4617 21097 4629 21131
rect 4663 21128 4675 21131
rect 4982 21128 4988 21140
rect 4663 21100 4988 21128
rect 4663 21097 4675 21100
rect 4617 21091 4675 21097
rect 4982 21088 4988 21100
rect 5040 21088 5046 21140
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5258 21128 5264 21140
rect 5215 21100 5264 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 5534 21128 5540 21140
rect 5495 21100 5540 21128
rect 5534 21088 5540 21100
rect 5592 21088 5598 21140
rect 7098 21128 7104 21140
rect 7059 21100 7104 21128
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 7653 21131 7711 21137
rect 7653 21128 7665 21131
rect 7616 21100 7665 21128
rect 7616 21088 7622 21100
rect 7653 21097 7665 21100
rect 7699 21097 7711 21131
rect 8478 21128 8484 21140
rect 8439 21100 8484 21128
rect 7653 21091 7711 21097
rect 8478 21088 8484 21100
rect 8536 21088 8542 21140
rect 9306 21088 9312 21140
rect 9364 21128 9370 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 9364 21100 9413 21128
rect 9364 21088 9370 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 9401 21091 9459 21097
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 9916 21100 9965 21128
rect 9916 21088 9922 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 10042 21088 10048 21140
rect 10100 21128 10106 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 10100 21100 10333 21128
rect 10100 21088 10106 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10321 21091 10379 21097
rect 12529 21131 12587 21137
rect 12529 21097 12541 21131
rect 12575 21128 12587 21131
rect 12802 21128 12808 21140
rect 12575 21100 12808 21128
rect 12575 21097 12587 21100
rect 12529 21091 12587 21097
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 12952 21100 12997 21128
rect 13188 21100 13645 21128
rect 12952 21088 12958 21100
rect 4433 21063 4491 21069
rect 4433 21029 4445 21063
rect 4479 21060 4491 21063
rect 4522 21060 4528 21072
rect 4479 21032 4528 21060
rect 4479 21029 4491 21032
rect 4433 21023 4491 21029
rect 4522 21020 4528 21032
rect 4580 21060 4586 21072
rect 5552 21060 5580 21088
rect 4580 21032 5580 21060
rect 4580 21020 4586 21032
rect 5718 21020 5724 21072
rect 5776 21060 5782 21072
rect 5966 21063 6024 21069
rect 5966 21060 5978 21063
rect 5776 21032 5978 21060
rect 5776 21020 5782 21032
rect 5966 21029 5978 21032
rect 6012 21029 6024 21063
rect 5966 21023 6024 21029
rect 10686 21020 10692 21072
rect 10744 21069 10750 21072
rect 10744 21063 10808 21069
rect 10744 21029 10762 21063
rect 10796 21029 10808 21063
rect 10744 21023 10808 21029
rect 10744 21020 10750 21023
rect 10962 21020 10968 21072
rect 11020 21020 11026 21072
rect 12986 21020 12992 21072
rect 13044 21060 13050 21072
rect 13188 21060 13216 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 15010 21128 15016 21140
rect 14971 21100 15016 21128
rect 13633 21091 13691 21097
rect 15010 21088 15016 21100
rect 15068 21128 15074 21140
rect 15933 21131 15991 21137
rect 15933 21128 15945 21131
rect 15068 21100 15945 21128
rect 15068 21088 15074 21100
rect 15933 21097 15945 21100
rect 15979 21097 15991 21131
rect 21082 21128 21088 21140
rect 21043 21100 21088 21128
rect 15933 21091 15991 21097
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 13044 21032 13216 21060
rect 13044 21020 13050 21032
rect 13262 21020 13268 21072
rect 13320 21060 13326 21072
rect 13449 21063 13507 21069
rect 13449 21060 13461 21063
rect 13320 21032 13461 21060
rect 13320 21020 13326 21032
rect 13449 21029 13461 21032
rect 13495 21029 13507 21063
rect 17494 21060 17500 21072
rect 17455 21032 17500 21060
rect 13449 21023 13507 21029
rect 3513 20995 3571 21001
rect 3513 20961 3525 20995
rect 3559 20992 3571 20995
rect 3881 20995 3939 21001
rect 3881 20992 3893 20995
rect 3559 20964 3893 20992
rect 3559 20961 3571 20964
rect 3513 20955 3571 20961
rect 3881 20961 3893 20964
rect 3927 20992 3939 20995
rect 4709 20995 4767 21001
rect 4709 20992 4721 20995
rect 3927 20964 4721 20992
rect 3927 20961 3939 20964
rect 3881 20955 3939 20961
rect 4709 20961 4721 20964
rect 4755 20961 4767 20995
rect 4709 20955 4767 20961
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 10980 20992 11008 21020
rect 10551 20964 11008 20992
rect 13464 20992 13492 21023
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 18782 21060 18788 21072
rect 18743 21032 18788 21060
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 13814 20992 13820 21004
rect 13464 20964 13820 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 13814 20952 13820 20964
rect 13872 20952 13878 21004
rect 15470 20952 15476 21004
rect 15528 20992 15534 21004
rect 15749 20995 15807 21001
rect 15749 20992 15761 20995
rect 15528 20964 15761 20992
rect 15528 20952 15534 20964
rect 15749 20961 15761 20964
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 16853 20995 16911 21001
rect 16853 20961 16865 20995
rect 16899 20992 16911 20995
rect 17586 20992 17592 21004
rect 16899 20964 17592 20992
rect 16899 20961 16911 20964
rect 16853 20955 16911 20961
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 18509 20995 18567 21001
rect 18509 20992 18521 20995
rect 17972 20964 18521 20992
rect 1486 20924 1492 20936
rect 1447 20896 1492 20924
rect 1486 20884 1492 20896
rect 1544 20884 1550 20936
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20893 5779 20927
rect 5721 20887 5779 20893
rect 4154 20856 4160 20868
rect 4115 20828 4160 20856
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 5736 20788 5764 20887
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 13722 20924 13728 20936
rect 12492 20896 13728 20924
rect 12492 20884 12498 20896
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 17092 20896 17417 20924
rect 17092 20884 17098 20896
rect 17405 20893 17417 20896
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 12526 20816 12532 20868
rect 12584 20856 12590 20868
rect 13262 20856 13268 20868
rect 12584 20828 13268 20856
rect 12584 20816 12590 20828
rect 13262 20816 13268 20828
rect 13320 20816 13326 20868
rect 15473 20859 15531 20865
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 17972 20856 18000 20964
rect 18509 20961 18521 20964
rect 18555 20992 18567 20995
rect 19058 20992 19064 21004
rect 18555 20964 19064 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 21082 20992 21088 21004
rect 20947 20964 21088 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 15519 20828 18000 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 6638 20788 6644 20800
rect 5736 20760 6644 20788
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8846 20788 8852 20800
rect 8352 20760 8852 20788
rect 8352 20748 8358 20760
rect 8846 20748 8852 20760
rect 8904 20788 8910 20800
rect 8941 20791 8999 20797
rect 8941 20788 8953 20791
rect 8904 20760 8953 20788
rect 8904 20748 8910 20760
rect 8941 20757 8953 20760
rect 8987 20757 8999 20791
rect 8941 20751 8999 20757
rect 11885 20791 11943 20797
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 12342 20788 12348 20800
rect 11931 20760 12348 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 12342 20748 12348 20760
rect 12400 20748 12406 20800
rect 13170 20788 13176 20800
rect 13131 20760 13176 20788
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 14090 20788 14096 20800
rect 14051 20760 14096 20788
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14550 20788 14556 20800
rect 14463 20760 14556 20788
rect 14550 20748 14556 20760
rect 14608 20788 14614 20800
rect 15286 20788 15292 20800
rect 14608 20760 15292 20788
rect 14608 20748 14614 20760
rect 15286 20748 15292 20760
rect 15344 20748 15350 20800
rect 17037 20791 17095 20797
rect 17037 20757 17049 20791
rect 17083 20788 17095 20791
rect 17954 20788 17960 20800
rect 17083 20760 17960 20788
rect 17083 20757 17095 20760
rect 17037 20751 17095 20757
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18690 20788 18696 20800
rect 18187 20760 18696 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2590 20584 2596 20596
rect 1995 20556 2596 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 2590 20544 2596 20556
rect 2648 20544 2654 20596
rect 3789 20587 3847 20593
rect 3789 20553 3801 20587
rect 3835 20584 3847 20587
rect 4982 20584 4988 20596
rect 3835 20556 4988 20584
rect 3835 20553 3847 20556
rect 3789 20547 3847 20553
rect 4982 20544 4988 20556
rect 5040 20544 5046 20596
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 5629 20587 5687 20593
rect 5629 20584 5641 20587
rect 5592 20556 5641 20584
rect 5592 20544 5598 20556
rect 5629 20553 5641 20556
rect 5675 20553 5687 20587
rect 10686 20584 10692 20596
rect 10647 20556 10692 20584
rect 5629 20547 5687 20553
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 11112 20556 11253 20584
rect 11112 20544 11118 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 12434 20584 12440 20596
rect 11931 20556 12440 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 3421 20519 3479 20525
rect 3421 20485 3433 20519
rect 3467 20516 3479 20519
rect 4246 20516 4252 20528
rect 3467 20488 4252 20516
rect 3467 20485 3479 20488
rect 3421 20479 3479 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 11256 20516 11284 20547
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 13872 20556 14381 20584
rect 13872 20544 13878 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14369 20547 14427 20553
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 16485 20587 16543 20593
rect 16485 20584 16497 20587
rect 16080 20556 16497 20584
rect 16080 20544 16086 20556
rect 16485 20553 16497 20556
rect 16531 20553 16543 20587
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 16485 20547 16543 20553
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 19058 20584 19064 20596
rect 19019 20556 19064 20584
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 11256 20488 12173 20516
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12161 20479 12219 20485
rect 18141 20519 18199 20525
rect 18141 20485 18153 20519
rect 18187 20485 18199 20519
rect 18141 20479 18199 20485
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20448 2559 20451
rect 2682 20448 2688 20460
rect 2547 20420 2688 20448
rect 2547 20417 2559 20420
rect 2501 20411 2559 20417
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9306 20448 9312 20460
rect 9263 20420 9312 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 2222 20380 2228 20392
rect 2183 20352 2228 20380
rect 2222 20340 2228 20352
rect 2280 20380 2286 20392
rect 7098 20389 7104 20392
rect 2869 20383 2927 20389
rect 2869 20380 2881 20383
rect 2280 20352 2881 20380
rect 2280 20340 2286 20352
rect 2869 20349 2881 20352
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 4157 20383 4215 20389
rect 4157 20349 4169 20383
rect 4203 20380 4215 20383
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 4203 20352 4261 20380
rect 4203 20349 4215 20352
rect 4157 20343 4215 20349
rect 4249 20349 4261 20352
rect 4295 20380 4307 20383
rect 6825 20383 6883 20389
rect 4295 20352 6316 20380
rect 4295 20349 4307 20352
rect 4249 20343 4307 20349
rect 1670 20272 1676 20324
rect 1728 20312 1734 20324
rect 2409 20315 2467 20321
rect 2409 20312 2421 20315
rect 1728 20284 2421 20312
rect 1728 20272 1734 20284
rect 2409 20281 2421 20284
rect 2455 20281 2467 20315
rect 2409 20275 2467 20281
rect 3786 20272 3792 20324
rect 3844 20312 3850 20324
rect 6288 20321 6316 20352
rect 6825 20349 6837 20383
rect 6871 20349 6883 20383
rect 7092 20380 7104 20389
rect 7059 20352 7104 20380
rect 6825 20343 6883 20349
rect 7092 20343 7104 20352
rect 4494 20315 4552 20321
rect 4494 20312 4506 20315
rect 3844 20284 4506 20312
rect 3844 20272 3850 20284
rect 4494 20281 4506 20284
rect 4540 20281 4552 20315
rect 4494 20275 4552 20281
rect 6273 20315 6331 20321
rect 6273 20281 6285 20315
rect 6319 20312 6331 20315
rect 6638 20312 6644 20324
rect 6319 20284 6644 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 6638 20272 6644 20284
rect 6696 20312 6702 20324
rect 6840 20312 6868 20343
rect 7098 20340 7104 20343
rect 7156 20340 7162 20392
rect 9232 20380 9260 20411
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 7208 20352 9260 20380
rect 12176 20380 12204 20479
rect 12342 20380 12348 20392
rect 12176 20352 12348 20380
rect 7208 20312 7236 20352
rect 12342 20340 12348 20352
rect 12400 20380 12406 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12400 20352 12449 20380
rect 12400 20340 12406 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 15105 20383 15163 20389
rect 15105 20380 15117 20383
rect 15059 20352 15117 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 15105 20349 15117 20352
rect 15151 20380 15163 20383
rect 16206 20380 16212 20392
rect 15151 20352 16212 20380
rect 15151 20349 15163 20352
rect 15105 20343 15163 20349
rect 16206 20340 16212 20352
rect 16264 20340 16270 20392
rect 18156 20380 18184 20479
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19797 20451 19855 20457
rect 19797 20448 19809 20451
rect 19392 20420 19809 20448
rect 19392 20408 19398 20420
rect 19797 20417 19809 20420
rect 19843 20417 19855 20451
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 19797 20411 19855 20417
rect 21082 20408 21088 20420
rect 21140 20448 21146 20460
rect 21637 20451 21695 20457
rect 21637 20448 21649 20451
rect 21140 20420 21649 20448
rect 21140 20408 21146 20420
rect 21637 20417 21649 20420
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 18156 20352 19625 20380
rect 19613 20349 19625 20352
rect 19659 20380 19671 20383
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 19659 20352 20361 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 20349 20349 20361 20352
rect 20395 20349 20407 20383
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20349 20343 20407 20349
rect 20732 20352 20913 20380
rect 6696 20284 7236 20312
rect 6696 20272 6702 20284
rect 8938 20272 8944 20324
rect 8996 20312 9002 20324
rect 9398 20312 9404 20324
rect 8996 20284 9404 20312
rect 8996 20272 9002 20284
rect 9398 20272 9404 20284
rect 9456 20312 9462 20324
rect 9554 20315 9612 20321
rect 9554 20312 9566 20315
rect 9456 20284 9566 20312
rect 9456 20272 9462 20284
rect 9554 20281 9566 20284
rect 9600 20281 9612 20315
rect 9554 20275 9612 20281
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 12682 20315 12740 20321
rect 12682 20312 12694 20315
rect 12584 20284 12694 20312
rect 12584 20272 12590 20284
rect 12682 20281 12694 20284
rect 12728 20281 12740 20315
rect 12682 20275 12740 20281
rect 14642 20272 14648 20324
rect 14700 20312 14706 20324
rect 15378 20321 15384 20324
rect 15350 20315 15384 20321
rect 15350 20312 15362 20315
rect 14700 20284 15362 20312
rect 14700 20272 14706 20284
rect 15350 20281 15362 20284
rect 15436 20312 15442 20324
rect 18417 20315 18475 20321
rect 15436 20284 15498 20312
rect 15350 20275 15384 20281
rect 15378 20272 15384 20275
rect 15436 20272 15442 20284
rect 18417 20281 18429 20315
rect 18463 20281 18475 20315
rect 18417 20275 18475 20281
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 8168 20216 8217 20244
rect 8168 20204 8174 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 8205 20207 8263 20213
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17770 20244 17776 20256
rect 17731 20216 17776 20244
rect 17770 20204 17776 20216
rect 17828 20244 17834 20256
rect 18432 20244 18460 20275
rect 20732 20256 20760 20352
rect 20901 20349 20913 20352
rect 20947 20349 20959 20383
rect 20901 20343 20959 20349
rect 18598 20244 18604 20256
rect 17828 20216 18460 20244
rect 18559 20216 18604 20244
rect 17828 20204 17834 20216
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 20714 20244 20720 20256
rect 20675 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2314 20000 2320 20052
rect 2372 20040 2378 20052
rect 2498 20040 2504 20052
rect 2372 20012 2504 20040
rect 2372 20000 2378 20012
rect 2498 20000 2504 20012
rect 2556 20040 2562 20052
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2556 20012 2605 20040
rect 2556 20000 2562 20012
rect 2593 20009 2605 20012
rect 2639 20009 2651 20043
rect 2593 20003 2651 20009
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3510 20040 3516 20052
rect 3191 20012 3516 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 2682 19972 2688 19984
rect 2595 19944 2688 19972
rect 2682 19932 2688 19944
rect 2740 19972 2746 19984
rect 3160 19972 3188 20003
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3786 20040 3792 20052
rect 3747 20012 3792 20040
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 4239 20043 4297 20049
rect 4239 20009 4251 20043
rect 4285 20040 4297 20043
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 4285 20012 6285 20040
rect 4285 20009 4297 20012
rect 4239 20003 4297 20009
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7098 20040 7104 20052
rect 6963 20012 7104 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 4522 19972 4528 19984
rect 2740 19944 3188 19972
rect 4483 19944 4528 19972
rect 2740 19932 2746 19944
rect 4522 19932 4528 19944
rect 4580 19932 4586 19984
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19972 4767 19975
rect 4982 19972 4988 19984
rect 4755 19944 4988 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 5534 19972 5540 19984
rect 5495 19944 5540 19972
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 6288 19972 6316 20003
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 8021 20043 8079 20049
rect 8021 20040 8033 20043
rect 7708 20012 8033 20040
rect 7708 20000 7714 20012
rect 8021 20009 8033 20012
rect 8067 20009 8079 20043
rect 9398 20040 9404 20052
rect 9359 20012 9404 20040
rect 8021 20003 8079 20009
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 12526 20040 12532 20052
rect 12487 20012 12532 20040
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13780 20012 14105 20040
rect 13780 20000 13786 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14700 20012 15025 20040
rect 14700 20000 14706 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 17586 20040 17592 20052
rect 17547 20012 17592 20040
rect 15013 20003 15071 20009
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18012 20012 18521 20040
rect 18012 20000 18018 20012
rect 18509 20009 18521 20012
rect 18555 20040 18567 20043
rect 18598 20040 18604 20052
rect 18555 20012 18604 20040
rect 18555 20009 18567 20012
rect 18509 20003 18567 20009
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 21266 20040 21272 20052
rect 21227 20012 21272 20040
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 22465 20043 22523 20049
rect 22465 20009 22477 20043
rect 22511 20040 22523 20043
rect 23382 20040 23388 20052
rect 22511 20012 23388 20040
rect 22511 20009 22523 20012
rect 22465 20003 22523 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 7193 19975 7251 19981
rect 7193 19972 7205 19975
rect 6288 19944 7205 19972
rect 7193 19941 7205 19944
rect 7239 19941 7251 19975
rect 11698 19972 11704 19984
rect 11659 19944 11704 19972
rect 7193 19935 7251 19941
rect 11698 19932 11704 19944
rect 11756 19932 11762 19984
rect 12980 19975 13038 19981
rect 12980 19972 12992 19975
rect 12176 19944 12992 19972
rect 1854 19864 1860 19916
rect 1912 19904 1918 19916
rect 2409 19907 2467 19913
rect 2409 19904 2421 19907
rect 1912 19876 2421 19904
rect 1912 19864 1918 19876
rect 2409 19873 2421 19876
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 5442 19864 5448 19916
rect 5500 19904 5506 19916
rect 6089 19907 6147 19913
rect 6089 19904 6101 19907
rect 5500 19876 6101 19904
rect 5500 19864 5506 19876
rect 6089 19873 6101 19876
rect 6135 19904 6147 19907
rect 8481 19907 8539 19913
rect 8481 19904 8493 19907
rect 6135 19876 8493 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 8481 19873 8493 19876
rect 8527 19873 8539 19907
rect 11514 19904 11520 19916
rect 11475 19876 11520 19904
rect 8481 19867 8539 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 12176 19848 12204 19944
rect 12980 19941 12992 19944
rect 13026 19972 13038 19975
rect 13814 19972 13820 19984
rect 13026 19944 13820 19972
rect 13026 19941 13038 19944
rect 12980 19935 13038 19941
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 15933 19975 15991 19981
rect 15933 19941 15945 19975
rect 15979 19972 15991 19975
rect 16022 19972 16028 19984
rect 15979 19944 16028 19972
rect 15979 19941 15991 19944
rect 15933 19935 15991 19941
rect 16022 19932 16028 19944
rect 16080 19972 16086 19984
rect 16454 19975 16512 19981
rect 16454 19972 16466 19975
rect 16080 19944 16466 19972
rect 16080 19932 16086 19944
rect 16454 19941 16466 19944
rect 16500 19972 16512 19975
rect 16574 19972 16580 19984
rect 16500 19944 16580 19972
rect 16500 19941 16512 19944
rect 16454 19935 16512 19941
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 17604 19972 17632 20000
rect 18138 19972 18144 19984
rect 17604 19944 18144 19972
rect 18138 19932 18144 19944
rect 18196 19932 18202 19984
rect 19337 19975 19395 19981
rect 19337 19941 19349 19975
rect 19383 19972 19395 19975
rect 20438 19972 20444 19984
rect 19383 19944 20444 19972
rect 19383 19941 19395 19944
rect 19337 19935 19395 19941
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 19058 19904 19064 19916
rect 19019 19876 19064 19904
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 21082 19904 21088 19916
rect 21043 19876 21088 19904
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 22281 19907 22339 19913
rect 22281 19873 22293 19907
rect 22327 19904 22339 19907
rect 22830 19904 22836 19916
rect 22327 19876 22836 19904
rect 22327 19873 22339 19876
rect 22281 19867 22339 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19836 4859 19839
rect 5166 19836 5172 19848
rect 4847 19808 5172 19836
rect 4847 19805 4859 19808
rect 4801 19799 4859 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 6362 19836 6368 19848
rect 6323 19808 6368 19836
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 7926 19836 7932 19848
rect 7887 19808 7932 19836
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 8110 19836 8116 19848
rect 8071 19808 8116 19836
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 10502 19836 10508 19848
rect 10183 19808 10508 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 11793 19839 11851 19845
rect 11793 19805 11805 19839
rect 11839 19836 11851 19839
rect 12158 19836 12164 19848
rect 11839 19808 12164 19836
rect 11839 19805 11851 19808
rect 11793 19799 11851 19805
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 12710 19836 12716 19848
rect 12400 19808 12716 19836
rect 12400 19796 12406 19808
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 16206 19836 16212 19848
rect 16167 19808 16212 19836
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 2133 19771 2191 19777
rect 2133 19737 2145 19771
rect 2179 19768 2191 19771
rect 2590 19768 2596 19780
rect 2179 19740 2596 19768
rect 2179 19737 2191 19740
rect 2133 19731 2191 19737
rect 2590 19728 2596 19740
rect 2648 19768 2654 19780
rect 3142 19768 3148 19780
rect 2648 19740 3148 19768
rect 2648 19728 2654 19740
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 5810 19768 5816 19780
rect 5771 19740 5816 19768
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 7561 19771 7619 19777
rect 7561 19737 7573 19771
rect 7607 19768 7619 19771
rect 8202 19768 8208 19780
rect 7607 19740 8208 19768
rect 7607 19737 7619 19740
rect 7561 19731 7619 19737
rect 8202 19728 8208 19740
rect 8260 19728 8266 19780
rect 11241 19771 11299 19777
rect 11241 19737 11253 19771
rect 11287 19768 11299 19771
rect 11287 19740 12480 19768
rect 11287 19737 11299 19740
rect 11241 19731 11299 19737
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 1673 19703 1731 19709
rect 1673 19700 1685 19703
rect 1544 19672 1685 19700
rect 1544 19660 1550 19672
rect 1673 19669 1685 19672
rect 1719 19700 1731 19703
rect 1946 19700 1952 19712
rect 1719 19672 1952 19700
rect 1719 19669 1731 19672
rect 1673 19663 1731 19669
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 5074 19660 5080 19712
rect 5132 19700 5138 19712
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 5132 19672 5181 19700
rect 5132 19660 5138 19672
rect 5169 19669 5181 19672
rect 5215 19669 5227 19703
rect 12452 19700 12480 19740
rect 12986 19700 12992 19712
rect 12452 19672 12992 19700
rect 5169 19663 5227 19669
rect 12986 19660 12992 19672
rect 13044 19700 13050 19712
rect 14645 19703 14703 19709
rect 14645 19700 14657 19703
rect 13044 19672 14657 19700
rect 13044 19660 13050 19672
rect 14645 19669 14657 19672
rect 14691 19669 14703 19703
rect 15470 19700 15476 19712
rect 15431 19672 15476 19700
rect 14645 19663 14703 19669
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 4065 19499 4123 19505
rect 4065 19465 4077 19499
rect 4111 19496 4123 19499
rect 4982 19496 4988 19508
rect 4111 19468 4988 19496
rect 4111 19465 4123 19468
rect 4065 19459 4123 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5997 19499 6055 19505
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 6362 19496 6368 19508
rect 6043 19468 6368 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 7561 19499 7619 19505
rect 7561 19465 7573 19499
rect 7607 19496 7619 19499
rect 7926 19496 7932 19508
rect 7607 19468 7932 19496
rect 7607 19465 7619 19468
rect 7561 19459 7619 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 9398 19456 9404 19508
rect 9456 19496 9462 19508
rect 9585 19499 9643 19505
rect 9585 19496 9597 19499
rect 9456 19468 9597 19496
rect 9456 19456 9462 19468
rect 9585 19465 9597 19468
rect 9631 19465 9643 19499
rect 10502 19496 10508 19508
rect 10463 19468 10508 19496
rect 9585 19459 9643 19465
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 11514 19456 11520 19508
rect 11572 19496 11578 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11572 19468 11713 19496
rect 11572 19456 11578 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 15378 19496 15384 19508
rect 15339 19468 15384 19496
rect 11701 19459 11759 19465
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 21082 19456 21088 19508
rect 21140 19496 21146 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 21140 19468 21373 19496
rect 21140 19456 21146 19468
rect 21361 19465 21373 19468
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 4522 19388 4528 19440
rect 4580 19428 4586 19440
rect 5537 19431 5595 19437
rect 5537 19428 5549 19431
rect 4580 19400 5549 19428
rect 4580 19388 4586 19400
rect 5537 19397 5549 19400
rect 5583 19397 5595 19431
rect 5537 19391 5595 19397
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 8110 19428 8116 19440
rect 6687 19400 8116 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 8110 19388 8116 19400
rect 8168 19388 8174 19440
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 2041 19363 2099 19369
rect 2041 19360 2053 19363
rect 2004 19332 2053 19360
rect 2004 19320 2010 19332
rect 2041 19329 2053 19332
rect 2087 19329 2099 19363
rect 5074 19360 5080 19372
rect 5035 19332 5080 19360
rect 2041 19323 2099 19329
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12768 19332 12817 19360
rect 12768 19320 12774 19332
rect 12805 19329 12817 19332
rect 12851 19360 12863 19363
rect 16945 19363 17003 19369
rect 12851 19332 13952 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 13924 19304 13952 19332
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17770 19360 17776 19372
rect 16991 19332 17776 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19116 19332 19288 19360
rect 19116 19320 19122 19332
rect 2308 19295 2366 19301
rect 2308 19261 2320 19295
rect 2354 19292 2366 19295
rect 2682 19292 2688 19304
rect 2354 19264 2688 19292
rect 2354 19261 2366 19264
rect 2308 19255 2366 19261
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 4599 19295 4657 19301
rect 4599 19261 4611 19295
rect 4645 19292 4657 19295
rect 5442 19292 5448 19304
rect 4645 19264 5448 19292
rect 4645 19261 4657 19264
rect 4599 19255 4657 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 10134 19292 10140 19304
rect 10095 19264 10140 19292
rect 8205 19255 8263 19261
rect 5166 19224 5172 19236
rect 5079 19196 5172 19224
rect 5166 19184 5172 19196
rect 5224 19224 5230 19236
rect 5994 19224 6000 19236
rect 5224 19196 6000 19224
rect 5224 19184 5230 19196
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 6825 19227 6883 19233
rect 6825 19193 6837 19227
rect 6871 19224 6883 19227
rect 7190 19224 7196 19236
rect 6871 19196 7196 19224
rect 6871 19193 6883 19196
rect 6825 19187 6883 19193
rect 7190 19184 7196 19196
rect 7248 19184 7254 19236
rect 1854 19156 1860 19168
rect 1815 19128 1860 19156
rect 1854 19116 1860 19128
rect 1912 19116 1918 19168
rect 3421 19159 3479 19165
rect 3421 19125 3433 19159
rect 3467 19156 3479 19159
rect 3786 19156 3792 19168
rect 3467 19128 3792 19156
rect 3467 19125 3479 19128
rect 3421 19119 3479 19125
rect 3786 19116 3792 19128
rect 3844 19116 3850 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 4212 19128 4353 19156
rect 4212 19116 4218 19128
rect 4341 19125 4353 19128
rect 4387 19156 4399 19159
rect 5077 19159 5135 19165
rect 5077 19156 5089 19159
rect 4387 19128 5089 19156
rect 4387 19125 4399 19128
rect 4341 19119 4399 19125
rect 5077 19125 5089 19128
rect 5123 19125 5135 19159
rect 5077 19119 5135 19125
rect 8113 19159 8171 19165
rect 8113 19125 8125 19159
rect 8159 19156 8171 19159
rect 8220 19156 8248 19255
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 10502 19252 10508 19304
rect 10560 19292 10566 19304
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 10560 19264 11069 19292
rect 10560 19252 10566 19264
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 11330 19292 11336 19304
rect 11243 19264 11336 19292
rect 11057 19255 11115 19261
rect 11330 19252 11336 19264
rect 11388 19292 11394 19304
rect 12342 19292 12348 19304
rect 11388 19264 12348 19292
rect 11388 19252 11394 19264
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12986 19292 12992 19304
rect 12947 19264 12992 19292
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13722 19292 13728 19304
rect 13587 19264 13728 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13906 19292 13912 19304
rect 13819 19264 13912 19292
rect 13906 19252 13912 19264
rect 13964 19292 13970 19304
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13964 19264 14013 19292
rect 13964 19252 13970 19264
rect 14001 19261 14013 19264
rect 14047 19292 14059 19295
rect 16574 19292 16580 19304
rect 14047 19264 16252 19292
rect 16535 19264 16580 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 8450 19227 8508 19233
rect 8450 19224 8462 19227
rect 8352 19196 8462 19224
rect 8352 19184 8358 19196
rect 8450 19193 8462 19196
rect 8496 19193 8508 19227
rect 10152 19224 10180 19252
rect 11241 19227 11299 19233
rect 11241 19224 11253 19227
rect 10152 19196 11253 19224
rect 8450 19187 8508 19193
rect 11241 19193 11253 19196
rect 11287 19193 11299 19227
rect 13740 19224 13768 19252
rect 16224 19236 16252 19264
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 14246 19227 14304 19233
rect 14246 19224 14258 19227
rect 13740 19196 14258 19224
rect 11241 19187 11299 19193
rect 14246 19193 14258 19196
rect 14292 19193 14304 19227
rect 14246 19187 14304 19193
rect 16206 19184 16212 19236
rect 16264 19224 16270 19236
rect 16301 19227 16359 19233
rect 16301 19224 16313 19227
rect 16264 19196 16313 19224
rect 16264 19184 16270 19196
rect 16301 19193 16313 19196
rect 16347 19224 16359 19227
rect 17770 19224 17776 19236
rect 16347 19196 17776 19224
rect 16347 19193 16359 19196
rect 16301 19187 16359 19193
rect 17770 19184 17776 19196
rect 17828 19224 17834 19236
rect 17865 19227 17923 19233
rect 17865 19224 17877 19227
rect 17828 19196 17877 19224
rect 17828 19184 17834 19196
rect 17865 19193 17877 19196
rect 17911 19224 17923 19227
rect 18064 19224 18092 19255
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18305 19295 18363 19301
rect 18305 19292 18317 19295
rect 18196 19264 18317 19292
rect 18196 19252 18202 19264
rect 18305 19261 18317 19264
rect 18351 19261 18363 19295
rect 19260 19292 19288 19332
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19260 19264 19993 19292
rect 18305 19255 18363 19261
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 20625 19295 20683 19301
rect 20625 19292 20637 19295
rect 19981 19255 20039 19261
rect 20456 19264 20637 19292
rect 18414 19224 18420 19236
rect 17911 19196 18420 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 18414 19184 18420 19196
rect 18472 19184 18478 19236
rect 20456 19168 20484 19264
rect 20625 19261 20637 19264
rect 20671 19261 20683 19295
rect 20625 19255 20683 19261
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 21913 19295 21971 19301
rect 21913 19292 21925 19295
rect 20947 19264 21925 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 21913 19261 21925 19264
rect 21959 19292 21971 19295
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 21959 19264 22477 19292
rect 21959 19261 21971 19264
rect 21913 19255 21971 19261
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 9490 19156 9496 19168
rect 8159 19128 9496 19156
rect 8159 19125 8171 19128
rect 8113 19119 8171 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10771 19159 10829 19165
rect 10771 19125 10783 19159
rect 10817 19156 10829 19159
rect 10962 19156 10968 19168
rect 10817 19128 10968 19156
rect 10817 19125 10829 19128
rect 10771 19119 10829 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 12158 19156 12164 19168
rect 12119 19128 12164 19156
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 18690 19116 18696 19168
rect 18748 19156 18754 19168
rect 19429 19159 19487 19165
rect 19429 19156 19441 19159
rect 18748 19128 19441 19156
rect 18748 19116 18754 19128
rect 19429 19125 19441 19128
rect 19475 19125 19487 19159
rect 20438 19156 20444 19168
rect 20399 19128 20444 19156
rect 19429 19119 19487 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 22097 19159 22155 19165
rect 22097 19125 22109 19159
rect 22143 19156 22155 19159
rect 22186 19156 22192 19168
rect 22143 19128 22192 19156
rect 22143 19125 22155 19128
rect 22097 19119 22155 19125
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 22830 19156 22836 19168
rect 22791 19128 22836 19156
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2590 18952 2596 18964
rect 2551 18924 2596 18952
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 5721 18955 5779 18961
rect 5721 18952 5733 18955
rect 5592 18924 5733 18952
rect 5592 18912 5598 18924
rect 5721 18921 5733 18924
rect 5767 18952 5779 18955
rect 6362 18952 6368 18964
rect 5767 18924 6368 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8260 18924 8309 18952
rect 8260 18912 8266 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 8297 18915 8355 18921
rect 10781 18955 10839 18961
rect 10781 18921 10793 18955
rect 10827 18952 10839 18955
rect 11330 18952 11336 18964
rect 10827 18924 11336 18952
rect 10827 18921 10839 18924
rect 10781 18915 10839 18921
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 11609 18955 11667 18961
rect 11609 18921 11621 18955
rect 11655 18952 11667 18955
rect 12158 18952 12164 18964
rect 11655 18924 12164 18952
rect 11655 18921 11667 18924
rect 11609 18915 11667 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 19150 18952 19156 18964
rect 19111 18924 19156 18952
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 22922 18952 22928 18964
rect 22883 18924 22928 18952
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 1578 18844 1584 18896
rect 1636 18884 1642 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 1636 18856 2421 18884
rect 1636 18844 1642 18856
rect 2409 18853 2421 18856
rect 2455 18884 2467 18887
rect 2682 18884 2688 18896
rect 2455 18856 2688 18884
rect 2455 18853 2467 18856
rect 2409 18847 2467 18853
rect 2682 18844 2688 18856
rect 2740 18844 2746 18896
rect 4614 18893 4620 18896
rect 4608 18884 4620 18893
rect 4575 18856 4620 18884
rect 4608 18847 4620 18856
rect 4614 18844 4620 18847
rect 4672 18844 4678 18896
rect 7377 18887 7435 18893
rect 7377 18853 7389 18887
rect 7423 18884 7435 18887
rect 7926 18884 7932 18896
rect 7423 18856 7932 18884
rect 7423 18853 7435 18856
rect 7377 18847 7435 18853
rect 7926 18844 7932 18856
rect 7984 18844 7990 18896
rect 10229 18887 10287 18893
rect 10229 18853 10241 18887
rect 10275 18853 10287 18887
rect 10229 18847 10287 18853
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 11698 18884 11704 18896
rect 11287 18856 11704 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18816 1731 18819
rect 2038 18816 2044 18828
rect 1719 18788 2044 18816
rect 1719 18785 1731 18788
rect 1673 18779 1731 18785
rect 2038 18776 2044 18788
rect 2096 18816 2102 18828
rect 2866 18816 2872 18828
rect 2096 18788 2872 18816
rect 2096 18776 2102 18788
rect 2866 18776 2872 18788
rect 2924 18816 2930 18828
rect 3234 18816 3240 18828
rect 2924 18788 3240 18816
rect 2924 18776 2930 18788
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18816 4399 18819
rect 4982 18816 4988 18828
rect 4387 18788 4988 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 7190 18816 7196 18828
rect 7151 18788 7196 18816
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 9030 18816 9036 18828
rect 8619 18788 9036 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 9030 18776 9036 18788
rect 9088 18816 9094 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9088 18788 10057 18816
rect 9088 18776 9094 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18748 2743 18751
rect 3786 18748 3792 18760
rect 2731 18720 3792 18748
rect 2731 18717 2743 18720
rect 2685 18711 2743 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 7466 18748 7472 18760
rect 7427 18720 7472 18748
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 2130 18680 2136 18692
rect 2091 18652 2136 18680
rect 2130 18640 2136 18652
rect 2188 18640 2194 18692
rect 6914 18680 6920 18692
rect 6875 18652 6920 18680
rect 6914 18640 6920 18652
rect 6972 18640 6978 18692
rect 9766 18680 9772 18692
rect 9727 18652 9772 18680
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 3142 18612 3148 18624
rect 3103 18584 3148 18612
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3292 18584 3433 18612
rect 3292 18572 3298 18584
rect 3421 18581 3433 18584
rect 3467 18581 3479 18615
rect 3786 18612 3792 18624
rect 3747 18584 3792 18612
rect 3421 18575 3479 18581
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 6052 18584 6285 18612
rect 6052 18572 6058 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6730 18612 6736 18624
rect 6691 18584 6736 18612
rect 6273 18575 6331 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 7650 18572 7656 18624
rect 7708 18612 7714 18624
rect 7929 18615 7987 18621
rect 7929 18612 7941 18615
rect 7708 18584 7941 18612
rect 7708 18572 7714 18584
rect 7929 18581 7941 18584
rect 7975 18612 7987 18615
rect 8110 18612 8116 18624
rect 7975 18584 8116 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 8352 18584 9413 18612
rect 8352 18572 8358 18584
rect 9401 18581 9413 18584
rect 9447 18612 9459 18615
rect 10244 18612 10272 18847
rect 11698 18844 11704 18856
rect 11756 18884 11762 18896
rect 12250 18884 12256 18896
rect 11756 18856 12256 18884
rect 11756 18844 11762 18856
rect 12250 18844 12256 18856
rect 12308 18884 12314 18896
rect 12345 18887 12403 18893
rect 12345 18884 12357 18887
rect 12308 18856 12357 18884
rect 12308 18844 12314 18856
rect 12345 18853 12357 18856
rect 12391 18853 12403 18887
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 12345 18847 12403 18853
rect 13096 18856 13277 18884
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11848 18788 12173 18816
rect 11848 18776 11854 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 11054 18748 11060 18760
rect 10367 18720 11060 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12492 18720 12537 18748
rect 12492 18708 12498 18720
rect 11885 18683 11943 18689
rect 11885 18649 11897 18683
rect 11931 18680 11943 18683
rect 13096 18680 13124 18856
rect 13265 18853 13277 18856
rect 13311 18884 13323 18887
rect 13909 18887 13967 18893
rect 13909 18884 13921 18887
rect 13311 18856 13921 18884
rect 13311 18853 13323 18856
rect 13265 18847 13323 18853
rect 13909 18853 13921 18856
rect 13955 18853 13967 18887
rect 13909 18847 13967 18853
rect 15286 18844 15292 18896
rect 15344 18884 15350 18896
rect 15841 18887 15899 18893
rect 15841 18884 15853 18887
rect 15344 18856 15853 18884
rect 15344 18844 15350 18856
rect 15841 18853 15853 18856
rect 15887 18884 15899 18887
rect 15930 18884 15936 18896
rect 15887 18856 15936 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 18040 18887 18098 18893
rect 18040 18853 18052 18887
rect 18086 18884 18098 18887
rect 18322 18884 18328 18896
rect 18086 18856 18328 18884
rect 18086 18853 18098 18856
rect 18040 18847 18098 18853
rect 18322 18844 18328 18856
rect 18380 18884 18386 18896
rect 18690 18884 18696 18896
rect 18380 18856 18696 18884
rect 18380 18844 18386 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 21177 18887 21235 18893
rect 21177 18884 21189 18887
rect 21140 18856 21189 18884
rect 21140 18844 21146 18856
rect 21177 18853 21189 18856
rect 21223 18853 21235 18887
rect 21177 18847 21235 18853
rect 13170 18776 13176 18828
rect 13228 18816 13234 18828
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 13228 18788 13737 18816
rect 13228 18776 13234 18788
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 15620 18788 15669 18816
rect 15620 18776 15626 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 17770 18816 17776 18828
rect 17731 18788 17776 18816
rect 15657 18779 15715 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 20898 18816 20904 18828
rect 20859 18788 20904 18816
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 22738 18816 22744 18828
rect 22699 18788 22744 18816
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 13998 18748 14004 18760
rect 13959 18720 14004 18748
rect 13998 18708 14004 18720
rect 14056 18748 14062 18760
rect 14369 18751 14427 18757
rect 14369 18748 14381 18751
rect 14056 18720 14381 18748
rect 14056 18708 14062 18720
rect 14369 18717 14381 18720
rect 14415 18717 14427 18751
rect 14369 18711 14427 18717
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15344 18720 15945 18748
rect 15344 18708 15350 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 11931 18652 13124 18680
rect 15381 18683 15439 18689
rect 11931 18649 11943 18652
rect 11885 18643 11943 18649
rect 15381 18649 15393 18683
rect 15427 18680 15439 18683
rect 16666 18680 16672 18692
rect 15427 18652 16672 18680
rect 15427 18649 15439 18652
rect 15381 18643 15439 18649
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 13446 18612 13452 18624
rect 9447 18584 10272 18612
rect 13407 18584 13452 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 4525 18411 4583 18417
rect 4525 18377 4537 18411
rect 4571 18408 4583 18411
rect 4614 18408 4620 18420
rect 4571 18380 4620 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 4614 18368 4620 18380
rect 4672 18408 4678 18420
rect 5258 18408 5264 18420
rect 4672 18380 5264 18408
rect 4672 18368 4678 18380
rect 5258 18368 5264 18380
rect 5316 18408 5322 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 5316 18380 5549 18408
rect 5316 18368 5322 18380
rect 5537 18377 5549 18380
rect 5583 18408 5595 18411
rect 5994 18408 6000 18420
rect 5583 18380 6000 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6273 18411 6331 18417
rect 6273 18377 6285 18411
rect 6319 18408 6331 18411
rect 7190 18408 7196 18420
rect 6319 18380 7196 18408
rect 6319 18377 6331 18380
rect 6273 18371 6331 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 13170 18408 13176 18420
rect 12636 18380 13176 18408
rect 1489 18343 1547 18349
rect 1489 18309 1501 18343
rect 1535 18309 1547 18343
rect 1489 18303 1547 18309
rect 1504 18204 1532 18303
rect 1946 18300 1952 18352
rect 2004 18340 2010 18352
rect 2004 18312 2544 18340
rect 2004 18300 2010 18312
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2516 18281 2544 18312
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 2547 18244 3096 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2958 18204 2964 18216
rect 1504 18176 2964 18204
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 3068 18213 3096 18244
rect 5074 18232 5080 18284
rect 5132 18272 5138 18284
rect 12636 18281 12664 18380
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 13541 18411 13599 18417
rect 13541 18377 13553 18411
rect 13587 18408 13599 18411
rect 13906 18408 13912 18420
rect 13587 18380 13912 18408
rect 13587 18377 13599 18380
rect 13541 18371 13599 18377
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5132 18244 5641 18272
rect 5132 18232 5138 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18241 12679 18275
rect 12621 18235 12679 18241
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13648 18281 13676 18380
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15286 18408 15292 18420
rect 15059 18380 15292 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 15930 18408 15936 18420
rect 15891 18380 15936 18408
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16206 18408 16212 18420
rect 16167 18380 16212 18408
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 17770 18408 17776 18420
rect 17731 18380 17776 18408
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 18322 18408 18328 18420
rect 18283 18380 18328 18408
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 20898 18408 20904 18420
rect 20859 18380 20904 18408
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 13044 18244 13645 18272
rect 13044 18232 13050 18244
rect 13633 18241 13645 18244
rect 13679 18241 13691 18275
rect 13633 18235 13691 18241
rect 21545 18275 21603 18281
rect 21545 18241 21557 18275
rect 21591 18272 21603 18275
rect 22830 18272 22836 18284
rect 21591 18244 22836 18272
rect 21591 18241 21603 18244
rect 21545 18235 21603 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18204 3111 18207
rect 3142 18204 3148 18216
rect 3099 18176 3148 18204
rect 3099 18173 3111 18176
rect 3053 18167 3111 18173
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 6638 18204 6644 18216
rect 6551 18176 6644 18204
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 3234 18136 3240 18148
rect 1811 18108 3240 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 3234 18096 3240 18108
rect 3292 18096 3298 18148
rect 3412 18139 3470 18145
rect 3412 18105 3424 18139
rect 3458 18136 3470 18139
rect 3786 18136 3792 18148
rect 3458 18108 3792 18136
rect 3458 18105 3470 18108
rect 3412 18099 3470 18105
rect 3786 18096 3792 18108
rect 3844 18136 3850 18148
rect 4154 18136 4160 18148
rect 3844 18108 4160 18136
rect 3844 18096 3850 18108
rect 4154 18096 4160 18108
rect 4212 18096 4218 18148
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 1949 18071 2007 18077
rect 1949 18068 1961 18071
rect 1912 18040 1961 18068
rect 1912 18028 1918 18040
rect 1949 18037 1961 18040
rect 1995 18037 2007 18071
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 1949 18031 2007 18037
rect 5074 18028 5080 18040
rect 5132 18068 5138 18080
rect 6564 18077 6592 18176
rect 6638 18164 6644 18176
rect 6696 18204 6702 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6696 18176 6837 18204
rect 6696 18164 6702 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18173 9551 18207
rect 21266 18204 21272 18216
rect 21227 18176 21272 18204
rect 9493 18167 9551 18173
rect 6730 18096 6736 18148
rect 6788 18136 6794 18148
rect 7070 18139 7128 18145
rect 7070 18136 7082 18139
rect 6788 18108 7082 18136
rect 6788 18096 6794 18108
rect 7070 18105 7082 18108
rect 7116 18105 7128 18139
rect 7070 18099 7128 18105
rect 9508 18080 9536 18167
rect 21266 18164 21272 18176
rect 21324 18204 21330 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21324 18176 22017 18204
rect 21324 18164 21330 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 9582 18096 9588 18148
rect 9640 18136 9646 18148
rect 9760 18139 9818 18145
rect 9760 18136 9772 18139
rect 9640 18108 9772 18136
rect 9640 18096 9646 18108
rect 9760 18105 9772 18108
rect 9806 18136 9818 18139
rect 13900 18139 13958 18145
rect 9806 18108 11100 18136
rect 9806 18105 9818 18108
rect 9760 18099 9818 18105
rect 11072 18080 11100 18108
rect 13900 18105 13912 18139
rect 13946 18136 13958 18139
rect 13998 18136 14004 18148
rect 13946 18108 14004 18136
rect 13946 18105 13958 18108
rect 13900 18099 13958 18105
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 16298 18136 16304 18148
rect 15344 18108 16304 18136
rect 15344 18096 15350 18108
rect 16298 18096 16304 18108
rect 16356 18136 16362 18148
rect 16485 18139 16543 18145
rect 16485 18136 16497 18139
rect 16356 18108 16497 18136
rect 16356 18096 16362 18108
rect 16485 18105 16497 18108
rect 16531 18105 16543 18139
rect 16666 18136 16672 18148
rect 16627 18108 16672 18136
rect 16485 18099 16543 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 16758 18096 16764 18148
rect 16816 18136 16822 18148
rect 17129 18139 17187 18145
rect 17129 18136 17141 18139
rect 16816 18108 17141 18136
rect 16816 18096 16822 18108
rect 17129 18105 17141 18108
rect 17175 18105 17187 18139
rect 17129 18099 17187 18105
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 5132 18040 6561 18068
rect 5132 18028 5138 18040
rect 6549 18037 6561 18040
rect 6595 18037 6607 18071
rect 6549 18031 6607 18037
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 7524 18040 8217 18068
rect 7524 18028 7530 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8205 18031 8263 18037
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9490 18068 9496 18080
rect 9447 18040 9496 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 10870 18068 10876 18080
rect 10831 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11425 18071 11483 18077
rect 11425 18068 11437 18071
rect 11112 18040 11437 18068
rect 11112 18028 11118 18040
rect 11425 18037 11437 18040
rect 11471 18037 11483 18071
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11425 18031 11483 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 15562 18068 15568 18080
rect 15523 18040 15568 18068
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22738 18068 22744 18080
rect 22152 18040 22744 18068
rect 22152 18028 22158 18040
rect 22738 18028 22744 18040
rect 22796 18028 22802 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 2832 17836 3341 17864
rect 2832 17824 2838 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4212 17836 4813 17864
rect 4212 17824 4218 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 4801 17827 4859 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6730 17864 6736 17876
rect 6691 17836 6736 17864
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17864 7530 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7524 17836 7665 17864
rect 7524 17824 7530 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 9122 17864 9128 17876
rect 8435 17836 9128 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 1946 17796 1952 17808
rect 1412 17768 1952 17796
rect 1412 17737 1440 17768
rect 1946 17756 1952 17768
rect 2004 17756 2010 17808
rect 2958 17756 2964 17808
rect 3016 17796 3022 17808
rect 4341 17799 4399 17805
rect 3016 17768 4108 17796
rect 3016 17756 3022 17768
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1397 17691 1455 17697
rect 1664 17731 1722 17737
rect 1664 17697 1676 17731
rect 1710 17728 1722 17731
rect 2406 17728 2412 17740
rect 1710 17700 2412 17728
rect 1710 17697 1722 17700
rect 1664 17691 1722 17697
rect 2406 17688 2412 17700
rect 2464 17728 2470 17740
rect 4080 17737 4108 17768
rect 4341 17765 4353 17799
rect 4387 17796 4399 17799
rect 5350 17796 5356 17808
rect 4387 17768 5356 17796
rect 4387 17765 4399 17768
rect 4341 17759 4399 17765
rect 5350 17756 5356 17768
rect 5408 17756 5414 17808
rect 5534 17756 5540 17808
rect 5592 17805 5598 17808
rect 5592 17799 5656 17805
rect 5592 17765 5610 17799
rect 5644 17765 5656 17799
rect 5592 17759 5656 17765
rect 5592 17756 5598 17759
rect 7006 17756 7012 17808
rect 7064 17796 7070 17808
rect 8404 17796 8432 17827
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 9582 17864 9588 17876
rect 9539 17836 9588 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11885 17867 11943 17873
rect 11885 17833 11897 17867
rect 11931 17864 11943 17867
rect 12434 17864 12440 17876
rect 11931 17836 12440 17864
rect 11931 17833 11943 17836
rect 11885 17827 11943 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 14642 17824 14648 17876
rect 14700 17864 14706 17876
rect 15105 17867 15163 17873
rect 15105 17864 15117 17867
rect 14700 17836 15117 17864
rect 14700 17824 14706 17836
rect 15105 17833 15117 17836
rect 15151 17864 15163 17867
rect 15194 17864 15200 17876
rect 15151 17836 15200 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 16669 17867 16727 17873
rect 16669 17833 16681 17867
rect 16715 17864 16727 17867
rect 16758 17864 16764 17876
rect 16715 17836 16764 17864
rect 16715 17833 16727 17836
rect 16669 17827 16727 17833
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 7064 17768 8432 17796
rect 15212 17796 15240 17824
rect 15534 17799 15592 17805
rect 15534 17796 15546 17799
rect 15212 17768 15546 17796
rect 7064 17756 7070 17768
rect 15534 17765 15546 17768
rect 15580 17765 15592 17799
rect 22002 17796 22008 17808
rect 21963 17768 22008 17796
rect 15534 17759 15592 17765
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 3697 17731 3755 17737
rect 3697 17728 3709 17731
rect 2464 17700 3709 17728
rect 2464 17688 2470 17700
rect 3697 17697 3709 17700
rect 3743 17697 3755 17731
rect 3697 17691 3755 17697
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 6454 17728 6460 17740
rect 4111 17700 6460 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 8481 17731 8539 17737
rect 8481 17728 8493 17731
rect 6788 17700 8493 17728
rect 6788 17688 6794 17700
rect 8481 17697 8493 17700
rect 8527 17697 8539 17731
rect 8481 17691 8539 17697
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 9950 17737 9956 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9640 17700 9689 17728
rect 9640 17688 9646 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9944 17728 9956 17737
rect 9911 17700 9956 17728
rect 9677 17691 9735 17697
rect 9944 17691 9956 17700
rect 9950 17688 9956 17691
rect 10008 17688 10014 17740
rect 11514 17688 11520 17740
rect 11572 17728 11578 17740
rect 12417 17731 12475 17737
rect 12417 17728 12429 17731
rect 11572 17700 12429 17728
rect 11572 17688 11578 17700
rect 12417 17697 12429 17700
rect 12463 17697 12475 17731
rect 12417 17691 12475 17697
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 15378 17728 15384 17740
rect 15335 17700 15384 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 15378 17688 15384 17700
rect 15436 17728 15442 17740
rect 16114 17728 16120 17740
rect 15436 17700 16120 17728
rect 15436 17688 15442 17700
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 21726 17728 21732 17740
rect 21687 17700 21732 17728
rect 21726 17688 21732 17700
rect 21784 17688 21790 17740
rect 5074 17620 5080 17672
rect 5132 17660 5138 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 5132 17632 5365 17660
rect 5132 17620 5138 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7432 17632 8309 17660
rect 7432 17620 7438 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 8297 17623 8355 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 17770 17660 17776 17672
rect 17731 17632 17776 17660
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 2777 17595 2835 17601
rect 2777 17561 2789 17595
rect 2823 17592 2835 17595
rect 2866 17592 2872 17604
rect 2823 17564 2872 17592
rect 2823 17561 2835 17564
rect 2777 17555 2835 17561
rect 2866 17552 2872 17564
rect 2924 17552 2930 17604
rect 7926 17592 7932 17604
rect 7887 17564 7932 17592
rect 7926 17552 7932 17564
rect 7984 17592 7990 17604
rect 8849 17595 8907 17601
rect 8849 17592 8861 17595
rect 7984 17564 8861 17592
rect 7984 17552 7990 17564
rect 8849 17561 8861 17564
rect 8895 17561 8907 17595
rect 8849 17555 8907 17561
rect 13538 17524 13544 17536
rect 13499 17496 13544 17524
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 14056 17496 14105 17524
rect 14056 17484 14062 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14093 17487 14151 17493
rect 18325 17527 18383 17533
rect 18325 17493 18337 17527
rect 18371 17524 18383 17527
rect 18598 17524 18604 17536
rect 18371 17496 18604 17524
rect 18371 17493 18383 17496
rect 18325 17487 18383 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 3142 17280 3148 17332
rect 3200 17320 3206 17332
rect 3237 17323 3295 17329
rect 3237 17320 3249 17323
rect 3200 17292 3249 17320
rect 3200 17280 3206 17292
rect 3237 17289 3249 17292
rect 3283 17320 3295 17323
rect 5074 17320 5080 17332
rect 3283 17292 5080 17320
rect 3283 17289 3295 17292
rect 3237 17283 3295 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5592 17292 5733 17320
rect 5592 17280 5598 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 6454 17320 6460 17332
rect 6415 17292 6460 17320
rect 5721 17283 5779 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 7006 17320 7012 17332
rect 6967 17292 7012 17320
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7834 17320 7840 17332
rect 7156 17292 7840 17320
rect 7156 17280 7162 17292
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 10870 17320 10876 17332
rect 10704 17292 10876 17320
rect 1854 17252 1860 17264
rect 1815 17224 1860 17252
rect 1854 17212 1860 17224
rect 1912 17212 1918 17264
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 4433 17255 4491 17261
rect 4433 17252 4445 17255
rect 4212 17224 4445 17252
rect 4212 17212 4218 17224
rect 4433 17221 4445 17224
rect 4479 17252 4491 17255
rect 5442 17252 5448 17264
rect 4479 17224 5448 17252
rect 4479 17221 4491 17224
rect 4433 17215 4491 17221
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 10134 17252 10140 17264
rect 10095 17224 10140 17252
rect 10134 17212 10140 17224
rect 10192 17212 10198 17264
rect 2406 17184 2412 17196
rect 2367 17156 2412 17184
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 3329 17187 3387 17193
rect 3329 17184 3341 17187
rect 3292 17156 3341 17184
rect 3292 17144 3298 17156
rect 3329 17153 3341 17156
rect 3375 17153 3387 17187
rect 6638 17184 6644 17196
rect 3329 17147 3387 17153
rect 3804 17156 6644 17184
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2869 17119 2927 17125
rect 1719 17088 2360 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2332 17060 2360 17088
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3694 17116 3700 17128
rect 2915 17088 3700 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 2133 17051 2191 17057
rect 2133 17017 2145 17051
rect 2179 17017 2191 17051
rect 2314 17048 2320 17060
rect 2275 17020 2320 17048
rect 2133 17011 2191 17017
rect 2148 16980 2176 17011
rect 2314 17008 2320 17020
rect 2372 17008 2378 17060
rect 2884 16980 2912 17079
rect 3694 17076 3700 17088
rect 3752 17116 3758 17128
rect 3804 17116 3832 17156
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 9582 17184 9588 17196
rect 9495 17156 9588 17184
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 3752 17088 3832 17116
rect 3896 17088 4997 17116
rect 3752 17076 3758 17088
rect 3896 16992 3924 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 7374 17116 7380 17128
rect 5316 17088 7380 17116
rect 5316 17076 5322 17088
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7558 17116 7564 17128
rect 7519 17088 7564 17116
rect 7558 17076 7564 17088
rect 7616 17116 7622 17128
rect 9508 17125 9536 17156
rect 9582 17144 9588 17156
rect 9640 17184 9646 17196
rect 10704 17193 10732 17292
rect 10870 17280 10876 17292
rect 10928 17320 10934 17332
rect 11149 17323 11207 17329
rect 11149 17320 11161 17323
rect 10928 17292 11161 17320
rect 10928 17280 10934 17292
rect 11149 17289 11161 17292
rect 11195 17320 11207 17323
rect 11514 17320 11520 17332
rect 11195 17292 11520 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 13630 17320 13636 17332
rect 12860 17292 13636 17320
rect 12860 17280 12866 17292
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 14642 17320 14648 17332
rect 14603 17292 14648 17320
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15013 17323 15071 17329
rect 15013 17289 15025 17323
rect 15059 17320 15071 17323
rect 15378 17320 15384 17332
rect 15059 17292 15384 17320
rect 15059 17289 15071 17292
rect 15013 17283 15071 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17320 17834 17332
rect 21726 17320 21732 17332
rect 17828 17292 18552 17320
rect 21687 17292 21732 17320
rect 17828 17280 17834 17292
rect 10689 17187 10747 17193
rect 9640 17156 10640 17184
rect 9640 17144 9646 17156
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 7616 17088 9505 17116
rect 7616 17076 7622 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 10612 17116 10640 17156
rect 10689 17153 10701 17187
rect 10735 17153 10747 17187
rect 15396 17184 15424 17280
rect 18138 17252 18144 17264
rect 18099 17224 18144 17252
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 18524 17193 18552 17292
rect 21726 17280 21732 17292
rect 21784 17280 21790 17332
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 15396 17156 15485 17184
rect 10689 17147 10747 17153
rect 15473 17153 15485 17156
rect 15519 17153 15531 17187
rect 15473 17147 15531 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17153 18567 17187
rect 18509 17147 18567 17153
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 9916 17088 10548 17116
rect 10612 17088 11805 17116
rect 9916 17076 9922 17088
rect 4706 17048 4712 17060
rect 4667 17020 4712 17048
rect 4706 17008 4712 17020
rect 4764 17008 4770 17060
rect 4890 17048 4896 17060
rect 4851 17020 4896 17048
rect 4890 17008 4896 17020
rect 4948 17008 4954 17060
rect 6086 17048 6092 17060
rect 6047 17020 6092 17048
rect 6086 17008 6092 17020
rect 6144 17008 6150 17060
rect 7466 17008 7472 17060
rect 7524 17048 7530 17060
rect 7806 17051 7864 17057
rect 7806 17048 7818 17051
rect 7524 17020 7818 17048
rect 7524 17008 7530 17020
rect 7806 17017 7818 17020
rect 7852 17017 7864 17051
rect 7806 17011 7864 17017
rect 10413 17051 10471 17057
rect 10413 17017 10425 17051
rect 10459 17017 10471 17051
rect 10520 17048 10548 17088
rect 11793 17085 11805 17088
rect 11839 17116 11851 17119
rect 12158 17116 12164 17128
rect 11839 17088 12164 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 12158 17076 12164 17088
rect 12216 17116 12222 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12216 17088 12449 17116
rect 12216 17076 12222 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 12704 17119 12762 17125
rect 12704 17116 12716 17119
rect 12584 17088 12716 17116
rect 12584 17076 12590 17088
rect 12704 17085 12716 17088
rect 12750 17116 12762 17119
rect 13538 17116 13544 17128
rect 12750 17088 13544 17116
rect 12750 17085 12762 17088
rect 12704 17079 12762 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 15746 17125 15752 17128
rect 15740 17116 15752 17125
rect 15659 17088 15752 17116
rect 15740 17079 15752 17088
rect 15804 17116 15810 17128
rect 16758 17116 16764 17128
rect 15804 17088 16764 17116
rect 15746 17076 15752 17079
rect 15804 17076 15810 17088
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 10520 17020 10609 17048
rect 10413 17011 10471 17017
rect 10597 17017 10609 17020
rect 10643 17017 10655 17051
rect 18693 17051 18751 17057
rect 18693 17048 18705 17051
rect 10597 17011 10655 17017
rect 17420 17020 18705 17048
rect 3878 16980 3884 16992
rect 2148 16952 2912 16980
rect 3839 16952 3884 16980
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4908 16980 4936 17008
rect 4295 16952 4936 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 5074 16940 5080 16992
rect 5132 16980 5138 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 5132 16952 5365 16980
rect 5132 16940 5138 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8941 16983 8999 16989
rect 8941 16980 8953 16983
rect 8352 16952 8953 16980
rect 8352 16940 8358 16952
rect 8941 16949 8953 16952
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 9861 16983 9919 16989
rect 9861 16980 9873 16983
rect 9824 16952 9873 16980
rect 9824 16940 9830 16952
rect 9861 16949 9873 16952
rect 9907 16980 9919 16983
rect 10428 16980 10456 17011
rect 17420 16992 17448 17020
rect 18693 17017 18705 17020
rect 18739 17017 18751 17051
rect 18693 17011 18751 17017
rect 9907 16952 10456 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 12492 16952 13829 16980
rect 12492 16940 12498 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 16850 16980 16856 16992
rect 16811 16952 16856 16980
rect 13817 16943 13875 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 17402 16980 17408 16992
rect 17363 16952 17408 16980
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 18598 16980 18604 16992
rect 18559 16952 18604 16980
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2406 16736 2412 16788
rect 2464 16776 2470 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2464 16748 2881 16776
rect 2464 16736 2470 16748
rect 2869 16745 2881 16748
rect 2915 16776 2927 16779
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 2915 16748 3801 16776
rect 2915 16745 2927 16748
rect 2869 16739 2927 16745
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 6788 16748 7205 16776
rect 6788 16736 6794 16748
rect 7193 16745 7205 16748
rect 7239 16745 7251 16779
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7193 16739 7251 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8011 16779 8069 16785
rect 8011 16745 8023 16779
rect 8057 16776 8069 16779
rect 8202 16776 8208 16788
rect 8057 16748 8208 16776
rect 8057 16745 8069 16748
rect 8011 16739 8069 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 9916 16748 10057 16776
rect 9916 16736 9922 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10045 16739 10103 16745
rect 10863 16779 10921 16785
rect 10863 16745 10875 16779
rect 10909 16776 10921 16779
rect 10962 16776 10968 16788
rect 10909 16748 10968 16776
rect 10909 16745 10921 16748
rect 10863 16739 10921 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11606 16776 11612 16788
rect 11440 16748 11612 16776
rect 3326 16668 3332 16720
rect 3384 16708 3390 16720
rect 4341 16711 4399 16717
rect 4341 16708 4353 16711
rect 3384 16680 4353 16708
rect 3384 16668 3390 16680
rect 4341 16677 4353 16680
rect 4387 16708 4399 16711
rect 4706 16708 4712 16720
rect 4387 16680 4712 16708
rect 4387 16677 4399 16680
rect 4341 16671 4399 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 8110 16668 8116 16720
rect 8168 16708 8174 16720
rect 8478 16708 8484 16720
rect 8168 16680 8484 16708
rect 8168 16668 8174 16680
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 8588 16680 9812 16708
rect 1756 16643 1814 16649
rect 1756 16609 1768 16643
rect 1802 16640 1814 16643
rect 2590 16640 2596 16652
rect 1802 16612 2596 16640
rect 1802 16609 1814 16612
rect 1756 16603 1814 16609
rect 2590 16600 2596 16612
rect 2648 16640 2654 16652
rect 3421 16643 3479 16649
rect 3421 16640 3433 16643
rect 2648 16612 3433 16640
rect 2648 16600 2654 16612
rect 3421 16609 3433 16612
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 5074 16600 5080 16652
rect 5132 16600 5138 16652
rect 5258 16649 5264 16652
rect 5252 16640 5264 16649
rect 5219 16612 5264 16640
rect 5252 16603 5264 16612
rect 5258 16600 5264 16603
rect 5316 16600 5322 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8588 16649 8616 16680
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8352 16612 8585 16640
rect 8352 16600 8358 16612
rect 8573 16609 8585 16612
rect 8619 16609 8631 16643
rect 8573 16603 8631 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9674 16640 9680 16652
rect 9539 16612 9680 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9784 16640 9812 16680
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 10778 16708 10784 16720
rect 10192 16680 10784 16708
rect 10192 16668 10198 16680
rect 10778 16668 10784 16680
rect 10836 16708 10842 16720
rect 11440 16717 11468 16748
rect 11606 16736 11612 16748
rect 11664 16776 11670 16788
rect 12526 16776 12532 16788
rect 11664 16748 12532 16776
rect 11664 16736 11670 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15746 16776 15752 16788
rect 15707 16748 15752 16776
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17957 16779 18015 16785
rect 17957 16776 17969 16779
rect 17460 16748 17969 16776
rect 17460 16736 17466 16748
rect 17957 16745 17969 16748
rect 18003 16745 18015 16779
rect 17957 16739 18015 16745
rect 11333 16711 11391 16717
rect 11333 16708 11345 16711
rect 10836 16680 11345 16708
rect 10836 16668 10842 16680
rect 11333 16677 11345 16680
rect 11379 16677 11391 16711
rect 11333 16671 11391 16677
rect 11425 16711 11483 16717
rect 11425 16677 11437 16711
rect 11471 16677 11483 16711
rect 11425 16671 11483 16677
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 12866 16711 12924 16717
rect 12866 16708 12878 16711
rect 12492 16680 12878 16708
rect 12492 16668 12498 16680
rect 12866 16677 12878 16680
rect 12912 16677 12924 16711
rect 12866 16671 12924 16677
rect 12986 16668 12992 16720
rect 13044 16668 13050 16720
rect 9950 16640 9956 16652
rect 9784 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10413 16643 10471 16649
rect 10413 16640 10425 16643
rect 10008 16612 10425 16640
rect 10008 16600 10014 16612
rect 10413 16609 10425 16612
rect 10459 16609 10471 16643
rect 11146 16640 11152 16652
rect 11107 16612 11152 16640
rect 10413 16603 10471 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 12158 16600 12164 16652
rect 12216 16640 12222 16652
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12216 16612 12633 16640
rect 12216 16600 12222 16612
rect 12621 16609 12633 16612
rect 12667 16640 12679 16643
rect 13004 16640 13032 16668
rect 12667 16612 13032 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16574 16640 16580 16652
rect 16172 16612 16580 16640
rect 16172 16600 16178 16612
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 16850 16649 16856 16652
rect 16844 16640 16856 16649
rect 16811 16612 16856 16640
rect 16844 16603 16856 16612
rect 16850 16600 16856 16603
rect 16908 16600 16914 16652
rect 1489 16575 1547 16581
rect 1489 16541 1501 16575
rect 1535 16541 1547 16575
rect 1489 16535 1547 16541
rect 1504 16436 1532 16535
rect 4890 16532 4896 16584
rect 4948 16572 4954 16584
rect 4985 16575 5043 16581
rect 4985 16572 4997 16575
rect 4948 16544 4997 16572
rect 4948 16532 4954 16544
rect 4985 16541 4997 16544
rect 5031 16572 5043 16575
rect 5092 16572 5120 16600
rect 8386 16572 8392 16584
rect 5031 16544 5120 16572
rect 8347 16544 8392 16572
rect 5031 16541 5043 16544
rect 4985 16535 5043 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 2130 16436 2136 16448
rect 1504 16408 2136 16436
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4672 16408 4721 16436
rect 4672 16396 4678 16408
rect 4709 16405 4721 16408
rect 4755 16405 4767 16439
rect 6362 16436 6368 16448
rect 6323 16408 6368 16436
rect 4709 16399 4767 16405
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 2188 16204 2237 16232
rect 2188 16192 2194 16204
rect 2225 16201 2237 16204
rect 2271 16232 2283 16235
rect 3142 16232 3148 16244
rect 2271 16204 3148 16232
rect 2271 16201 2283 16204
rect 2225 16195 2283 16201
rect 3142 16192 3148 16204
rect 3200 16192 3206 16244
rect 7745 16235 7803 16241
rect 7745 16201 7757 16235
rect 7791 16232 7803 16235
rect 8202 16232 8208 16244
rect 7791 16204 8208 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8536 16204 8677 16232
rect 8536 16192 8542 16204
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 9582 16232 9588 16244
rect 9543 16204 9588 16232
rect 8665 16195 8723 16201
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 11606 16232 11612 16244
rect 11567 16204 11612 16232
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 12986 16232 12992 16244
rect 12299 16204 12992 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 16022 16232 16028 16244
rect 15983 16204 16028 16232
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 16632 16204 16957 16232
rect 16632 16192 16638 16204
rect 16945 16201 16957 16204
rect 16991 16201 17003 16235
rect 16945 16195 17003 16201
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16164 2835 16167
rect 3973 16167 4031 16173
rect 3973 16164 3985 16167
rect 2823 16136 3985 16164
rect 2823 16133 2835 16136
rect 2777 16127 2835 16133
rect 3973 16133 3985 16136
rect 4019 16133 4031 16167
rect 3973 16127 4031 16133
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2792 16028 2820 16127
rect 5442 16124 5448 16176
rect 5500 16164 5506 16176
rect 6181 16167 6239 16173
rect 6181 16164 6193 16167
rect 5500 16136 6193 16164
rect 5500 16124 5506 16136
rect 6181 16133 6193 16136
rect 6227 16133 6239 16167
rect 6181 16127 6239 16133
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 3878 16096 3884 16108
rect 3835 16068 3884 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 3878 16056 3884 16068
rect 3936 16096 3942 16108
rect 9401 16099 9459 16105
rect 3936 16068 4384 16096
rect 3936 16056 3942 16068
rect 1443 16000 2820 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 4062 15988 4068 16040
rect 4120 15988 4126 16040
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 15997 4307 16031
rect 4356 16028 4384 16068
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10042 16096 10048 16108
rect 9447 16068 10048 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10919 16068 11069 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 11146 16096 11152 16108
rect 11103 16068 11152 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 13004 16096 13032 16192
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 13004 16068 13093 16096
rect 13081 16065 13093 16068
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 16577 16099 16635 16105
rect 16577 16096 16589 16099
rect 15519 16068 16589 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16577 16065 16589 16068
rect 16623 16096 16635 16099
rect 16850 16096 16856 16108
rect 16623 16068 16856 16096
rect 16623 16065 16635 16068
rect 16577 16059 16635 16065
rect 16850 16056 16856 16068
rect 16908 16096 16914 16108
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 16908 16068 17325 16096
rect 16908 16056 16914 16068
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 4516 16031 4574 16037
rect 4516 16028 4528 16031
rect 4356 16000 4528 16028
rect 4249 15991 4307 15997
rect 4516 15997 4528 16000
rect 4562 16028 4574 16031
rect 8662 16028 8668 16040
rect 4562 16000 8668 16028
rect 4562 15997 4574 16000
rect 4516 15991 4574 15997
rect 1673 15963 1731 15969
rect 1673 15929 1685 15963
rect 1719 15960 1731 15963
rect 1946 15960 1952 15972
rect 1719 15932 1952 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 1946 15920 1952 15932
rect 2004 15920 2010 15972
rect 2593 15963 2651 15969
rect 2593 15929 2605 15963
rect 2639 15960 2651 15963
rect 2958 15960 2964 15972
rect 2639 15932 2964 15960
rect 2639 15929 2651 15932
rect 2593 15923 2651 15929
rect 2958 15920 2964 15932
rect 3016 15960 3022 15972
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 3016 15932 3065 15960
rect 3016 15920 3022 15932
rect 3053 15929 3065 15932
rect 3099 15929 3111 15963
rect 3326 15960 3332 15972
rect 3287 15932 3332 15960
rect 3053 15923 3111 15929
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 4080 15960 4108 15988
rect 3620 15932 4108 15960
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3620 15892 3648 15932
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 4264 15960 4292 15991
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 4212 15932 4292 15960
rect 4614 15932 6561 15960
rect 4212 15920 4218 15932
rect 3283 15864 3648 15892
rect 3973 15895 4031 15901
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3973 15861 3985 15895
rect 4019 15892 4031 15895
rect 4614 15892 4642 15932
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 6549 15923 6607 15929
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 9640 15932 10149 15960
rect 9640 15920 9646 15932
rect 10137 15929 10149 15932
rect 10183 15929 10195 15963
rect 10137 15923 10195 15929
rect 13170 15920 13176 15972
rect 13228 15960 13234 15972
rect 13326 15963 13384 15969
rect 13326 15960 13338 15963
rect 13228 15932 13338 15960
rect 13228 15920 13234 15932
rect 13326 15929 13338 15932
rect 13372 15929 13384 15963
rect 13326 15923 13384 15929
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15929 16359 15963
rect 16482 15960 16488 15972
rect 16443 15932 16488 15960
rect 16301 15923 16359 15929
rect 5626 15892 5632 15904
rect 4019 15864 4642 15892
rect 5587 15864 5632 15892
rect 4019 15861 4031 15864
rect 3973 15855 4031 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7834 15892 7840 15904
rect 7795 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 10045 15895 10103 15901
rect 10045 15892 10057 15895
rect 9732 15864 10057 15892
rect 9732 15852 9738 15864
rect 10045 15861 10057 15864
rect 10091 15861 10103 15895
rect 14458 15892 14464 15904
rect 14419 15864 14464 15892
rect 10045 15855 10103 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15746 15892 15752 15904
rect 15707 15864 15752 15892
rect 15746 15852 15752 15864
rect 15804 15892 15810 15904
rect 16316 15892 16344 15923
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 15804 15864 16344 15892
rect 15804 15852 15810 15864
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 3326 15688 3332 15700
rect 3283 15660 3332 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 3326 15648 3332 15660
rect 3384 15688 3390 15700
rect 5258 15688 5264 15700
rect 3384 15660 5264 15688
rect 3384 15648 3390 15660
rect 5258 15648 5264 15660
rect 5316 15688 5322 15700
rect 5537 15691 5595 15697
rect 5537 15688 5549 15691
rect 5316 15660 5549 15688
rect 5316 15648 5322 15660
rect 5537 15657 5549 15660
rect 5583 15688 5595 15691
rect 5626 15688 5632 15700
rect 5583 15660 5632 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 10100 15660 11253 15688
rect 10100 15648 10106 15660
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 11241 15651 11299 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 12492 15660 12633 15688
rect 12492 15648 12498 15660
rect 12621 15657 12633 15660
rect 12667 15657 12679 15691
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 12621 15651 12679 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 16025 15691 16083 15697
rect 16025 15657 16037 15691
rect 16071 15688 16083 15691
rect 16482 15688 16488 15700
rect 16071 15660 16488 15688
rect 16071 15657 16083 15660
rect 16025 15651 16083 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 2498 15580 2504 15632
rect 2556 15620 2562 15632
rect 2685 15623 2743 15629
rect 2685 15620 2697 15623
rect 2556 15592 2697 15620
rect 2556 15580 2562 15592
rect 2685 15589 2697 15592
rect 2731 15589 2743 15623
rect 2685 15583 2743 15589
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 5350 15620 5356 15632
rect 4663 15592 5356 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 5350 15580 5356 15592
rect 5408 15580 5414 15632
rect 5896 15623 5954 15629
rect 5896 15589 5908 15623
rect 5942 15620 5954 15623
rect 5994 15620 6000 15632
rect 5942 15592 6000 15620
rect 5942 15589 5954 15592
rect 5896 15583 5954 15589
rect 5994 15580 6000 15592
rect 6052 15620 6058 15632
rect 6362 15620 6368 15632
rect 6052 15592 6368 15620
rect 6052 15580 6058 15592
rect 6362 15580 6368 15592
rect 6420 15580 6426 15632
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 10134 15620 10140 15632
rect 9548 15592 10140 15620
rect 9548 15580 9554 15592
rect 10134 15580 10140 15592
rect 10192 15620 10198 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 10192 15592 10241 15620
rect 10192 15580 10198 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10778 15620 10784 15632
rect 10739 15592 10784 15620
rect 10229 15583 10287 15589
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15552 1731 15555
rect 1719 15524 2820 15552
rect 1719 15521 1731 15524
rect 1673 15515 1731 15521
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2682 15484 2688 15496
rect 2087 15456 2688 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 2792 15493 2820 15524
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 4890 15552 4896 15564
rect 4212 15524 4896 15552
rect 4212 15512 4218 15524
rect 4890 15512 4896 15524
rect 4948 15552 4954 15564
rect 5169 15555 5227 15561
rect 5169 15552 5181 15555
rect 4948 15524 5181 15552
rect 4948 15512 4954 15524
rect 5169 15521 5181 15524
rect 5215 15552 5227 15555
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5215 15524 5641 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 5629 15521 5641 15524
rect 5675 15552 5687 15555
rect 6454 15552 6460 15564
rect 5675 15524 6460 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 9122 15552 9128 15564
rect 9035 15524 9128 15552
rect 9122 15512 9128 15524
rect 9180 15552 9186 15564
rect 10318 15552 10324 15564
rect 9180 15524 10324 15552
rect 9180 15512 9186 15524
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 2866 15484 2872 15496
rect 2823 15456 2872 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4764 15456 4809 15484
rect 4764 15444 4770 15456
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9916 15456 10149 15484
rect 9916 15444 9922 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 7006 15416 7012 15428
rect 6967 15388 7012 15416
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 9732 15388 9781 15416
rect 9732 15376 9738 15388
rect 9769 15385 9781 15388
rect 9815 15385 9827 15419
rect 9769 15379 9827 15385
rect 2222 15348 2228 15360
rect 2183 15320 2228 15348
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2498 15308 2504 15360
rect 2556 15348 2562 15360
rect 2682 15348 2688 15360
rect 2556 15320 2688 15348
rect 2556 15308 2562 15320
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 3878 15348 3884 15360
rect 3839 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 5166 15348 5172 15360
rect 4203 15320 5172 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9582 15348 9588 15360
rect 9539 15320 9588 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15144 4215 15147
rect 4706 15144 4712 15156
rect 4203 15116 4712 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5258 15144 5264 15156
rect 5219 15116 5264 15144
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 5408 15116 6561 15144
rect 5408 15104 5414 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 6549 15107 6607 15113
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 4724 15076 4752 15104
rect 6730 15076 6736 15088
rect 4724 15048 6736 15076
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 9766 15076 9772 15088
rect 9723 15048 9772 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 1394 14968 1400 15020
rect 1452 15008 1458 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1452 14980 1685 15008
rect 1452 14968 1458 14980
rect 1673 14977 1685 14980
rect 1719 15008 1731 15011
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1719 14980 2053 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2041 14977 2053 14980
rect 2087 15008 2099 15011
rect 2130 15008 2136 15020
rect 2087 14980 2136 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 4755 14980 5825 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5813 14977 5825 14980
rect 5859 15008 5871 15011
rect 5994 15008 6000 15020
rect 5859 14980 6000 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 2400 14943 2458 14949
rect 2400 14909 2412 14943
rect 2446 14940 2458 14943
rect 2866 14940 2872 14952
rect 2446 14912 2872 14940
rect 2446 14909 2458 14912
rect 2400 14903 2458 14909
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 7285 14943 7343 14949
rect 5123 14912 5764 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5258 14832 5264 14884
rect 5316 14872 5322 14884
rect 5736 14881 5764 14912
rect 7285 14909 7297 14943
rect 7331 14909 7343 14943
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 7285 14903 7343 14909
rect 9232 14912 9781 14940
rect 5537 14875 5595 14881
rect 5537 14872 5549 14875
rect 5316 14844 5549 14872
rect 5316 14832 5322 14844
rect 5537 14841 5549 14844
rect 5583 14841 5595 14875
rect 5537 14835 5595 14841
rect 5721 14875 5779 14881
rect 5721 14841 5733 14875
rect 5767 14872 5779 14875
rect 6086 14872 6092 14884
rect 5767 14844 6092 14872
rect 5767 14841 5779 14844
rect 5721 14835 5779 14841
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 6273 14807 6331 14813
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6454 14804 6460 14816
rect 6319 14776 6460 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6454 14764 6460 14776
rect 6512 14804 6518 14816
rect 7101 14807 7159 14813
rect 7101 14804 7113 14807
rect 6512 14776 7113 14804
rect 6512 14764 6518 14776
rect 7101 14773 7113 14776
rect 7147 14804 7159 14807
rect 7300 14804 7328 14903
rect 7374 14832 7380 14884
rect 7432 14872 7438 14884
rect 7530 14875 7588 14881
rect 7530 14872 7542 14875
rect 7432 14844 7542 14872
rect 7432 14832 7438 14844
rect 7530 14841 7542 14844
rect 7576 14841 7588 14875
rect 7530 14835 7588 14841
rect 9232 14813 9260 14912
rect 9769 14909 9781 14912
rect 9815 14940 9827 14943
rect 9858 14940 9864 14952
rect 9815 14912 9864 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10036 14943 10094 14949
rect 10036 14909 10048 14943
rect 10082 14940 10094 14943
rect 10318 14940 10324 14952
rect 10082 14912 10324 14940
rect 10082 14909 10094 14912
rect 10036 14903 10094 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 7147 14776 9229 14804
rect 7147 14773 7159 14776
rect 7101 14767 7159 14773
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 9732 14776 11161 14804
rect 9732 14764 9738 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2648 14572 2789 14600
rect 2648 14560 2654 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 3329 14603 3387 14609
rect 3329 14600 3341 14603
rect 2924 14572 3341 14600
rect 2924 14560 2930 14572
rect 3329 14569 3341 14572
rect 3375 14569 3387 14603
rect 3329 14563 3387 14569
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 3697 14603 3755 14609
rect 3697 14600 3709 14603
rect 3568 14572 3709 14600
rect 3568 14560 3574 14572
rect 3697 14569 3709 14572
rect 3743 14569 3755 14603
rect 3697 14563 3755 14569
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4304 14572 4629 14600
rect 4304 14560 4310 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 5721 14603 5779 14609
rect 5721 14569 5733 14603
rect 5767 14600 5779 14603
rect 5994 14600 6000 14612
rect 5767 14572 6000 14600
rect 5767 14569 5779 14572
rect 5721 14563 5779 14569
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 9122 14600 9128 14612
rect 7055 14572 8156 14600
rect 9083 14572 9128 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 3878 14492 3884 14544
rect 3936 14532 3942 14544
rect 4430 14532 4436 14544
rect 3936 14504 4436 14532
rect 3936 14492 3942 14504
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 6457 14535 6515 14541
rect 6457 14501 6469 14535
rect 6503 14532 6515 14535
rect 6503 14504 7604 14532
rect 6503 14501 6515 14504
rect 6457 14495 6515 14501
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1670 14473 1676 14476
rect 1664 14464 1676 14473
rect 1631 14436 1676 14464
rect 1664 14427 1676 14436
rect 1670 14424 1676 14427
rect 1728 14424 1734 14476
rect 5258 14464 5264 14476
rect 5219 14436 5264 14464
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5994 14424 6000 14476
rect 6052 14464 6058 14476
rect 6273 14467 6331 14473
rect 6273 14464 6285 14467
rect 6052 14436 6285 14464
rect 6052 14424 6058 14436
rect 6273 14433 6285 14436
rect 6319 14433 6331 14467
rect 6273 14427 6331 14433
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4396 14368 4721 14396
rect 4396 14356 4402 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14396 6607 14399
rect 7374 14396 7380 14408
rect 6595 14368 7380 14396
rect 6595 14365 6607 14368
rect 6549 14359 6607 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 4157 14331 4215 14337
rect 4157 14297 4169 14331
rect 4203 14328 4215 14331
rect 5350 14328 5356 14340
rect 4203 14300 5356 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 7576 14337 7604 14504
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 7708 14504 7849 14532
rect 7708 14492 7714 14504
rect 7837 14501 7849 14504
rect 7883 14501 7895 14535
rect 7837 14495 7895 14501
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 8021 14535 8079 14541
rect 8021 14532 8033 14535
rect 7984 14504 8033 14532
rect 7984 14492 7990 14504
rect 8021 14501 8033 14504
rect 8067 14501 8079 14535
rect 8021 14495 8079 14501
rect 8128 14405 8156 14572
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9490 14600 9496 14612
rect 9451 14572 9496 14600
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 14090 14492 14096 14544
rect 14148 14532 14154 14544
rect 14274 14532 14280 14544
rect 14148 14504 14280 14532
rect 14148 14492 14154 14504
rect 14274 14492 14280 14504
rect 14332 14492 14338 14544
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 10209 14467 10267 14473
rect 10209 14464 10221 14467
rect 9732 14436 10221 14464
rect 9732 14424 9738 14436
rect 10209 14433 10221 14436
rect 10255 14433 10267 14467
rect 10209 14427 10267 14433
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9916 14368 9965 14396
rect 9916 14356 9922 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 7561 14331 7619 14337
rect 7561 14297 7573 14331
rect 7607 14328 7619 14331
rect 8481 14331 8539 14337
rect 8481 14328 8493 14331
rect 7607 14300 8493 14328
rect 7607 14297 7619 14300
rect 7561 14291 7619 14297
rect 8481 14297 8493 14300
rect 8527 14297 8539 14331
rect 8481 14291 8539 14297
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 3476 14232 6009 14260
rect 3476 14220 3482 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 5997 14223 6055 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 11330 14260 11336 14272
rect 11291 14232 11336 14260
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 4488 14028 4629 14056
rect 4488 14016 4494 14028
rect 4617 14025 4629 14028
rect 4663 14025 4675 14059
rect 4617 14019 4675 14025
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6086 14056 6092 14068
rect 5675 14028 6092 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 1486 13988 1492 14000
rect 1447 13960 1492 13988
rect 1486 13948 1492 13960
rect 1544 13948 1550 14000
rect 3050 13988 3056 14000
rect 3011 13960 3056 13988
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3973 13991 4031 13997
rect 3973 13988 3985 13991
rect 3200 13960 3985 13988
rect 3200 13948 3206 13960
rect 3973 13957 3985 13960
rect 4019 13957 4031 13991
rect 3973 13951 4031 13957
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2590 13920 2596 13932
rect 2087 13892 2596 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3568 13892 3617 13920
rect 3568 13880 3574 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 3988 13852 4016 13951
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4948 13892 5181 13920
rect 4948 13880 4954 13892
rect 5169 13889 5181 13892
rect 5215 13920 5227 13923
rect 5644 13920 5672 14019
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14056 6423 14059
rect 7374 14056 7380 14068
rect 6411 14028 7380 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 7374 14016 7380 14028
rect 7432 14056 7438 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 7432 14028 9045 14056
rect 7432 14016 7438 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 9033 14019 9091 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 7193 13991 7251 13997
rect 7193 13957 7205 13991
rect 7239 13988 7251 13991
rect 7282 13988 7288 14000
rect 7239 13960 7288 13988
rect 7239 13957 7251 13960
rect 7193 13951 7251 13957
rect 7282 13948 7288 13960
rect 7340 13988 7346 14000
rect 7650 13988 7656 14000
rect 7340 13960 7656 13988
rect 7340 13948 7346 13960
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 9858 13948 9864 14000
rect 9916 13988 9922 14000
rect 10321 13991 10379 13997
rect 10321 13988 10333 13991
rect 9916 13960 10333 13988
rect 9916 13948 9922 13960
rect 10321 13957 10333 13960
rect 10367 13957 10379 13991
rect 10321 13951 10379 13957
rect 7558 13920 7564 13932
rect 5215 13892 5672 13920
rect 7519 13892 7564 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 4430 13852 4436 13864
rect 2547 13824 3372 13852
rect 3988 13824 4436 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 3344 13796 3372 13824
rect 4430 13812 4436 13824
rect 4488 13852 4494 13864
rect 5994 13852 6000 13864
rect 4488 13824 4936 13852
rect 5955 13824 6000 13852
rect 4488 13812 4494 13824
rect 1762 13784 1768 13796
rect 1723 13756 1768 13784
rect 1762 13744 1768 13756
rect 1820 13744 1826 13796
rect 3050 13784 3056 13796
rect 2792 13756 3056 13784
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2792 13716 2820 13756
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3326 13784 3332 13796
rect 3287 13756 3332 13784
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 3513 13787 3571 13793
rect 3513 13753 3525 13787
rect 3559 13784 3571 13787
rect 3602 13784 3608 13796
rect 3559 13756 3608 13784
rect 3559 13753 3571 13756
rect 3513 13747 3571 13753
rect 1995 13688 2820 13716
rect 2869 13719 2927 13725
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2869 13685 2881 13719
rect 2915 13716 2927 13719
rect 3528 13716 3556 13747
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 4908 13793 4936 13824
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6454 13812 6460 13864
rect 6512 13852 6518 13864
rect 7653 13855 7711 13861
rect 7653 13852 7665 13855
rect 6512 13824 7665 13852
rect 6512 13812 6518 13824
rect 7653 13821 7665 13824
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 7920 13855 7978 13861
rect 7920 13821 7932 13855
rect 7966 13852 7978 13855
rect 8202 13852 8208 13864
rect 7966 13824 8208 13852
rect 7966 13821 7978 13824
rect 7920 13815 7978 13821
rect 4893 13787 4951 13793
rect 4893 13753 4905 13787
rect 4939 13753 4951 13787
rect 7668 13784 7696 13815
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 10134 13852 10140 13864
rect 10095 13824 10140 13852
rect 10134 13812 10140 13824
rect 10192 13852 10198 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10192 13824 10701 13852
rect 10192 13812 10198 13824
rect 10689 13821 10701 13824
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 8110 13784 8116 13796
rect 7668 13756 8116 13784
rect 4893 13747 4951 13753
rect 8110 13744 8116 13756
rect 8168 13744 8174 13796
rect 2915 13688 3556 13716
rect 4433 13719 4491 13725
rect 2915 13685 2927 13688
rect 2869 13679 2927 13685
rect 4433 13685 4445 13719
rect 4479 13716 4491 13719
rect 5074 13716 5080 13728
rect 4479 13688 5080 13716
rect 4479 13685 4491 13688
rect 4433 13679 4491 13685
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 3234 13512 3240 13524
rect 2547 13484 3240 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4338 13512 4344 13524
rect 3927 13484 4344 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4338 13472 4344 13484
rect 4396 13512 4402 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 4396 13484 6009 13512
rect 4396 13472 4402 13484
rect 5997 13481 6009 13484
rect 6043 13512 6055 13515
rect 6178 13512 6184 13524
rect 6043 13484 6184 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 6788 13484 6837 13512
rect 6788 13472 6794 13484
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8260 13484 8585 13512
rect 8260 13472 8266 13484
rect 8573 13481 8585 13484
rect 8619 13512 8631 13515
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 8619 13484 11069 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 1949 13447 2007 13453
rect 1949 13413 1961 13447
rect 1995 13444 2007 13447
rect 2130 13444 2136 13456
rect 1995 13416 2136 13444
rect 1995 13413 2007 13416
rect 1949 13407 2007 13413
rect 2130 13404 2136 13416
rect 2188 13404 2194 13456
rect 4890 13453 4896 13456
rect 4249 13447 4307 13453
rect 4249 13413 4261 13447
rect 4295 13444 4307 13447
rect 4884 13444 4896 13453
rect 4295 13416 4896 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 4884 13407 4896 13416
rect 4890 13404 4896 13407
rect 4948 13404 4954 13456
rect 7650 13444 7656 13456
rect 7611 13416 7656 13444
rect 7650 13404 7656 13416
rect 7708 13444 7714 13456
rect 8849 13447 8907 13453
rect 8849 13444 8861 13447
rect 7708 13416 8861 13444
rect 7708 13404 7714 13416
rect 8849 13413 8861 13416
rect 8895 13413 8907 13447
rect 8849 13407 8907 13413
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 1854 13376 1860 13388
rect 1811 13348 1860 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 1854 13336 1860 13348
rect 1912 13376 1918 13388
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 1912 13348 2973 13376
rect 1912 13336 1918 13348
rect 2961 13345 2973 13348
rect 3007 13345 3019 13379
rect 2961 13339 3019 13345
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7834 13376 7840 13388
rect 7515 13348 7840 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 9944 13379 10002 13385
rect 9944 13376 9956 13379
rect 9824 13348 9956 13376
rect 9824 13336 9830 13348
rect 9944 13345 9956 13348
rect 9990 13376 10002 13379
rect 10502 13376 10508 13388
rect 9990 13348 10508 13376
rect 9990 13345 10002 13348
rect 9944 13339 10002 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1728 13280 2053 13308
rect 1728 13268 1734 13280
rect 2041 13277 2053 13280
rect 2087 13308 2099 13311
rect 3510 13308 3516 13320
rect 2087 13280 3516 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13240 1547 13243
rect 1762 13240 1768 13252
rect 1535 13212 1768 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 1762 13200 1768 13212
rect 1820 13240 1826 13252
rect 2498 13240 2504 13252
rect 1820 13212 2504 13240
rect 1820 13200 1826 13212
rect 2498 13200 2504 13212
rect 2556 13200 2562 13252
rect 2866 13172 2872 13184
rect 2827 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 4632 13172 4660 13271
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 6236 13280 7757 13308
rect 6236 13268 6242 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 7190 13240 7196 13252
rect 7151 13212 7196 13240
rect 7190 13200 7196 13212
rect 7248 13200 7254 13252
rect 4982 13172 4988 13184
rect 4632 13144 4988 13172
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 8110 13172 8116 13184
rect 8071 13144 8116 13172
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 9692 13172 9720 13271
rect 10042 13172 10048 13184
rect 9692 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4062 12968 4068 12980
rect 4019 12940 4068 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4948 12940 5273 12968
rect 4948 12928 4954 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 5261 12931 5319 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12968 10655 12971
rect 10962 12968 10968 12980
rect 10643 12940 10968 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 9674 12900 9680 12912
rect 9635 12872 9680 12900
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 11333 12903 11391 12909
rect 11333 12900 11345 12903
rect 10744 12872 11345 12900
rect 10744 12860 10750 12872
rect 11333 12869 11345 12872
rect 11379 12869 11391 12903
rect 11333 12863 11391 12869
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3384 12804 3433 12832
rect 3384 12792 3390 12804
rect 3421 12801 3433 12804
rect 3467 12832 3479 12835
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 3467 12804 4445 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 4433 12801 4445 12804
rect 4479 12832 4491 12835
rect 4614 12832 4620 12844
rect 4479 12804 4620 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2924 12736 2973 12764
rect 2924 12724 2930 12736
rect 2961 12733 2973 12736
rect 3007 12764 3019 12767
rect 4890 12764 4896 12776
rect 3007 12736 4896 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 4540 12705 4568 12736
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12764 5506 12776
rect 5994 12764 6000 12776
rect 5500 12736 6000 12764
rect 5500 12724 5506 12736
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6564 12736 6837 12764
rect 2685 12699 2743 12705
rect 2685 12665 2697 12699
rect 2731 12665 2743 12699
rect 2685 12659 2743 12665
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12665 4583 12699
rect 4525 12659 4583 12665
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 6454 12696 6460 12708
rect 5767 12668 6460 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12628 1731 12631
rect 2130 12628 2136 12640
rect 1719 12600 2136 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 2130 12588 2136 12600
rect 2188 12628 2194 12640
rect 2700 12628 2728 12659
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 6564 12640 6592 12736
rect 6825 12733 6837 12736
rect 6871 12764 6883 12767
rect 8110 12764 8116 12776
rect 6871 12736 8116 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 11072 12764 11100 12792
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 11072 12736 11161 12764
rect 11149 12733 11161 12736
rect 11195 12764 11207 12767
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 11195 12736 11713 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11701 12733 11713 12736
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7070 12699 7128 12705
rect 7070 12696 7082 12699
rect 6788 12668 7082 12696
rect 6788 12656 6794 12668
rect 7070 12665 7082 12668
rect 7116 12665 7128 12699
rect 9953 12699 10011 12705
rect 9953 12696 9965 12699
rect 7070 12659 7128 12665
rect 9048 12668 9965 12696
rect 9048 12640 9076 12668
rect 9953 12665 9965 12668
rect 9999 12665 10011 12699
rect 9953 12659 10011 12665
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10275 12668 10977 12696
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 10965 12665 10977 12668
rect 11011 12696 11023 12699
rect 11054 12696 11060 12708
rect 11011 12668 11060 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 2866 12628 2872 12640
rect 2188 12600 2728 12628
rect 2779 12600 2872 12628
rect 2188 12588 2194 12600
rect 2866 12588 2872 12600
rect 2924 12628 2930 12640
rect 3234 12628 3240 12640
rect 2924 12600 3240 12628
rect 2924 12588 2930 12600
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3789 12631 3847 12637
rect 3789 12597 3801 12631
rect 3835 12628 3847 12631
rect 4433 12631 4491 12637
rect 4433 12628 4445 12631
rect 3835 12600 4445 12628
rect 3835 12597 3847 12600
rect 3789 12591 3847 12597
rect 4433 12597 4445 12600
rect 4479 12628 4491 12631
rect 4798 12628 4804 12640
rect 4479 12600 4804 12628
rect 4479 12597 4491 12600
rect 4433 12591 4491 12597
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 9539 12600 10149 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 10137 12597 10149 12600
rect 10183 12628 10195 12631
rect 11146 12628 11152 12640
rect 10183 12600 11152 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 2590 12424 2596 12436
rect 2363 12396 2596 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 2832 12396 3433 12424
rect 2832 12384 2838 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3421 12387 3479 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4062 12424 4068 12436
rect 3927 12396 4068 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4706 12424 4712 12436
rect 4667 12396 4712 12424
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 6641 12427 6699 12433
rect 6641 12393 6653 12427
rect 6687 12424 6699 12427
rect 6730 12424 6736 12436
rect 6687 12396 6736 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7834 12424 7840 12436
rect 7331 12396 7840 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8846 12424 8852 12436
rect 8619 12396 8852 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8846 12384 8852 12396
rect 8904 12424 8910 12436
rect 9582 12424 9588 12436
rect 8904 12396 9588 12424
rect 8904 12384 8910 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 11020 12396 11437 12424
rect 11020 12384 11026 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 4154 12356 4160 12368
rect 3007 12328 4160 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 5528 12359 5586 12365
rect 5528 12325 5540 12359
rect 5574 12356 5586 12359
rect 6178 12356 6184 12368
rect 5574 12328 6184 12356
rect 5574 12325 5586 12328
rect 5528 12319 5586 12325
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 5040 12260 5273 12288
rect 5040 12248 5046 12260
rect 5261 12257 5273 12260
rect 5307 12288 5319 12291
rect 6546 12288 6552 12300
rect 5307 12260 6552 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8628 12260 8677 12288
rect 8628 12248 8634 12260
rect 8665 12257 8677 12260
rect 8711 12288 8723 12291
rect 9582 12288 9588 12300
rect 8711 12260 9588 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 10301 12291 10359 12297
rect 10301 12288 10313 12291
rect 9784 12260 10313 12288
rect 9784 12232 9812 12260
rect 10301 12257 10313 12260
rect 10347 12288 10359 12291
rect 11054 12288 11060 12300
rect 10347 12260 11060 12288
rect 10347 12257 10359 12260
rect 10301 12251 10359 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 2038 12220 2044 12232
rect 1443 12192 2044 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2958 12220 2964 12232
rect 2919 12192 2964 12220
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3602 12220 3608 12232
rect 3099 12192 3608 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 8202 12152 8208 12164
rect 7852 12124 8208 12152
rect 7852 12096 7880 12124
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 10060 12096 10088 12183
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 2682 12084 2688 12096
rect 2547 12056 2688 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4028 12056 4261 12084
rect 4028 12044 4034 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5258 12084 5264 12096
rect 5215 12056 5264 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 7834 12084 7840 12096
rect 7795 12056 7840 12084
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 9953 12087 10011 12093
rect 9953 12053 9965 12087
rect 9999 12084 10011 12087
rect 10042 12084 10048 12096
rect 9999 12056 10048 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 4798 11880 4804 11892
rect 3016 11852 4804 11880
rect 3016 11840 3022 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7285 11883 7343 11889
rect 7285 11849 7297 11883
rect 7331 11880 7343 11883
rect 8478 11880 8484 11892
rect 7331 11852 8484 11880
rect 7331 11849 7343 11852
rect 7285 11843 7343 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 4157 11815 4215 11821
rect 4157 11812 4169 11815
rect 4120 11784 4169 11812
rect 4120 11772 4126 11784
rect 4157 11781 4169 11784
rect 4203 11781 4215 11815
rect 4157 11775 4215 11781
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 6052 11784 6469 11812
rect 6052 11772 6058 11784
rect 6457 11781 6469 11784
rect 6503 11781 6515 11815
rect 6457 11775 6515 11781
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 2179 11648 2237 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2225 11645 2237 11648
rect 2271 11676 2283 11679
rect 3234 11676 3240 11688
rect 2271 11648 3240 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 4764 11648 5089 11676
rect 4764 11636 4770 11648
rect 5077 11645 5089 11648
rect 5123 11645 5135 11679
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 5077 11639 5135 11645
rect 7576 11648 7757 11676
rect 2492 11611 2550 11617
rect 2492 11577 2504 11611
rect 2538 11608 2550 11611
rect 2590 11608 2596 11620
rect 2538 11580 2596 11608
rect 2538 11577 2550 11580
rect 2492 11571 2550 11577
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 5350 11608 5356 11620
rect 5311 11580 5356 11608
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 5074 11540 5080 11552
rect 4663 11512 5080 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5074 11500 5080 11512
rect 5132 11540 5138 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 5132 11512 5273 11540
rect 5132 11500 5138 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 6546 11540 6552 11552
rect 5859 11512 6552 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 6546 11500 6552 11512
rect 6604 11540 6610 11552
rect 7006 11540 7012 11552
rect 6604 11512 7012 11540
rect 6604 11500 6610 11512
rect 7006 11500 7012 11512
rect 7064 11540 7070 11552
rect 7576 11549 7604 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 10226 11676 10232 11688
rect 10187 11648 10232 11676
rect 7745 11639 7803 11645
rect 10226 11636 10232 11648
rect 10284 11676 10290 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10284 11648 10793 11676
rect 10284 11636 10290 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 7990 11611 8048 11617
rect 7990 11608 8002 11611
rect 7760 11580 8002 11608
rect 7760 11552 7788 11580
rect 7990 11577 8002 11580
rect 8036 11577 8048 11611
rect 7990 11571 8048 11577
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 7064 11512 7573 11540
rect 7064 11500 7070 11512
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7561 11503 7619 11509
rect 7742 11500 7748 11552
rect 7800 11500 7806 11552
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 9582 11540 9588 11552
rect 9171 11512 9588 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 10192 11512 10425 11540
rect 10192 11500 10198 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2501 11339 2559 11345
rect 2501 11336 2513 11339
rect 1728 11308 2513 11336
rect 1728 11296 1734 11308
rect 2501 11305 2513 11308
rect 2547 11336 2559 11339
rect 2866 11336 2872 11348
rect 2547 11308 2872 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3697 11339 3755 11345
rect 3697 11336 3709 11339
rect 3108 11308 3709 11336
rect 3108 11296 3114 11308
rect 3697 11305 3709 11308
rect 3743 11305 3755 11339
rect 3697 11299 3755 11305
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 4856 11308 6561 11336
rect 4856 11296 4862 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7926 11336 7932 11348
rect 6972 11308 7932 11336
rect 6972 11296 6978 11308
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8570 11336 8576 11348
rect 8527 11308 8576 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 11609 11339 11667 11345
rect 11609 11336 11621 11339
rect 9824 11308 11621 11336
rect 9824 11296 9830 11308
rect 11609 11305 11621 11308
rect 11655 11305 11667 11339
rect 11609 11299 11667 11305
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 4617 11271 4675 11277
rect 1811 11240 2636 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 2608 11212 2636 11240
rect 4617 11237 4629 11271
rect 4663 11268 4675 11271
rect 4706 11268 4712 11280
rect 4663 11240 4712 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 12912 11268 12940 11299
rect 9732 11240 12940 11268
rect 9732 11228 9738 11240
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 2130 11200 2136 11212
rect 1912 11172 2136 11200
rect 1912 11160 1918 11172
rect 2130 11160 2136 11172
rect 2188 11200 2194 11212
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 2188 11172 2329 11200
rect 2188 11160 2194 11172
rect 2317 11169 2329 11172
rect 2363 11169 2375 11203
rect 2590 11200 2596 11212
rect 2503 11172 2596 11200
rect 2317 11163 2375 11169
rect 2590 11160 2596 11172
rect 2648 11200 2654 11212
rect 3053 11203 3111 11209
rect 3053 11200 3065 11203
rect 2648 11172 3065 11200
rect 2648 11160 2654 11172
rect 3053 11169 3065 11172
rect 3099 11200 3111 11203
rect 3099 11172 4752 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4724 11141 4752 11172
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5500 11172 5641 11200
rect 5500 11160 5506 11172
rect 5629 11169 5641 11172
rect 5675 11200 5687 11203
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5675 11172 6193 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 6181 11169 6193 11172
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7800 11172 8033 11200
rect 7800 11160 7806 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 10496 11203 10554 11209
rect 10496 11169 10508 11203
rect 10542 11200 10554 11203
rect 11054 11200 11060 11212
rect 10542 11172 11060 11200
rect 10542 11169 10554 11172
rect 10496 11163 10554 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12710 11200 12716 11212
rect 12671 11172 12716 11200
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4798 11132 4804 11144
rect 4755 11104 4804 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 4798 11092 4804 11104
rect 4856 11132 4862 11144
rect 5350 11132 5356 11144
rect 4856 11104 5356 11132
rect 4856 11092 4862 11104
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 6696 11104 7941 11132
rect 6696 11092 6702 11104
rect 7929 11101 7941 11104
rect 7975 11132 7987 11135
rect 8294 11132 8300 11144
rect 7975 11104 8300 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10226 11132 10232 11144
rect 10100 11104 10232 11132
rect 10100 11092 10106 11104
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 2222 11064 2228 11076
rect 2087 11036 2228 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 2222 11024 2228 11036
rect 2280 11024 2286 11076
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 2832 11036 3341 11064
rect 2832 11024 2838 11036
rect 3329 11033 3341 11036
rect 3375 11064 3387 11067
rect 3602 11064 3608 11076
rect 3375 11036 3608 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 4154 11064 4160 11076
rect 4115 11036 4160 11064
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5442 11064 5448 11076
rect 5307 11036 5448 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5810 11064 5816 11076
rect 5771 11036 5816 11064
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7006 10996 7012 11008
rect 6967 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7466 10996 7472 11008
rect 7427 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 4706 10792 4712 10804
rect 4203 10764 4712 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6822 10792 6828 10804
rect 6687 10764 6828 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 7800 10764 8953 10792
rect 7800 10752 7806 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11606 10792 11612 10804
rect 11112 10764 11612 10792
rect 11112 10752 11118 10764
rect 11606 10752 11612 10764
rect 11664 10792 11670 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11664 10764 11805 10792
rect 11664 10752 11670 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12768 10764 12909 10792
rect 12768 10752 12774 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 5258 10724 5264 10736
rect 5219 10696 5264 10724
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 8386 10724 8392 10736
rect 8347 10696 8392 10724
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5718 10656 5724 10668
rect 5500 10628 5724 10656
rect 5500 10616 5506 10628
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 2406 10597 2412 10600
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10557 2191 10591
rect 2400 10588 2412 10597
rect 2319 10560 2412 10588
rect 2133 10551 2191 10557
rect 2400 10551 2412 10560
rect 2464 10588 2470 10600
rect 2774 10588 2780 10600
rect 2464 10560 2780 10588
rect 2148 10520 2176 10551
rect 2406 10548 2412 10551
rect 2464 10548 2470 10560
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 6362 10588 6368 10600
rect 5736 10560 6368 10588
rect 3234 10520 3240 10532
rect 2148 10492 3240 10520
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 5077 10523 5135 10529
rect 5077 10489 5089 10523
rect 5123 10520 5135 10523
rect 5442 10520 5448 10532
rect 5123 10492 5448 10520
rect 5123 10489 5135 10492
rect 5077 10483 5135 10489
rect 5442 10480 5448 10492
rect 5500 10520 5506 10532
rect 5736 10529 5764 10560
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7006 10588 7012 10600
rect 6919 10560 7012 10588
rect 7006 10548 7012 10560
rect 7064 10588 7070 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 7064 10560 9413 10588
rect 7064 10548 7070 10560
rect 9401 10557 9413 10560
rect 9447 10588 9459 10591
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9447 10560 9505 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9493 10557 9505 10560
rect 9539 10588 9551 10591
rect 9539 10560 9904 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 9876 10532 9904 10560
rect 5721 10523 5779 10529
rect 5721 10520 5733 10523
rect 5500 10492 5733 10520
rect 5500 10480 5506 10492
rect 5721 10489 5733 10492
rect 5767 10489 5779 10523
rect 5721 10483 5779 10489
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 5994 10520 6000 10532
rect 5859 10492 6000 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 7276 10523 7334 10529
rect 7276 10520 7288 10523
rect 6319 10492 7288 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 7276 10489 7288 10492
rect 7322 10520 7334 10523
rect 7926 10520 7932 10532
rect 7322 10492 7932 10520
rect 7322 10489 7334 10492
rect 7276 10483 7334 10489
rect 7926 10480 7932 10492
rect 7984 10520 7990 10532
rect 7984 10492 9444 10520
rect 7984 10480 7990 10492
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1912 10424 1961 10452
rect 1912 10412 1918 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 1949 10415 2007 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 4614 10452 4620 10464
rect 4571 10424 4620 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 9416 10452 9444 10492
rect 9674 10480 9680 10532
rect 9732 10529 9738 10532
rect 9732 10523 9796 10529
rect 9732 10489 9750 10523
rect 9784 10489 9796 10523
rect 9732 10483 9796 10489
rect 9732 10480 9738 10483
rect 9858 10480 9864 10532
rect 9916 10520 9922 10532
rect 10226 10520 10232 10532
rect 9916 10492 10232 10520
rect 9916 10480 9922 10492
rect 10226 10480 10232 10492
rect 10284 10520 10290 10532
rect 11425 10523 11483 10529
rect 11425 10520 11437 10523
rect 10284 10492 11437 10520
rect 10284 10480 10290 10492
rect 11425 10489 11437 10492
rect 11471 10489 11483 10523
rect 11425 10483 11483 10489
rect 12434 10480 12440 10532
rect 12492 10520 12498 10532
rect 12492 10492 12537 10520
rect 12492 10480 12498 10492
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 9416 10424 10885 10452
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 2406 10248 2412 10260
rect 1719 10220 2412 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 2556 10220 3157 10248
rect 2556 10208 2562 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4062 10248 4068 10260
rect 3651 10220 4068 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4798 10248 4804 10260
rect 4387 10220 4804 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7466 10248 7472 10260
rect 7055 10220 7472 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 9861 10211 9919 10217
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 2682 10180 2688 10192
rect 2363 10152 2688 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 3234 10180 3240 10192
rect 2915 10152 3240 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 3234 10140 3240 10152
rect 3292 10180 3298 10192
rect 4982 10180 4988 10192
rect 3292 10152 4988 10180
rect 3292 10140 3298 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 7653 10183 7711 10189
rect 7653 10149 7665 10183
rect 7699 10180 7711 10183
rect 8202 10180 8208 10192
rect 7699 10152 8208 10180
rect 7699 10149 7711 10152
rect 7653 10143 7711 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 7340 10084 7481 10112
rect 7340 10072 7346 10084
rect 7469 10081 7481 10084
rect 7515 10112 7527 10115
rect 7558 10112 7564 10124
rect 7515 10084 7564 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 10496 10115 10554 10121
rect 10496 10081 10508 10115
rect 10542 10112 10554 10115
rect 10870 10112 10876 10124
rect 10542 10084 10876 10112
rect 10542 10081 10554 10084
rect 10496 10075 10554 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3510 10044 3516 10056
rect 2455 10016 3516 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4967 10047 5025 10053
rect 4967 10044 4979 10047
rect 4120 10016 4979 10044
rect 4120 10004 4126 10016
rect 4967 10013 4979 10016
rect 5013 10013 5025 10047
rect 5442 10044 5448 10056
rect 5403 10016 5448 10044
rect 4967 10007 5025 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 5537 10007 5595 10013
rect 5552 9976 5580 10007
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 9916 10016 10241 10044
rect 9916 10004 9922 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 4816 9948 5580 9976
rect 4816 9920 4844 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 2130 9908 2136 9920
rect 1903 9880 2136 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 4798 9908 4804 9920
rect 4759 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5994 9908 6000 9920
rect 5955 9880 6000 9908
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 7282 9908 7288 9920
rect 7239 9880 7288 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 8386 9908 8392 9920
rect 8251 9880 8392 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 9122 9908 9128 9920
rect 8619 9880 9128 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 3142 9704 3148 9716
rect 3103 9676 3148 9704
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 5261 9707 5319 9713
rect 5261 9673 5273 9707
rect 5307 9704 5319 9707
rect 5350 9704 5356 9716
rect 5307 9676 5356 9704
rect 5307 9673 5319 9676
rect 5261 9667 5319 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 7742 9704 7748 9716
rect 6840 9676 7748 9704
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 2314 9636 2320 9648
rect 1811 9608 2320 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 2314 9596 2320 9608
rect 2372 9636 2378 9648
rect 2958 9636 2964 9648
rect 2372 9608 2964 9636
rect 2372 9596 2378 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 5534 9636 5540 9648
rect 5495 9608 5540 9636
rect 5534 9596 5540 9608
rect 5592 9636 5598 9648
rect 6273 9639 6331 9645
rect 5592 9608 5764 9636
rect 5592 9596 5598 9608
rect 5736 9577 5764 9608
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 6840 9636 6868 9676
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 14274 9704 14280 9716
rect 14148 9676 14280 9704
rect 14148 9664 14154 9676
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 6319 9608 6868 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 7558 9596 7564 9648
rect 7616 9596 7622 9648
rect 8570 9636 8576 9648
rect 8531 9608 8576 9636
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 10321 9639 10379 9645
rect 10321 9605 10333 9639
rect 10367 9636 10379 9639
rect 11698 9636 11704 9648
rect 10367 9608 11704 9636
rect 10367 9605 10379 9608
rect 10321 9599 10379 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 5721 9571 5779 9577
rect 2823 9540 3372 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2406 9500 2412 9512
rect 2363 9472 2412 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 3200 9472 3249 9500
rect 3200 9460 3206 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3344 9500 3372 9540
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7190 9568 7196 9580
rect 6687 9540 7196 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7190 9528 7196 9540
rect 7248 9568 7254 9580
rect 7576 9568 7604 9596
rect 7248 9540 7604 9568
rect 7248 9528 7254 9540
rect 8386 9528 8392 9580
rect 8444 9568 8450 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8444 9540 8953 9568
rect 8444 9528 8450 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 9122 9568 9128 9580
rect 9083 9540 9128 9568
rect 8941 9531 8999 9537
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 10870 9568 10876 9580
rect 10831 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9568 10934 9580
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 10928 9540 11253 9568
rect 10928 9528 10934 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 3510 9509 3516 9512
rect 3504 9500 3516 9509
rect 3344 9472 3516 9500
rect 3237 9463 3295 9469
rect 3504 9463 3516 9472
rect 3510 9460 3516 9463
rect 3568 9460 3574 9512
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7800 9472 8033 9500
rect 7800 9460 7806 9472
rect 8021 9469 8033 9472
rect 8067 9500 8079 9503
rect 8202 9500 8208 9512
rect 8067 9472 8208 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8202 9460 8208 9472
rect 8260 9500 8266 9512
rect 10137 9503 10195 9509
rect 8260 9472 9812 9500
rect 8260 9460 8266 9472
rect 2222 9432 2228 9444
rect 2183 9404 2228 9432
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 7282 9432 7288 9444
rect 7243 9404 7288 9432
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 7466 9432 7472 9444
rect 7427 9404 7472 9432
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 7561 9435 7619 9441
rect 7561 9401 7573 9435
rect 7607 9432 7619 9435
rect 7834 9432 7840 9444
rect 7607 9404 7840 9432
rect 7607 9401 7619 9404
rect 7561 9395 7619 9401
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 9030 9432 9036 9444
rect 8991 9404 9036 9432
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 9784 9441 9812 9472
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10183 9472 10824 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 9769 9435 9827 9441
rect 9769 9401 9781 9435
rect 9815 9432 9827 9435
rect 10597 9435 10655 9441
rect 10597 9432 10609 9435
rect 9815 9404 10609 9432
rect 9815 9401 9827 9404
rect 9769 9395 9827 9401
rect 10597 9401 10609 9404
rect 10643 9432 10655 9435
rect 10686 9432 10692 9444
rect 10643 9404 10692 9432
rect 10643 9401 10655 9404
rect 10597 9395 10655 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 10796 9441 10824 9472
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 11238 9432 11244 9444
rect 10827 9404 11244 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4890 9364 4896 9376
rect 4663 9336 4896 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 6999 9367 7057 9373
rect 6999 9333 7011 9367
rect 7045 9364 7057 9367
rect 7650 9364 7656 9376
rect 7045 9336 7656 9364
rect 7045 9333 7057 9336
rect 6999 9327 7057 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 9048 9364 9076 9392
rect 8435 9336 9076 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 11848 9336 12449 9364
rect 11848 9324 11854 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 2096 9132 2145 9160
rect 2096 9120 2102 9132
rect 2133 9129 2145 9132
rect 2179 9129 2191 9163
rect 2133 9123 2191 9129
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2501 9163 2559 9169
rect 2501 9160 2513 9163
rect 2464 9132 2513 9160
rect 2464 9120 2470 9132
rect 2501 9129 2513 9132
rect 2547 9129 2559 9163
rect 2501 9123 2559 9129
rect 3329 9163 3387 9169
rect 3329 9129 3341 9163
rect 3375 9160 3387 9163
rect 3510 9160 3516 9172
rect 3375 9132 3516 9160
rect 3375 9129 3387 9132
rect 3329 9123 3387 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 7282 9160 7288 9172
rect 6687 9132 7288 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7484 9132 8125 9160
rect 2222 9052 2228 9104
rect 2280 9092 2286 9104
rect 3605 9095 3663 9101
rect 3605 9092 3617 9095
rect 2280 9064 3617 9092
rect 2280 9052 2286 9064
rect 3605 9061 3617 9064
rect 3651 9061 3663 9095
rect 3605 9055 3663 9061
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7484 9101 7512 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8113 9123 8171 9129
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8444 9132 8493 9160
rect 8444 9120 8450 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 8481 9123 8539 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9824 9132 10241 9160
rect 9824 9120 9830 9132
rect 10229 9129 10241 9132
rect 10275 9160 10287 9163
rect 10686 9160 10692 9172
rect 10275 9132 10692 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10928 9132 11069 9160
rect 10928 9120 10934 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11057 9123 11115 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11756 9132 11805 9160
rect 11756 9120 11762 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 11793 9123 11851 9129
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 7432 9064 7481 9092
rect 7432 9052 7438 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 7650 9092 7656 9104
rect 7611 9064 7656 9092
rect 7469 9055 7527 9061
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 7745 9095 7803 9101
rect 7745 9061 7757 9095
rect 7791 9092 7803 9095
rect 7926 9092 7932 9104
rect 7791 9064 7932 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11885 9095 11943 9101
rect 11885 9092 11897 9095
rect 11664 9064 11897 9092
rect 11664 9052 11670 9064
rect 11885 9061 11897 9064
rect 11931 9061 11943 9095
rect 11885 9055 11943 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1486 9024 1492 9036
rect 1443 8996 1492 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1486 8984 1492 8996
rect 1544 8984 1550 9036
rect 1946 8984 1952 9036
rect 2004 9024 2010 9036
rect 2314 9024 2320 9036
rect 2004 8996 2320 9024
rect 2004 8984 2010 8996
rect 2314 8984 2320 8996
rect 2372 9024 2378 9036
rect 2685 9027 2743 9033
rect 2685 9024 2697 9027
rect 2372 8996 2697 9024
rect 2372 8984 2378 8996
rect 2685 8993 2697 8996
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 3200 8996 4629 9024
rect 3200 8984 3206 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 4706 9024 4712 9036
rect 4663 8996 4712 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4890 9033 4896 9036
rect 4884 9024 4896 9033
rect 4851 8996 4896 9024
rect 4884 8987 4896 8996
rect 4890 8984 4896 8987
rect 4948 8984 4954 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 7834 9024 7840 9036
rect 7055 8996 7840 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 10008 8996 10333 9024
rect 10008 8984 10014 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 10226 8956 10232 8968
rect 10187 8928 10232 8956
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 2866 8820 2872 8832
rect 2827 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 4798 8820 4804 8832
rect 4571 8792 4804 8820
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 4798 8780 4804 8792
rect 4856 8820 4862 8832
rect 5994 8820 6000 8832
rect 4856 8792 6000 8820
rect 4856 8780 4862 8792
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 7064 8792 7205 8820
rect 7064 8780 7070 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 9490 8820 9496 8832
rect 9451 8792 9496 8820
rect 7193 8783 7251 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9769 8823 9827 8829
rect 9769 8789 9781 8823
rect 9815 8820 9827 8823
rect 10134 8820 10140 8832
rect 9815 8792 10140 8820
rect 9815 8789 9827 8792
rect 9769 8783 9827 8789
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11330 8820 11336 8832
rect 11291 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1820 8588 1961 8616
rect 1820 8576 1826 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 1949 8579 2007 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7708 8588 8217 8616
rect 7708 8576 7714 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 8352 8588 8585 8616
rect 8352 8576 8358 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 8573 8579 8631 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10226 8616 10232 8628
rect 9876 8588 10232 8616
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 2832 8520 3709 8548
rect 2832 8508 2838 8520
rect 3697 8517 3709 8520
rect 3743 8517 3755 8551
rect 3697 8511 3755 8517
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6917 8551 6975 8557
rect 6917 8548 6929 8551
rect 5592 8520 6929 8548
rect 5592 8508 5598 8520
rect 6917 8517 6929 8520
rect 6963 8517 6975 8551
rect 7926 8548 7932 8560
rect 7887 8520 7932 8548
rect 6917 8511 6975 8517
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 9876 8548 9904 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 10928 8588 11253 8616
rect 10928 8576 10934 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11241 8579 11299 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 9447 8520 9904 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 11756 8520 12173 8548
rect 11756 8508 11762 8520
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 4062 8480 4068 8492
rect 4023 8452 4068 8480
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4948 8452 4997 8480
rect 4948 8440 4954 8452
rect 4985 8449 4997 8452
rect 5031 8480 5043 8483
rect 5031 8452 6316 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1762 8412 1768 8424
rect 1443 8384 1768 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 3513 8415 3571 8421
rect 2547 8384 3188 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 3160 8288 3188 8384
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 4246 8412 4252 8424
rect 3559 8384 4252 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5813 8415 5871 8421
rect 5813 8412 5825 8415
rect 5132 8384 5825 8412
rect 5132 8372 5138 8384
rect 5813 8381 5825 8384
rect 5859 8412 5871 8415
rect 5994 8412 6000 8424
rect 5859 8384 6000 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 5534 8344 5540 8356
rect 5495 8316 5540 8344
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5718 8344 5724 8356
rect 5679 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6288 8353 6316 8452
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 7248 8452 7297 8480
rect 7248 8440 7254 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7742 8412 7748 8424
rect 6687 8384 7748 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 8076 8384 8401 8412
rect 8076 8372 8082 8384
rect 8389 8381 8401 8384
rect 8435 8412 8447 8415
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8435 8384 8953 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 9824 8384 9873 8412
rect 9824 8372 9830 8384
rect 9861 8381 9873 8384
rect 9907 8381 9919 8415
rect 9861 8375 9919 8381
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 6319 8316 7481 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7469 8313 7481 8316
rect 7515 8344 7527 8347
rect 9122 8344 9128 8356
rect 7515 8316 9128 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 10106 8347 10164 8353
rect 10106 8344 10118 8347
rect 9548 8316 10118 8344
rect 9548 8304 9554 8316
rect 10106 8313 10118 8316
rect 10152 8344 10164 8347
rect 10962 8344 10968 8356
rect 10152 8316 10968 8344
rect 10152 8313 10164 8316
rect 10106 8307 10164 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 2682 8276 2688 8288
rect 2643 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 4157 8279 4215 8285
rect 4157 8276 4169 8279
rect 3568 8248 4169 8276
rect 3568 8236 3574 8248
rect 4157 8245 4169 8248
rect 4203 8276 4215 8279
rect 5243 8279 5301 8285
rect 5243 8276 5255 8279
rect 4203 8248 5255 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 5243 8245 5255 8248
rect 5289 8245 5301 8279
rect 5243 8239 5301 8245
rect 7377 8279 7435 8285
rect 7377 8245 7389 8279
rect 7423 8276 7435 8279
rect 7742 8276 7748 8288
rect 7423 8248 7748 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 1544 8044 2421 8072
rect 1544 8032 1550 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 3016 8044 3157 8072
rect 3016 8032 3022 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3145 8035 3203 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4246 8072 4252 8084
rect 4207 8044 4252 8072
rect 4246 8032 4252 8044
rect 4304 8072 4310 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 4304 8044 5917 8072
rect 4304 8032 4310 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7190 8072 7196 8084
rect 6963 8044 7196 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11606 8072 11612 8084
rect 11567 8044 11612 8072
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 3050 8004 3056 8016
rect 2915 7976 3056 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 4706 7964 4712 8016
rect 4764 7964 4770 8016
rect 7742 8004 7748 8016
rect 7703 7976 7748 8004
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 9950 8013 9956 8016
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9944 8004 9956 8013
rect 9171 7976 9956 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 9944 7967 9956 7976
rect 9950 7964 9956 7967
rect 10008 7964 10014 8016
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2498 7936 2504 7948
rect 1719 7908 2504 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 2774 7936 2780 7948
rect 2556 7908 2780 7936
rect 2556 7896 2562 7908
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 3844 7908 4537 7936
rect 3844 7896 3850 7908
rect 4525 7905 4537 7908
rect 4571 7936 4583 7939
rect 4724 7936 4752 7964
rect 4571 7908 4752 7936
rect 4792 7939 4850 7945
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4792 7905 4804 7939
rect 4838 7936 4850 7939
rect 5074 7936 5080 7948
rect 4838 7908 5080 7936
rect 4838 7905 4850 7908
rect 4792 7899 4850 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 6696 7908 7573 7936
rect 6696 7896 6702 7908
rect 7561 7905 7573 7908
rect 7607 7936 7619 7939
rect 8202 7936 8208 7948
rect 7607 7908 8208 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9539 7908 9689 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 9677 7905 9689 7908
rect 9723 7936 9735 7939
rect 9766 7936 9772 7948
rect 9723 7908 9772 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9766 7896 9772 7908
rect 9824 7936 9830 7948
rect 10686 7936 10692 7948
rect 9824 7908 10692 7936
rect 9824 7896 9830 7908
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 7834 7868 7840 7880
rect 7795 7840 7840 7868
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 6549 7803 6607 7809
rect 6549 7769 6561 7803
rect 6595 7800 6607 7803
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6595 7772 7297 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 7285 7769 7297 7772
rect 7331 7800 7343 7803
rect 7374 7800 7380 7812
rect 7331 7772 7380 7800
rect 7331 7769 7343 7772
rect 7285 7763 7343 7769
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 8573 7735 8631 7741
rect 8573 7732 8585 7735
rect 8536 7704 8585 7732
rect 8536 7692 8542 7704
rect 8573 7701 8585 7704
rect 8619 7701 8631 7735
rect 8573 7695 8631 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2590 7528 2596 7540
rect 2547 7500 2596 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2516 7324 2544 7491
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3234 7528 3240 7540
rect 2915 7500 3240 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 2976 7333 3004 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3786 7528 3792 7540
rect 3747 7500 3792 7528
rect 3786 7488 3792 7500
rect 3844 7528 3850 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3844 7500 4077 7528
rect 3844 7488 3850 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 4065 7491 4123 7497
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4080 7392 4108 7491
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7800 7500 7849 7528
rect 7800 7488 7806 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 9950 7528 9956 7540
rect 9911 7500 9956 7528
rect 7837 7491 7895 7497
rect 9950 7488 9956 7500
rect 10008 7528 10014 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10008 7500 10885 7528
rect 10008 7488 10014 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 6914 7460 6920 7472
rect 6875 7432 6920 7460
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4080 7364 4261 7392
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 8435 7364 8616 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 1719 7296 2544 7324
rect 2961 7327 3019 7333
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2961 7293 2973 7327
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 4505 7327 4563 7333
rect 4505 7324 4517 7327
rect 4396 7296 4517 7324
rect 4396 7284 4402 7296
rect 4505 7293 4517 7296
rect 4551 7293 4563 7327
rect 4505 7287 4563 7293
rect 6273 7327 6331 7333
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 6319 7296 7481 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 7469 7293 7481 7296
rect 7515 7324 7527 7327
rect 8478 7324 8484 7336
rect 7515 7296 8484 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8588 7333 8616 7364
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7324 8631 7327
rect 9766 7324 9772 7336
rect 8619 7296 9772 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2314 7256 2320 7268
rect 1995 7228 2320 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 7190 7256 7196 7268
rect 7151 7228 7196 7256
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 7374 7256 7380 7268
rect 7335 7228 7380 7256
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 8496 7256 8524 7284
rect 8818 7259 8876 7265
rect 8818 7256 8830 7259
rect 8496 7228 8830 7256
rect 8818 7225 8830 7228
rect 8864 7225 8876 7259
rect 8818 7219 8876 7225
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5592 7160 5641 7188
rect 5592 7148 5598 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 10686 7188 10692 7200
rect 10643 7160 10692 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2498 6984 2504 6996
rect 2459 6956 2504 6984
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5074 6984 5080 6996
rect 5035 6956 5080 6984
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7190 6984 7196 6996
rect 6963 6956 7196 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 8478 6984 8484 6996
rect 8439 6956 8484 6984
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 4246 6876 4252 6928
rect 4304 6916 4310 6928
rect 4617 6919 4675 6925
rect 4617 6916 4629 6919
rect 4304 6888 4629 6916
rect 4304 6876 4310 6888
rect 4617 6885 4629 6888
rect 4663 6885 4675 6919
rect 7368 6919 7426 6925
rect 7368 6916 7380 6919
rect 4617 6879 4675 6885
rect 7300 6888 7380 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6817 1731 6851
rect 1673 6811 1731 6817
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2866 6848 2872 6860
rect 1995 6820 2872 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 1688 6780 1716 6811
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3786 6848 3792 6860
rect 3007 6820 3792 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3786 6808 3792 6820
rect 3844 6848 3850 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 3844 6820 4445 6848
rect 3844 6808 3850 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4580 6820 4721 6848
rect 4580 6808 4586 6820
rect 4709 6817 4721 6820
rect 4755 6848 4767 6851
rect 5442 6848 5448 6860
rect 4755 6820 5448 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5718 6848 5724 6860
rect 5675 6820 5724 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 2038 6780 2044 6792
rect 1688 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5644 6780 5672 6811
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7300 6848 7328 6888
rect 7368 6885 7380 6888
rect 7414 6916 7426 6919
rect 7834 6916 7840 6928
rect 7414 6888 7840 6916
rect 7414 6885 7426 6888
rect 7368 6879 7426 6885
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 10229 6919 10287 6925
rect 10229 6885 10241 6919
rect 10275 6885 10287 6919
rect 10229 6879 10287 6885
rect 10042 6848 10048 6860
rect 6595 6820 7328 6848
rect 10003 6820 10048 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10244 6848 10272 6879
rect 10192 6820 10272 6848
rect 10192 6808 10198 6820
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10962 6848 10968 6860
rect 10376 6820 10968 6848
rect 10376 6808 10382 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 5592 6752 5672 6780
rect 5592 6740 5598 6752
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6880 6752 7113 6780
rect 6880 6740 6886 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 3881 6715 3939 6721
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 4522 6712 4528 6724
rect 3927 6684 4528 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4522 6672 4528 6684
rect 4580 6672 4586 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 5813 6715 5871 6721
rect 5813 6712 5825 6715
rect 5684 6684 5825 6712
rect 5684 6672 5690 6684
rect 5813 6681 5825 6684
rect 5859 6681 5871 6715
rect 5813 6675 5871 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3970 6644 3976 6656
rect 2915 6616 3976 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6086 6644 6092 6656
rect 5583 6616 6092 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 3694 6440 3700 6452
rect 3655 6412 3700 6440
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4246 6440 4252 6452
rect 4203 6412 4252 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7892 6412 8217 6440
rect 7892 6400 7898 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 8205 6403 8263 6409
rect 9324 6412 9873 6440
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 3712 6372 3740 6400
rect 2832 6344 2877 6372
rect 3712 6344 4292 6372
rect 2832 6332 2838 6344
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3200 6276 3249 6304
rect 3200 6264 3206 6276
rect 3237 6273 3249 6276
rect 3283 6304 3295 6307
rect 4154 6304 4160 6316
rect 3283 6276 4160 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4264 6313 4292 6344
rect 9324 6313 9352 6412
rect 9861 6409 9873 6412
rect 9907 6440 9919 6443
rect 10042 6440 10048 6452
rect 9907 6412 10048 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10192 6412 10517 6440
rect 10192 6400 10198 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10229 6375 10287 6381
rect 10229 6341 10241 6375
rect 10275 6372 10287 6375
rect 10318 6372 10324 6384
rect 10275 6344 10324 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 10318 6332 10324 6344
rect 10376 6332 10382 6384
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1854 6236 1860 6248
rect 1443 6208 1860 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 2038 6236 2044 6248
rect 1999 6208 2044 6236
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6236 2651 6239
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 2639 6208 3341 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 3329 6199 3387 6205
rect 3344 6168 3372 6199
rect 4264 6168 4292 6267
rect 4522 6245 4528 6248
rect 4516 6236 4528 6245
rect 4483 6208 4528 6236
rect 4516 6199 4528 6208
rect 4522 6196 4528 6199
rect 4580 6196 4586 6248
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 4632 6208 6561 6236
rect 4632 6168 4660 6208
rect 6549 6205 6561 6208
rect 6595 6236 6607 6239
rect 6822 6236 6828 6248
rect 6595 6208 6828 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 3344 6140 4200 6168
rect 4264 6140 4660 6168
rect 6196 6140 7082 6168
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 3234 6100 3240 6112
rect 3195 6072 3240 6100
rect 1581 6063 1639 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 4172 6100 4200 6140
rect 6196 6109 6224 6140
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 7070 6131 7128 6137
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 4172 6072 5641 6100
rect 5629 6069 5641 6072
rect 5675 6100 5687 6103
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 5675 6072 6193 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 6181 6063 6239 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 1854 5896 1860 5908
rect 1719 5868 1860 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3786 5896 3792 5908
rect 3747 5868 3792 5896
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5592 5868 5641 5896
rect 5592 5856 5598 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 6822 5896 6828 5908
rect 6783 5868 6828 5896
rect 5629 5859 5687 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7190 5896 7196 5908
rect 7055 5868 7196 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7834 5896 7840 5908
rect 7607 5868 7840 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 4706 5828 4712 5840
rect 4667 5800 4712 5828
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2498 5760 2504 5772
rect 1811 5732 2504 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3970 5760 3976 5772
rect 3559 5732 3976 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3970 5720 3976 5732
rect 4028 5760 4034 5772
rect 4522 5760 4528 5772
rect 4028 5732 4528 5760
rect 4028 5720 4034 5732
rect 4522 5720 4528 5732
rect 4580 5760 4586 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4580 5732 4813 5760
rect 4580 5720 4586 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 3234 5624 3240 5636
rect 2823 5596 3240 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 3234 5584 3240 5596
rect 3292 5624 3298 5636
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 3292 5596 4261 5624
rect 3292 5584 3298 5596
rect 4249 5593 4261 5596
rect 4295 5593 4307 5627
rect 4249 5587 4307 5593
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 3970 5352 3976 5364
rect 3931 5324 3976 5352
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4706 5352 4712 5364
rect 4667 5324 4712 5352
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 1995 5188 4108 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 2038 5148 2044 5160
rect 1719 5120 2044 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 4080 5157 4108 5188
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2924 5120 2973 5148
rect 2924 5108 2930 5120
rect 2961 5117 2973 5120
rect 3007 5148 3019 5151
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3007 5120 3525 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4154 5148 4160 5160
rect 4111 5120 4160 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 4246 5012 4252 5024
rect 4207 4984 4252 5012
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4672 4984 4997 5012
rect 4672 4972 4678 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4212 4780 4261 4808
rect 4212 4768 4218 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1946 4672 1952 4684
rect 1443 4644 1952 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2498 4672 2504 4684
rect 2459 4644 2504 4672
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3234 4604 3240 4616
rect 2823 4576 3240 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2038 4468 2044 4480
rect 1999 4440 2044 4468
rect 2038 4428 2044 4440
rect 2096 4428 2102 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1946 4264 1952 4276
rect 1719 4236 1952 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1946 4224 1952 4236
rect 2004 4224 2010 4276
rect 3602 4264 3608 4276
rect 3563 4236 3608 4264
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 2556 4168 2728 4196
rect 2556 4156 2562 4168
rect 2700 4128 2728 4168
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2700 4100 3249 4128
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2148 3924 2176 4023
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 2372 4032 3433 4060
rect 2372 4020 2378 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3467 4032 3985 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 2409 3995 2467 4001
rect 2409 3961 2421 3995
rect 2455 3992 2467 3995
rect 2682 3992 2688 4004
rect 2455 3964 2688 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 2682 3952 2688 3964
rect 2740 3952 2746 4004
rect 2958 3992 2964 4004
rect 2919 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 2976 3924 3004 3952
rect 2148 3896 3004 3924
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1673 3723 1731 3729
rect 1673 3720 1685 3723
rect 1544 3692 1685 3720
rect 1544 3680 1550 3692
rect 1673 3689 1685 3692
rect 1719 3720 1731 3723
rect 2130 3720 2136 3732
rect 1719 3692 2136 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2222 3584 2228 3596
rect 1811 3556 2228 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3234 3176 3240 3188
rect 3195 3148 3240 3176
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1486 2972 1492 2984
rect 1443 2944 1492 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 3234 2972 3240 2984
rect 2731 2944 3240 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 2498 2904 2504 2916
rect 1719 2876 2504 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1964 2496 1992 2592
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 4617 2567 4675 2573
rect 4617 2564 4629 2567
rect 2832 2536 4629 2564
rect 2832 2524 2838 2536
rect 2498 2496 2504 2508
rect 1443 2468 1992 2496
rect 2459 2468 2504 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2498 2456 2504 2468
rect 2556 2496 2562 2508
rect 4080 2505 4108 2536
rect 4617 2533 4629 2536
rect 4663 2533 4675 2567
rect 4617 2527 4675 2533
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 2556 2468 3065 2496
rect 2556 2456 2562 2468
rect 3053 2465 3065 2468
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2682 2292 2688 2304
rect 2643 2264 2688 2292
rect 2682 2252 2688 2264
rect 2740 2252 2746 2304
rect 4246 2292 4252 2304
rect 4207 2264 4252 2292
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 4068 26528 4120 26580
rect 7288 26528 7340 26580
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2044 25440 2096 25492
rect 2688 25440 2740 25492
rect 1584 25372 1636 25424
rect 8208 25372 8260 25424
rect 10232 25372 10284 25424
rect 1768 25347 1820 25356
rect 1768 25313 1777 25347
rect 1777 25313 1811 25347
rect 1811 25313 1820 25347
rect 1768 25304 1820 25313
rect 8300 25304 8352 25356
rect 10140 25304 10192 25356
rect 3424 25236 3476 25288
rect 8576 25279 8628 25288
rect 8576 25245 8585 25279
rect 8585 25245 8619 25279
rect 8619 25245 8628 25279
rect 8576 25236 8628 25245
rect 10416 25279 10468 25288
rect 2780 25168 2832 25220
rect 3056 25168 3108 25220
rect 9404 25168 9456 25220
rect 10416 25245 10425 25279
rect 10425 25245 10459 25279
rect 10459 25245 10468 25279
rect 10416 25236 10468 25245
rect 12808 25236 12860 25288
rect 23664 25168 23716 25220
rect 24308 25168 24360 25220
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 9312 25100 9364 25152
rect 15292 25100 15344 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 848 24896 900 24948
rect 2780 24896 2832 24948
rect 3884 24896 3936 24948
rect 10232 24939 10284 24948
rect 10232 24905 10241 24939
rect 10241 24905 10275 24939
rect 10275 24905 10284 24939
rect 10232 24896 10284 24905
rect 2688 24828 2740 24880
rect 9680 24828 9732 24880
rect 10416 24828 10468 24880
rect 10968 24828 11020 24880
rect 3424 24803 3476 24812
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2596 24556 2648 24608
rect 3424 24769 3433 24803
rect 3433 24769 3467 24803
rect 3467 24769 3476 24803
rect 3424 24760 3476 24769
rect 6000 24760 6052 24812
rect 6552 24760 6604 24812
rect 10140 24760 10192 24812
rect 12992 24828 13044 24880
rect 12900 24760 12952 24812
rect 2780 24667 2832 24676
rect 2780 24633 2789 24667
rect 2789 24633 2823 24667
rect 2823 24633 2832 24667
rect 3056 24667 3108 24676
rect 2780 24624 2832 24633
rect 3056 24633 3065 24667
rect 3065 24633 3099 24667
rect 3099 24633 3108 24667
rect 3056 24624 3108 24633
rect 6092 24692 6144 24744
rect 8116 24735 8168 24744
rect 8116 24701 8125 24735
rect 8125 24701 8159 24735
rect 8159 24701 8168 24735
rect 8116 24692 8168 24701
rect 12440 24692 12492 24744
rect 15568 24692 15620 24744
rect 8300 24624 8352 24676
rect 8944 24667 8996 24676
rect 8944 24633 8953 24667
rect 8953 24633 8987 24667
rect 8987 24633 8996 24667
rect 8944 24624 8996 24633
rect 9312 24624 9364 24676
rect 10048 24624 10100 24676
rect 10692 24667 10744 24676
rect 3884 24599 3936 24608
rect 3884 24565 3893 24599
rect 3893 24565 3927 24599
rect 3927 24565 3936 24599
rect 3884 24556 3936 24565
rect 5540 24556 5592 24608
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 10692 24633 10701 24667
rect 10701 24633 10735 24667
rect 10735 24633 10744 24667
rect 10692 24624 10744 24633
rect 12900 24667 12952 24676
rect 12900 24633 12909 24667
rect 12909 24633 12943 24667
rect 12943 24633 12952 24667
rect 12900 24624 12952 24633
rect 12992 24624 13044 24676
rect 13360 24624 13412 24676
rect 14372 24667 14424 24676
rect 14372 24633 14381 24667
rect 14381 24633 14415 24667
rect 14415 24633 14424 24667
rect 14372 24624 14424 24633
rect 13268 24556 13320 24608
rect 16488 24624 16540 24676
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1768 24352 1820 24404
rect 7564 24352 7616 24404
rect 8024 24352 8076 24404
rect 8576 24395 8628 24404
rect 8576 24361 8585 24395
rect 8585 24361 8619 24395
rect 8619 24361 8628 24395
rect 8576 24352 8628 24361
rect 9404 24395 9456 24404
rect 9404 24361 9413 24395
rect 9413 24361 9447 24395
rect 9447 24361 9456 24395
rect 9404 24352 9456 24361
rect 10140 24395 10192 24404
rect 10140 24361 10149 24395
rect 10149 24361 10183 24395
rect 10183 24361 10192 24395
rect 10140 24352 10192 24361
rect 10692 24352 10744 24404
rect 12440 24352 12492 24404
rect 13268 24352 13320 24404
rect 17040 24352 17092 24404
rect 25412 24352 25464 24404
rect 2872 24284 2924 24336
rect 2504 24259 2556 24268
rect 2504 24225 2529 24259
rect 2529 24225 2556 24259
rect 2504 24216 2556 24225
rect 6184 24284 6236 24336
rect 11612 24327 11664 24336
rect 11612 24293 11621 24327
rect 11621 24293 11655 24327
rect 11655 24293 11664 24327
rect 11612 24284 11664 24293
rect 6644 24216 6696 24268
rect 2780 24148 2832 24200
rect 3056 24191 3108 24200
rect 3056 24157 3065 24191
rect 3065 24157 3099 24191
rect 3099 24157 3108 24191
rect 3056 24148 3108 24157
rect 3424 24148 3476 24200
rect 4252 24148 4304 24200
rect 11520 24191 11572 24200
rect 11520 24157 11529 24191
rect 11529 24157 11563 24191
rect 11563 24157 11572 24191
rect 11520 24148 11572 24157
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 2412 24080 2464 24132
rect 6920 24080 6972 24132
rect 7748 24080 7800 24132
rect 21916 24327 21968 24336
rect 21916 24293 21950 24327
rect 21950 24293 21968 24327
rect 21916 24284 21968 24293
rect 12440 24216 12492 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16580 24259 16632 24268
rect 16580 24225 16589 24259
rect 16589 24225 16623 24259
rect 16623 24225 16632 24259
rect 16580 24216 16632 24225
rect 24032 24216 24084 24268
rect 21640 24191 21692 24200
rect 2320 24055 2372 24064
rect 2320 24021 2329 24055
rect 2329 24021 2363 24055
rect 2363 24021 2372 24055
rect 2320 24012 2372 24021
rect 2780 24012 2832 24064
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 4160 24012 4212 24064
rect 5356 24012 5408 24064
rect 8944 24012 8996 24064
rect 9864 24012 9916 24064
rect 21640 24157 21649 24191
rect 21649 24157 21683 24191
rect 21683 24157 21692 24191
rect 21640 24148 21692 24157
rect 23020 24123 23072 24132
rect 23020 24089 23029 24123
rect 23029 24089 23063 24123
rect 23063 24089 23072 24123
rect 23020 24080 23072 24089
rect 13452 24012 13504 24064
rect 23940 24055 23992 24064
rect 23940 24021 23949 24055
rect 23949 24021 23983 24055
rect 23983 24021 23992 24055
rect 23940 24012 23992 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2872 23808 2924 23860
rect 3516 23808 3568 23860
rect 8852 23808 8904 23860
rect 10140 23808 10192 23860
rect 11612 23808 11664 23860
rect 11704 23808 11756 23860
rect 13360 23808 13412 23860
rect 16580 23851 16632 23860
rect 16580 23817 16589 23851
rect 16589 23817 16623 23851
rect 16623 23817 16632 23851
rect 16580 23808 16632 23817
rect 21916 23808 21968 23860
rect 24124 23851 24176 23860
rect 24124 23817 24133 23851
rect 24133 23817 24167 23851
rect 24167 23817 24176 23851
rect 24124 23808 24176 23817
rect 26516 23808 26568 23860
rect 5448 23740 5500 23792
rect 6828 23740 6880 23792
rect 15936 23740 15988 23792
rect 1768 23672 1820 23724
rect 5356 23672 5408 23724
rect 6276 23672 6328 23724
rect 7380 23715 7432 23724
rect 7380 23681 7389 23715
rect 7389 23681 7423 23715
rect 7423 23681 7432 23715
rect 7380 23672 7432 23681
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 1676 23468 1728 23520
rect 3976 23604 4028 23656
rect 5540 23647 5592 23656
rect 5540 23613 5549 23647
rect 5549 23613 5583 23647
rect 5583 23613 5592 23647
rect 5540 23604 5592 23613
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 9220 23604 9272 23613
rect 3424 23536 3476 23588
rect 6184 23579 6236 23588
rect 6184 23545 6193 23579
rect 6193 23545 6227 23579
rect 6227 23545 6236 23579
rect 6184 23536 6236 23545
rect 9312 23536 9364 23588
rect 16028 23604 16080 23656
rect 16856 23647 16908 23656
rect 16856 23613 16865 23647
rect 16865 23613 16899 23647
rect 16899 23613 16908 23647
rect 16856 23604 16908 23613
rect 23480 23604 23532 23656
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24860 23604 24912 23656
rect 13452 23536 13504 23588
rect 16488 23536 16540 23588
rect 23572 23536 23624 23588
rect 24032 23536 24084 23588
rect 5356 23468 5408 23520
rect 6644 23511 6696 23520
rect 6644 23477 6653 23511
rect 6653 23477 6687 23511
rect 6687 23477 6696 23511
rect 6644 23468 6696 23477
rect 6920 23468 6972 23520
rect 11704 23468 11756 23520
rect 12716 23468 12768 23520
rect 12992 23511 13044 23520
rect 12992 23477 13001 23511
rect 13001 23477 13035 23511
rect 13035 23477 13044 23511
rect 12992 23468 13044 23477
rect 15292 23511 15344 23520
rect 15292 23477 15301 23511
rect 15301 23477 15335 23511
rect 15335 23477 15344 23511
rect 15292 23468 15344 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2412 23264 2464 23316
rect 2596 23264 2648 23316
rect 6000 23264 6052 23316
rect 6828 23264 6880 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12348 23264 12400 23316
rect 17592 23264 17644 23316
rect 17868 23307 17920 23316
rect 17868 23273 17877 23307
rect 17877 23273 17911 23307
rect 17911 23273 17920 23307
rect 17868 23264 17920 23273
rect 19064 23307 19116 23316
rect 19064 23273 19073 23307
rect 19073 23273 19107 23307
rect 19107 23273 19116 23307
rect 19064 23264 19116 23273
rect 3056 23196 3108 23248
rect 3516 23196 3568 23248
rect 6276 23196 6328 23248
rect 3976 23128 4028 23180
rect 5080 23128 5132 23180
rect 10140 23196 10192 23248
rect 15568 23239 15620 23248
rect 15568 23205 15577 23239
rect 15577 23205 15611 23239
rect 15611 23205 15620 23239
rect 15568 23196 15620 23205
rect 23480 23196 23532 23248
rect 24768 23196 24820 23248
rect 9220 23128 9272 23180
rect 10968 23128 11020 23180
rect 12716 23128 12768 23180
rect 15384 23128 15436 23180
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17684 23171 17736 23180
rect 17684 23137 17693 23171
rect 17693 23137 17727 23171
rect 17727 23137 17736 23171
rect 17684 23128 17736 23137
rect 18788 23128 18840 23180
rect 22100 23128 22152 23180
rect 23756 23128 23808 23180
rect 6184 23060 6236 23112
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 1584 22924 1636 22976
rect 2780 22967 2832 22976
rect 2780 22933 2789 22967
rect 2789 22933 2823 22967
rect 2823 22933 2832 22967
rect 3424 22967 3476 22976
rect 2780 22924 2832 22933
rect 3424 22933 3433 22967
rect 3433 22933 3467 22967
rect 3467 22933 3476 22967
rect 3424 22924 3476 22933
rect 7932 22967 7984 22976
rect 7932 22933 7941 22967
rect 7941 22933 7975 22967
rect 7975 22933 7984 22967
rect 7932 22924 7984 22933
rect 9312 22967 9364 22976
rect 9312 22933 9321 22967
rect 9321 22933 9355 22967
rect 9355 22933 9364 22967
rect 9312 22924 9364 22933
rect 13452 22924 13504 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2780 22720 2832 22772
rect 3608 22763 3660 22772
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 3056 22627 3108 22636
rect 3056 22593 3065 22627
rect 3065 22593 3099 22627
rect 3099 22593 3108 22627
rect 3056 22584 3108 22593
rect 3608 22729 3617 22763
rect 3617 22729 3651 22763
rect 3651 22729 3660 22763
rect 3608 22720 3660 22729
rect 3976 22720 4028 22772
rect 5172 22720 5224 22772
rect 6184 22720 6236 22772
rect 7380 22720 7432 22772
rect 9220 22763 9272 22772
rect 9220 22729 9229 22763
rect 9229 22729 9263 22763
rect 9263 22729 9272 22763
rect 9220 22720 9272 22729
rect 13360 22763 13412 22772
rect 13360 22729 13369 22763
rect 13369 22729 13403 22763
rect 13403 22729 13412 22763
rect 13360 22720 13412 22729
rect 15384 22720 15436 22772
rect 16580 22720 16632 22772
rect 18696 22720 18748 22772
rect 19524 22720 19576 22772
rect 7104 22652 7156 22704
rect 8208 22652 8260 22704
rect 5080 22627 5132 22636
rect 5080 22593 5089 22627
rect 5089 22593 5123 22627
rect 5123 22593 5132 22627
rect 5080 22584 5132 22593
rect 7932 22584 7984 22636
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 7104 22516 7156 22568
rect 7472 22559 7524 22568
rect 7472 22525 7481 22559
rect 7481 22525 7515 22559
rect 7515 22525 7524 22559
rect 7472 22516 7524 22525
rect 9588 22559 9640 22568
rect 9588 22525 9622 22559
rect 9622 22525 9640 22559
rect 2596 22491 2648 22500
rect 2596 22457 2605 22491
rect 2605 22457 2639 22491
rect 2639 22457 2648 22491
rect 2596 22448 2648 22457
rect 3884 22491 3936 22500
rect 3884 22457 3893 22491
rect 3893 22457 3927 22491
rect 3927 22457 3936 22491
rect 3884 22448 3936 22457
rect 4068 22491 4120 22500
rect 4068 22457 4077 22491
rect 4077 22457 4111 22491
rect 4111 22457 4120 22491
rect 4068 22448 4120 22457
rect 6276 22491 6328 22500
rect 6276 22457 6285 22491
rect 6285 22457 6319 22491
rect 6319 22457 6328 22491
rect 7380 22491 7432 22500
rect 6276 22448 6328 22457
rect 7380 22457 7389 22491
rect 7389 22457 7423 22491
rect 7423 22457 7432 22491
rect 7380 22448 7432 22457
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 2412 22380 2464 22432
rect 6000 22380 6052 22432
rect 9588 22516 9640 22525
rect 10140 22516 10192 22568
rect 23572 22584 23624 22636
rect 10968 22448 11020 22500
rect 12164 22448 12216 22500
rect 12992 22448 13044 22500
rect 17868 22516 17920 22568
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 16672 22448 16724 22500
rect 17684 22491 17736 22500
rect 17684 22457 17693 22491
rect 17693 22457 17727 22491
rect 17727 22457 17736 22491
rect 17684 22448 17736 22457
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 13268 22380 13320 22432
rect 13544 22380 13596 22432
rect 16212 22423 16264 22432
rect 16212 22389 16221 22423
rect 16221 22389 16255 22423
rect 16255 22389 16264 22423
rect 16212 22380 16264 22389
rect 17776 22380 17828 22432
rect 18788 22380 18840 22432
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 22100 22380 22152 22389
rect 23848 22423 23900 22432
rect 23848 22389 23857 22423
rect 23857 22389 23891 22423
rect 23891 22389 23900 22423
rect 23848 22380 23900 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2136 22176 2188 22228
rect 2596 22176 2648 22228
rect 3148 22176 3200 22228
rect 3976 22176 4028 22228
rect 5080 22176 5132 22228
rect 1492 22108 1544 22160
rect 5540 22108 5592 22160
rect 6828 22176 6880 22228
rect 7656 22176 7708 22228
rect 9588 22176 9640 22228
rect 7196 22151 7248 22160
rect 7196 22117 7205 22151
rect 7205 22117 7239 22151
rect 7239 22117 7248 22151
rect 7196 22108 7248 22117
rect 2136 22040 2188 22092
rect 5448 22040 5500 22092
rect 2688 21972 2740 22024
rect 2504 21947 2556 21956
rect 2504 21913 2513 21947
rect 2513 21913 2547 21947
rect 2547 21913 2556 21947
rect 2504 21904 2556 21913
rect 2596 21904 2648 21956
rect 4252 21972 4304 22024
rect 4620 21972 4672 22024
rect 6644 22040 6696 22092
rect 7472 22083 7524 22092
rect 7472 22049 7481 22083
rect 7481 22049 7515 22083
rect 7515 22049 7524 22083
rect 7472 22040 7524 22049
rect 7564 22040 7616 22092
rect 8852 22108 8904 22160
rect 9496 22108 9548 22160
rect 14556 22176 14608 22228
rect 9312 22040 9364 22092
rect 5724 21972 5776 22024
rect 10140 22015 10192 22024
rect 3148 21904 3200 21956
rect 5356 21947 5408 21956
rect 5356 21913 5365 21947
rect 5365 21913 5399 21947
rect 5399 21913 5408 21947
rect 5356 21904 5408 21913
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 11888 22040 11940 22092
rect 14004 22108 14056 22160
rect 16212 22108 16264 22160
rect 12716 22040 12768 22092
rect 13728 22040 13780 22092
rect 15476 22083 15528 22092
rect 15476 22049 15485 22083
rect 15485 22049 15519 22083
rect 15519 22049 15528 22083
rect 15476 22040 15528 22049
rect 6092 21904 6144 21956
rect 6920 21947 6972 21956
rect 6920 21913 6929 21947
rect 6929 21913 6963 21947
rect 6963 21913 6972 21947
rect 6920 21904 6972 21913
rect 10048 21904 10100 21956
rect 1860 21879 1912 21888
rect 1860 21845 1869 21879
rect 1869 21845 1903 21879
rect 1903 21845 1912 21879
rect 1860 21836 1912 21845
rect 2872 21836 2924 21888
rect 4436 21836 4488 21888
rect 4988 21836 5040 21888
rect 5172 21879 5224 21888
rect 5172 21845 5181 21879
rect 5181 21845 5215 21879
rect 5215 21845 5224 21879
rect 5172 21836 5224 21845
rect 6736 21879 6788 21888
rect 6736 21845 6745 21879
rect 6745 21845 6779 21879
rect 6779 21845 6788 21879
rect 6736 21836 6788 21845
rect 7380 21836 7432 21888
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 11704 21972 11756 22024
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 13360 21972 13412 22024
rect 17868 22040 17920 22092
rect 19340 22083 19392 22092
rect 17132 21972 17184 22024
rect 17776 21972 17828 22024
rect 19340 22049 19349 22083
rect 19349 22049 19383 22083
rect 19383 22049 19392 22083
rect 19340 22040 19392 22049
rect 12348 21904 12400 21956
rect 12992 21904 13044 21956
rect 20352 21904 20404 21956
rect 13544 21836 13596 21888
rect 14648 21879 14700 21888
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2136 21675 2188 21684
rect 2136 21641 2145 21675
rect 2145 21641 2179 21675
rect 2179 21641 2188 21675
rect 2136 21632 2188 21641
rect 3792 21632 3844 21684
rect 4528 21632 4580 21684
rect 4620 21607 4672 21616
rect 4620 21573 4629 21607
rect 4629 21573 4663 21607
rect 4663 21573 4672 21607
rect 4620 21564 4672 21573
rect 4988 21632 5040 21684
rect 6092 21675 6144 21684
rect 5448 21564 5500 21616
rect 6092 21641 6101 21675
rect 6101 21641 6135 21675
rect 6135 21641 6144 21675
rect 6092 21632 6144 21641
rect 6828 21632 6880 21684
rect 7196 21632 7248 21684
rect 7656 21632 7708 21684
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 11704 21675 11756 21684
rect 11704 21641 11713 21675
rect 11713 21641 11747 21675
rect 11747 21641 11756 21675
rect 11704 21632 11756 21641
rect 12900 21632 12952 21684
rect 15476 21675 15528 21684
rect 15476 21641 15485 21675
rect 15485 21641 15519 21675
rect 15519 21641 15528 21675
rect 15476 21632 15528 21641
rect 19984 21632 20036 21684
rect 20628 21675 20680 21684
rect 20628 21641 20637 21675
rect 20637 21641 20671 21675
rect 20671 21641 20680 21675
rect 20628 21632 20680 21641
rect 6920 21607 6972 21616
rect 6920 21573 6929 21607
rect 6929 21573 6963 21607
rect 6963 21573 6972 21607
rect 6920 21564 6972 21573
rect 8484 21607 8536 21616
rect 8484 21573 8493 21607
rect 8493 21573 8527 21607
rect 8527 21573 8536 21607
rect 8484 21564 8536 21573
rect 10140 21564 10192 21616
rect 12716 21564 12768 21616
rect 15016 21564 15068 21616
rect 19340 21564 19392 21616
rect 6736 21496 6788 21548
rect 7104 21496 7156 21548
rect 8944 21496 8996 21548
rect 10692 21496 10744 21548
rect 12900 21496 12952 21548
rect 13452 21496 13504 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 19156 21496 19208 21548
rect 1492 21360 1544 21412
rect 5172 21428 5224 21480
rect 5724 21471 5776 21480
rect 5724 21437 5733 21471
rect 5733 21437 5767 21471
rect 5767 21437 5776 21471
rect 5724 21428 5776 21437
rect 7564 21428 7616 21480
rect 9864 21428 9916 21480
rect 12808 21471 12860 21480
rect 2872 21403 2924 21412
rect 2872 21369 2906 21403
rect 2906 21369 2924 21403
rect 2872 21360 2924 21369
rect 5264 21360 5316 21412
rect 6000 21360 6052 21412
rect 7380 21403 7432 21412
rect 7380 21369 7389 21403
rect 7389 21369 7423 21403
rect 7423 21369 7432 21403
rect 7380 21360 7432 21369
rect 8484 21360 8536 21412
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 14004 21428 14056 21480
rect 12992 21403 13044 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 8852 21292 8904 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 12992 21369 13001 21403
rect 13001 21369 13035 21403
rect 13035 21369 13044 21403
rect 12992 21360 13044 21369
rect 14096 21360 14148 21412
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 20444 21471 20496 21480
rect 20444 21437 20453 21471
rect 20453 21437 20487 21471
rect 20487 21437 20496 21471
rect 20444 21428 20496 21437
rect 9772 21292 9824 21301
rect 11704 21292 11756 21344
rect 11888 21292 11940 21344
rect 13360 21292 13412 21344
rect 14556 21335 14608 21344
rect 14556 21301 14565 21335
rect 14565 21301 14599 21335
rect 14599 21301 14608 21335
rect 14556 21292 14608 21301
rect 15108 21335 15160 21344
rect 15108 21301 15117 21335
rect 15117 21301 15151 21335
rect 15151 21301 15160 21335
rect 15108 21292 15160 21301
rect 17776 21335 17828 21344
rect 17776 21301 17785 21335
rect 17785 21301 17819 21335
rect 17819 21301 17828 21335
rect 17776 21292 17828 21301
rect 19340 21292 19392 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2872 21131 2924 21140
rect 2872 21097 2881 21131
rect 2881 21097 2915 21131
rect 2915 21097 2924 21131
rect 2872 21088 2924 21097
rect 1860 21020 1912 21072
rect 4988 21088 5040 21140
rect 5264 21088 5316 21140
rect 5540 21131 5592 21140
rect 5540 21097 5549 21131
rect 5549 21097 5583 21131
rect 5583 21097 5592 21131
rect 5540 21088 5592 21097
rect 7104 21131 7156 21140
rect 7104 21097 7113 21131
rect 7113 21097 7147 21131
rect 7147 21097 7156 21131
rect 7104 21088 7156 21097
rect 7564 21088 7616 21140
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 9312 21088 9364 21140
rect 9864 21088 9916 21140
rect 10048 21088 10100 21140
rect 12808 21088 12860 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 4528 21020 4580 21072
rect 5724 21020 5776 21072
rect 10692 21020 10744 21072
rect 10968 21020 11020 21072
rect 12992 21020 13044 21072
rect 15016 21131 15068 21140
rect 15016 21097 15025 21131
rect 15025 21097 15059 21131
rect 15059 21097 15068 21131
rect 15016 21088 15068 21097
rect 21088 21131 21140 21140
rect 21088 21097 21097 21131
rect 21097 21097 21131 21131
rect 21131 21097 21140 21131
rect 21088 21088 21140 21097
rect 13268 21020 13320 21072
rect 17500 21063 17552 21072
rect 17500 21029 17509 21063
rect 17509 21029 17543 21063
rect 17543 21029 17552 21063
rect 17500 21020 17552 21029
rect 18788 21063 18840 21072
rect 18788 21029 18797 21063
rect 18797 21029 18831 21063
rect 18831 21029 18840 21063
rect 18788 21020 18840 21029
rect 13820 20952 13872 21004
rect 15476 20952 15528 21004
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 1492 20927 1544 20936
rect 1492 20893 1501 20927
rect 1501 20893 1535 20927
rect 1535 20893 1544 20927
rect 1492 20884 1544 20893
rect 4160 20859 4212 20868
rect 4160 20825 4169 20859
rect 4169 20825 4203 20859
rect 4203 20825 4212 20859
rect 4160 20816 4212 20825
rect 12440 20884 12492 20936
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 17040 20884 17092 20936
rect 12532 20816 12584 20868
rect 13268 20816 13320 20868
rect 19064 20952 19116 21004
rect 21088 20952 21140 21004
rect 6644 20748 6696 20800
rect 8300 20748 8352 20800
rect 8852 20748 8904 20800
rect 12348 20748 12400 20800
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 14556 20791 14608 20800
rect 14556 20757 14565 20791
rect 14565 20757 14599 20791
rect 14599 20757 14608 20791
rect 14556 20748 14608 20757
rect 15292 20748 15344 20800
rect 17960 20748 18012 20800
rect 18696 20748 18748 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 2596 20544 2648 20596
rect 4988 20544 5040 20596
rect 5540 20544 5592 20596
rect 10692 20587 10744 20596
rect 10692 20553 10701 20587
rect 10701 20553 10735 20587
rect 10735 20553 10744 20587
rect 10692 20544 10744 20553
rect 11060 20544 11112 20596
rect 4252 20476 4304 20528
rect 12440 20544 12492 20596
rect 13820 20544 13872 20596
rect 16028 20544 16080 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 19064 20587 19116 20596
rect 19064 20553 19073 20587
rect 19073 20553 19107 20587
rect 19107 20553 19116 20587
rect 19064 20544 19116 20553
rect 2688 20408 2740 20460
rect 9312 20451 9364 20460
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 1676 20272 1728 20324
rect 3792 20272 3844 20324
rect 7104 20383 7156 20392
rect 7104 20349 7138 20383
rect 7138 20349 7156 20383
rect 6644 20315 6696 20324
rect 6644 20281 6653 20315
rect 6653 20281 6687 20315
rect 6687 20281 6696 20315
rect 7104 20340 7156 20349
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 12348 20340 12400 20392
rect 16212 20340 16264 20392
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 19340 20408 19392 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 6644 20272 6696 20281
rect 8944 20272 8996 20324
rect 9404 20272 9456 20324
rect 12532 20272 12584 20324
rect 14648 20272 14700 20324
rect 15384 20315 15436 20324
rect 15384 20281 15396 20315
rect 15396 20281 15436 20315
rect 15384 20272 15436 20281
rect 8116 20204 8168 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 18604 20247 18656 20256
rect 17776 20204 17828 20213
rect 18604 20213 18613 20247
rect 18613 20213 18647 20247
rect 18647 20213 18656 20247
rect 18604 20204 18656 20213
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2320 20000 2372 20052
rect 2504 20000 2556 20052
rect 3516 20043 3568 20052
rect 2688 19975 2740 19984
rect 2688 19941 2697 19975
rect 2697 19941 2731 19975
rect 2731 19941 2740 19975
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 4528 19975 4580 19984
rect 2688 19932 2740 19941
rect 4528 19941 4537 19975
rect 4537 19941 4571 19975
rect 4571 19941 4580 19975
rect 4528 19932 4580 19941
rect 4988 19932 5040 19984
rect 5540 19975 5592 19984
rect 5540 19941 5549 19975
rect 5549 19941 5583 19975
rect 5583 19941 5592 19975
rect 5540 19932 5592 19941
rect 7104 20000 7156 20052
rect 7656 20000 7708 20052
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 12532 20043 12584 20052
rect 12532 20009 12541 20043
rect 12541 20009 12575 20043
rect 12575 20009 12584 20043
rect 12532 20000 12584 20009
rect 13728 20000 13780 20052
rect 14648 20000 14700 20052
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 17960 20000 18012 20052
rect 18604 20000 18656 20052
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 23388 20000 23440 20052
rect 11704 19975 11756 19984
rect 11704 19941 11713 19975
rect 11713 19941 11747 19975
rect 11747 19941 11756 19975
rect 11704 19932 11756 19941
rect 1860 19864 1912 19916
rect 5448 19864 5500 19916
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 13820 19932 13872 19984
rect 16028 19932 16080 19984
rect 16580 19932 16632 19984
rect 18144 19975 18196 19984
rect 18144 19941 18153 19975
rect 18153 19941 18187 19975
rect 18187 19941 18196 19975
rect 18144 19932 18196 19941
rect 20444 19932 20496 19984
rect 19064 19907 19116 19916
rect 19064 19873 19073 19907
rect 19073 19873 19107 19907
rect 19107 19873 19116 19907
rect 19064 19864 19116 19873
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 22836 19864 22888 19916
rect 5172 19796 5224 19848
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 8116 19839 8168 19848
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 10508 19796 10560 19848
rect 12164 19796 12216 19848
rect 12348 19796 12400 19848
rect 12716 19839 12768 19848
rect 12716 19805 12725 19839
rect 12725 19805 12759 19839
rect 12759 19805 12768 19839
rect 12716 19796 12768 19805
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 2596 19728 2648 19780
rect 3148 19728 3200 19780
rect 5816 19771 5868 19780
rect 5816 19737 5825 19771
rect 5825 19737 5859 19771
rect 5859 19737 5868 19771
rect 5816 19728 5868 19737
rect 8208 19728 8260 19780
rect 1492 19660 1544 19712
rect 1952 19660 2004 19712
rect 5080 19660 5132 19712
rect 12992 19660 13044 19712
rect 15476 19703 15528 19712
rect 15476 19669 15485 19703
rect 15485 19669 15519 19703
rect 15519 19669 15528 19703
rect 15476 19660 15528 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4988 19456 5040 19508
rect 6368 19456 6420 19508
rect 7932 19456 7984 19508
rect 9404 19456 9456 19508
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 11520 19456 11572 19508
rect 15384 19499 15436 19508
rect 15384 19465 15393 19499
rect 15393 19465 15427 19499
rect 15427 19465 15436 19499
rect 15384 19456 15436 19465
rect 21088 19456 21140 19508
rect 4528 19388 4580 19440
rect 8116 19388 8168 19440
rect 1952 19320 2004 19372
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 12716 19320 12768 19372
rect 17776 19320 17828 19372
rect 19064 19320 19116 19372
rect 2688 19252 2740 19304
rect 5448 19252 5500 19304
rect 10140 19295 10192 19304
rect 5172 19227 5224 19236
rect 5172 19193 5181 19227
rect 5181 19193 5215 19227
rect 5215 19193 5224 19227
rect 5172 19184 5224 19193
rect 6000 19184 6052 19236
rect 7196 19184 7248 19236
rect 1860 19159 1912 19168
rect 1860 19125 1869 19159
rect 1869 19125 1903 19159
rect 1903 19125 1912 19159
rect 1860 19116 1912 19125
rect 3792 19116 3844 19168
rect 4160 19116 4212 19168
rect 10140 19261 10149 19295
rect 10149 19261 10183 19295
rect 10183 19261 10192 19295
rect 10140 19252 10192 19261
rect 10508 19252 10560 19304
rect 11336 19295 11388 19304
rect 11336 19261 11345 19295
rect 11345 19261 11379 19295
rect 11379 19261 11388 19295
rect 11336 19252 11388 19261
rect 12348 19252 12400 19304
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 13728 19252 13780 19304
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 13912 19252 13964 19261
rect 16580 19295 16632 19304
rect 8300 19184 8352 19236
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 16212 19184 16264 19236
rect 17776 19184 17828 19236
rect 18144 19252 18196 19304
rect 18420 19184 18472 19236
rect 9496 19116 9548 19168
rect 10968 19116 11020 19168
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 18696 19116 18748 19168
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 22192 19116 22244 19168
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2596 18955 2648 18964
rect 2596 18921 2605 18955
rect 2605 18921 2639 18955
rect 2639 18921 2648 18955
rect 2596 18912 2648 18921
rect 5540 18912 5592 18964
rect 6368 18912 6420 18964
rect 8208 18912 8260 18964
rect 11336 18912 11388 18964
rect 12164 18912 12216 18964
rect 19156 18955 19208 18964
rect 19156 18921 19165 18955
rect 19165 18921 19199 18955
rect 19199 18921 19208 18955
rect 19156 18912 19208 18921
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 1584 18844 1636 18896
rect 2688 18844 2740 18896
rect 4620 18887 4672 18896
rect 4620 18853 4654 18887
rect 4654 18853 4672 18887
rect 4620 18844 4672 18853
rect 7932 18844 7984 18896
rect 2044 18776 2096 18828
rect 2872 18776 2924 18828
rect 3240 18776 3292 18828
rect 4988 18776 5040 18828
rect 7196 18819 7248 18828
rect 7196 18785 7205 18819
rect 7205 18785 7239 18819
rect 7239 18785 7248 18819
rect 7196 18776 7248 18785
rect 9036 18776 9088 18828
rect 3792 18708 3844 18760
rect 7472 18751 7524 18760
rect 7472 18717 7481 18751
rect 7481 18717 7515 18751
rect 7515 18717 7524 18751
rect 7472 18708 7524 18717
rect 2136 18683 2188 18692
rect 2136 18649 2145 18683
rect 2145 18649 2179 18683
rect 2179 18649 2188 18683
rect 2136 18640 2188 18649
rect 6920 18683 6972 18692
rect 6920 18649 6929 18683
rect 6929 18649 6963 18683
rect 6963 18649 6972 18683
rect 6920 18640 6972 18649
rect 9772 18683 9824 18692
rect 9772 18649 9781 18683
rect 9781 18649 9815 18683
rect 9815 18649 9824 18683
rect 9772 18640 9824 18649
rect 3148 18615 3200 18624
rect 3148 18581 3157 18615
rect 3157 18581 3191 18615
rect 3191 18581 3200 18615
rect 3148 18572 3200 18581
rect 3240 18572 3292 18624
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 6000 18572 6052 18624
rect 6736 18615 6788 18624
rect 6736 18581 6745 18615
rect 6745 18581 6779 18615
rect 6779 18581 6788 18615
rect 6736 18572 6788 18581
rect 7656 18572 7708 18624
rect 8116 18572 8168 18624
rect 8300 18572 8352 18624
rect 11704 18844 11756 18896
rect 12256 18844 12308 18896
rect 11796 18776 11848 18828
rect 11060 18708 11112 18760
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 15292 18844 15344 18896
rect 15936 18844 15988 18896
rect 18328 18844 18380 18896
rect 18696 18844 18748 18896
rect 21088 18844 21140 18896
rect 13176 18776 13228 18828
rect 15568 18776 15620 18828
rect 17776 18819 17828 18828
rect 17776 18785 17785 18819
rect 17785 18785 17819 18819
rect 17819 18785 17828 18819
rect 17776 18776 17828 18785
rect 20904 18819 20956 18828
rect 20904 18785 20913 18819
rect 20913 18785 20947 18819
rect 20947 18785 20956 18819
rect 20904 18776 20956 18785
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 14004 18751 14056 18760
rect 14004 18717 14013 18751
rect 14013 18717 14047 18751
rect 14047 18717 14056 18751
rect 14004 18708 14056 18717
rect 15292 18708 15344 18760
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 16672 18640 16724 18649
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 4620 18368 4672 18420
rect 5264 18368 5316 18420
rect 6000 18368 6052 18420
rect 7196 18368 7248 18420
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 13176 18411 13228 18420
rect 1952 18300 2004 18352
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 2964 18164 3016 18216
rect 5080 18232 5132 18284
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 12992 18232 13044 18284
rect 13912 18368 13964 18420
rect 15292 18368 15344 18420
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16212 18411 16264 18420
rect 16212 18377 16221 18411
rect 16221 18377 16255 18411
rect 16255 18377 16264 18411
rect 16212 18368 16264 18377
rect 17776 18411 17828 18420
rect 17776 18377 17785 18411
rect 17785 18377 17819 18411
rect 17819 18377 17828 18411
rect 17776 18368 17828 18377
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 22836 18232 22888 18284
rect 3148 18207 3200 18216
rect 3148 18173 3157 18207
rect 3157 18173 3191 18207
rect 3191 18173 3200 18207
rect 3148 18164 3200 18173
rect 3240 18096 3292 18148
rect 3792 18096 3844 18148
rect 4160 18096 4212 18148
rect 1860 18028 1912 18080
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 6644 18164 6696 18216
rect 21272 18207 21324 18216
rect 6736 18096 6788 18148
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 9588 18096 9640 18148
rect 14004 18096 14056 18148
rect 15292 18096 15344 18148
rect 16304 18096 16356 18148
rect 16672 18139 16724 18148
rect 16672 18105 16681 18139
rect 16681 18105 16715 18139
rect 16715 18105 16724 18139
rect 16672 18096 16724 18105
rect 16764 18139 16816 18148
rect 16764 18105 16773 18139
rect 16773 18105 16807 18139
rect 16807 18105 16816 18139
rect 16764 18096 16816 18105
rect 5080 18028 5132 18037
rect 7472 18028 7524 18080
rect 9496 18028 9548 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 11060 18028 11112 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 22100 18028 22152 18080
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2780 17824 2832 17876
rect 4160 17824 4212 17876
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 7472 17824 7524 17876
rect 1952 17756 2004 17808
rect 2964 17756 3016 17808
rect 2412 17688 2464 17740
rect 5356 17756 5408 17808
rect 5540 17756 5592 17808
rect 7012 17756 7064 17808
rect 9128 17824 9180 17876
rect 9588 17824 9640 17876
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 12440 17824 12492 17876
rect 14648 17824 14700 17876
rect 15200 17824 15252 17876
rect 16764 17824 16816 17876
rect 22008 17799 22060 17808
rect 22008 17765 22017 17799
rect 22017 17765 22051 17799
rect 22051 17765 22060 17799
rect 22008 17756 22060 17765
rect 6460 17688 6512 17740
rect 6736 17688 6788 17740
rect 9588 17688 9640 17740
rect 9956 17731 10008 17740
rect 9956 17697 9990 17731
rect 9990 17697 10008 17731
rect 9956 17688 10008 17697
rect 11520 17688 11572 17740
rect 15384 17688 15436 17740
rect 16120 17688 16172 17740
rect 21732 17731 21784 17740
rect 21732 17697 21741 17731
rect 21741 17697 21775 17731
rect 21775 17697 21784 17731
rect 21732 17688 21784 17697
rect 5080 17620 5132 17672
rect 7380 17620 7432 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 2872 17552 2924 17604
rect 7932 17595 7984 17604
rect 7932 17561 7941 17595
rect 7941 17561 7975 17595
rect 7975 17561 7984 17595
rect 7932 17552 7984 17561
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 14004 17484 14056 17536
rect 18604 17484 18656 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 3148 17280 3200 17332
rect 5080 17280 5132 17332
rect 5540 17280 5592 17332
rect 6460 17323 6512 17332
rect 6460 17289 6469 17323
rect 6469 17289 6503 17323
rect 6503 17289 6512 17323
rect 6460 17280 6512 17289
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 7104 17280 7156 17332
rect 7840 17280 7892 17332
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 4160 17212 4212 17264
rect 5448 17212 5500 17264
rect 10140 17255 10192 17264
rect 10140 17221 10149 17255
rect 10149 17221 10183 17255
rect 10183 17221 10192 17255
rect 10140 17212 10192 17221
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 3240 17144 3292 17196
rect 2320 17051 2372 17060
rect 2320 17017 2329 17051
rect 2329 17017 2363 17051
rect 2363 17017 2372 17051
rect 2320 17008 2372 17017
rect 3700 17076 3752 17128
rect 6644 17144 6696 17196
rect 5264 17076 5316 17128
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 9588 17144 9640 17196
rect 10876 17280 10928 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 12808 17280 12860 17332
rect 13636 17280 13688 17332
rect 14648 17323 14700 17332
rect 14648 17289 14657 17323
rect 14657 17289 14691 17323
rect 14691 17289 14700 17323
rect 14648 17280 14700 17289
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 21732 17323 21784 17332
rect 17776 17280 17828 17289
rect 7564 17076 7616 17085
rect 9864 17076 9916 17128
rect 18144 17255 18196 17264
rect 18144 17221 18153 17255
rect 18153 17221 18187 17255
rect 18187 17221 18196 17255
rect 18144 17212 18196 17221
rect 21732 17289 21741 17323
rect 21741 17289 21775 17323
rect 21775 17289 21784 17323
rect 21732 17280 21784 17289
rect 4712 17051 4764 17060
rect 4712 17017 4721 17051
rect 4721 17017 4755 17051
rect 4755 17017 4764 17051
rect 4712 17008 4764 17017
rect 4896 17051 4948 17060
rect 4896 17017 4905 17051
rect 4905 17017 4939 17051
rect 4939 17017 4948 17051
rect 4896 17008 4948 17017
rect 6092 17051 6144 17060
rect 6092 17017 6101 17051
rect 6101 17017 6135 17051
rect 6135 17017 6144 17051
rect 6092 17008 6144 17017
rect 7472 17008 7524 17060
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 12532 17076 12584 17128
rect 13544 17076 13596 17128
rect 15752 17119 15804 17128
rect 15752 17085 15786 17119
rect 15786 17085 15804 17119
rect 15752 17076 15804 17085
rect 16764 17076 16816 17128
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 5080 16940 5132 16992
rect 8300 16940 8352 16992
rect 9772 16940 9824 16992
rect 12440 16940 12492 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 18604 16983 18656 16992
rect 18604 16949 18613 16983
rect 18613 16949 18647 16983
rect 18647 16949 18656 16983
rect 18604 16940 18656 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2412 16736 2464 16788
rect 6736 16736 6788 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 8208 16736 8260 16788
rect 9864 16736 9916 16788
rect 10968 16736 11020 16788
rect 3332 16668 3384 16720
rect 4712 16668 4764 16720
rect 8116 16668 8168 16720
rect 8484 16711 8536 16720
rect 8484 16677 8493 16711
rect 8493 16677 8527 16711
rect 8527 16677 8536 16711
rect 8484 16668 8536 16677
rect 2596 16600 2648 16652
rect 5080 16600 5132 16652
rect 5264 16643 5316 16652
rect 5264 16609 5298 16643
rect 5298 16609 5316 16643
rect 5264 16600 5316 16609
rect 8300 16600 8352 16652
rect 9680 16600 9732 16652
rect 10140 16668 10192 16720
rect 10784 16668 10836 16720
rect 11612 16736 11664 16788
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 17408 16736 17460 16788
rect 12440 16668 12492 16720
rect 12992 16668 13044 16720
rect 9956 16600 10008 16652
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 12164 16600 12216 16652
rect 16120 16600 16172 16652
rect 16580 16643 16632 16652
rect 16580 16609 16589 16643
rect 16589 16609 16623 16643
rect 16623 16609 16632 16643
rect 16580 16600 16632 16609
rect 16856 16643 16908 16652
rect 16856 16609 16890 16643
rect 16890 16609 16908 16643
rect 16856 16600 16908 16609
rect 4896 16532 4948 16584
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 2136 16396 2188 16448
rect 4620 16396 4672 16448
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2136 16192 2188 16244
rect 3148 16192 3200 16244
rect 8208 16192 8260 16244
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 8484 16192 8536 16244
rect 9588 16235 9640 16244
rect 9588 16201 9597 16235
rect 9597 16201 9631 16235
rect 9631 16201 9640 16235
rect 9588 16192 9640 16201
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 12992 16235 13044 16244
rect 12992 16201 13001 16235
rect 13001 16201 13035 16235
rect 13035 16201 13044 16235
rect 12992 16192 13044 16201
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 16580 16192 16632 16244
rect 5448 16124 5500 16176
rect 3884 16056 3936 16108
rect 4068 15988 4120 16040
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 11152 16056 11204 16108
rect 16856 16056 16908 16108
rect 1952 15920 2004 15972
rect 2964 15920 3016 15972
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 4160 15963 4212 15972
rect 4160 15929 4169 15963
rect 4169 15929 4203 15963
rect 4203 15929 4212 15963
rect 8668 15988 8720 16040
rect 4160 15920 4212 15929
rect 9588 15920 9640 15972
rect 13176 15920 13228 15972
rect 16488 15963 16540 15972
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7840 15895 7892 15904
rect 7840 15861 7849 15895
rect 7849 15861 7883 15895
rect 7883 15861 7892 15895
rect 7840 15852 7892 15861
rect 9680 15852 9732 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 16488 15929 16497 15963
rect 16497 15929 16531 15963
rect 16531 15929 16540 15963
rect 16488 15920 16540 15929
rect 15752 15852 15804 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 3332 15648 3384 15700
rect 5264 15648 5316 15700
rect 5632 15648 5684 15700
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 10048 15648 10100 15700
rect 12440 15648 12492 15700
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 16488 15648 16540 15700
rect 2504 15580 2556 15632
rect 5356 15580 5408 15632
rect 6000 15580 6052 15632
rect 6368 15580 6420 15632
rect 9496 15580 9548 15632
rect 10140 15580 10192 15632
rect 10784 15623 10836 15632
rect 10784 15589 10793 15623
rect 10793 15589 10827 15623
rect 10827 15589 10836 15623
rect 10784 15580 10836 15589
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 4160 15512 4212 15564
rect 4896 15512 4948 15564
rect 6460 15512 6512 15564
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 10324 15555 10376 15564
rect 9128 15512 9180 15521
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 2872 15444 2924 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 9864 15444 9916 15496
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 9680 15376 9732 15428
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 2504 15308 2556 15360
rect 2688 15308 2740 15360
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 5172 15308 5224 15360
rect 9588 15308 9640 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 4712 15104 4764 15156
rect 5264 15147 5316 15156
rect 5264 15113 5273 15147
rect 5273 15113 5307 15147
rect 5307 15113 5316 15147
rect 5264 15104 5316 15113
rect 5356 15104 5408 15156
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 6736 15036 6788 15088
rect 9772 15036 9824 15088
rect 1400 14968 1452 15020
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 6000 14968 6052 15020
rect 2872 14900 2924 14952
rect 5264 14832 5316 14884
rect 6092 14832 6144 14884
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 6460 14764 6512 14816
rect 7380 14832 7432 14884
rect 9864 14900 9916 14952
rect 10324 14900 10376 14952
rect 9680 14764 9732 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2596 14560 2648 14612
rect 2872 14560 2924 14612
rect 3516 14560 3568 14612
rect 4252 14560 4304 14612
rect 6000 14560 6052 14612
rect 9128 14603 9180 14612
rect 3884 14492 3936 14544
rect 4436 14535 4488 14544
rect 4436 14501 4445 14535
rect 4445 14501 4479 14535
rect 4479 14501 4488 14535
rect 4436 14492 4488 14501
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 1676 14467 1728 14476
rect 1676 14433 1710 14467
rect 1710 14433 1728 14467
rect 1676 14424 1728 14433
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 6000 14424 6052 14476
rect 4344 14356 4396 14408
rect 7380 14356 7432 14408
rect 5356 14288 5408 14340
rect 7656 14492 7708 14544
rect 7932 14492 7984 14544
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 14096 14492 14148 14544
rect 14280 14492 14332 14544
rect 9680 14424 9732 14476
rect 8208 14356 8260 14408
rect 9864 14356 9916 14408
rect 3424 14220 3476 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4436 14016 4488 14068
rect 1492 13991 1544 14000
rect 1492 13957 1501 13991
rect 1501 13957 1535 13991
rect 1535 13957 1544 13991
rect 1492 13948 1544 13957
rect 3056 13991 3108 14000
rect 3056 13957 3065 13991
rect 3065 13957 3099 13991
rect 3099 13957 3108 13991
rect 3056 13948 3108 13957
rect 3148 13948 3200 14000
rect 2596 13880 2648 13932
rect 3516 13880 3568 13932
rect 4896 13880 4948 13932
rect 6092 14016 6144 14068
rect 7380 14016 7432 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 7288 13948 7340 14000
rect 7656 13948 7708 14000
rect 9864 13948 9916 14000
rect 7564 13923 7616 13932
rect 7564 13889 7573 13923
rect 7573 13889 7607 13923
rect 7607 13889 7616 13923
rect 7564 13880 7616 13889
rect 4436 13812 4488 13864
rect 6000 13855 6052 13864
rect 1768 13787 1820 13796
rect 1768 13753 1777 13787
rect 1777 13753 1811 13787
rect 1811 13753 1820 13787
rect 1768 13744 1820 13753
rect 3056 13744 3108 13796
rect 3332 13787 3384 13796
rect 3332 13753 3341 13787
rect 3341 13753 3375 13787
rect 3375 13753 3384 13787
rect 3332 13744 3384 13753
rect 3608 13744 3660 13796
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 6460 13812 6512 13864
rect 8208 13812 8260 13864
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 8116 13744 8168 13796
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3240 13472 3292 13524
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 4344 13472 4396 13524
rect 6184 13472 6236 13524
rect 6736 13472 6788 13524
rect 8208 13472 8260 13524
rect 2136 13404 2188 13456
rect 4896 13447 4948 13456
rect 4896 13413 4930 13447
rect 4930 13413 4948 13447
rect 4896 13404 4948 13413
rect 7656 13447 7708 13456
rect 7656 13413 7665 13447
rect 7665 13413 7699 13447
rect 7699 13413 7708 13447
rect 7656 13404 7708 13413
rect 1860 13336 1912 13388
rect 7840 13336 7892 13388
rect 9772 13336 9824 13388
rect 10508 13336 10560 13388
rect 1676 13268 1728 13320
rect 3516 13268 3568 13320
rect 1768 13200 1820 13252
rect 2504 13200 2556 13252
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 6184 13268 6236 13320
rect 7196 13243 7248 13252
rect 7196 13209 7205 13243
rect 7205 13209 7239 13243
rect 7239 13209 7248 13243
rect 7196 13200 7248 13209
rect 4988 13132 5040 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 10048 13132 10100 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 4068 12928 4120 12980
rect 4896 12928 4948 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 10508 12928 10560 12980
rect 10968 12928 11020 12980
rect 9680 12903 9732 12912
rect 9680 12869 9689 12903
rect 9689 12869 9723 12903
rect 9723 12869 9732 12903
rect 9680 12860 9732 12869
rect 10692 12860 10744 12912
rect 3332 12792 3384 12844
rect 4620 12792 4672 12844
rect 11060 12792 11112 12844
rect 2872 12724 2924 12776
rect 4896 12724 4948 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 6000 12724 6052 12776
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 6460 12656 6512 12708
rect 8116 12724 8168 12776
rect 6736 12656 6788 12708
rect 11060 12656 11112 12708
rect 2872 12631 2924 12640
rect 2136 12588 2188 12597
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 2872 12588 2924 12597
rect 3240 12588 3292 12640
rect 4804 12588 4856 12640
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 11152 12588 11204 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 2596 12384 2648 12436
rect 2780 12384 2832 12436
rect 4068 12384 4120 12436
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 6736 12384 6788 12436
rect 7840 12384 7892 12436
rect 8852 12384 8904 12436
rect 9588 12384 9640 12436
rect 10968 12384 11020 12436
rect 4160 12316 4212 12368
rect 6184 12316 6236 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 4988 12248 5040 12300
rect 6552 12248 6604 12300
rect 8576 12248 8628 12300
rect 9588 12248 9640 12300
rect 11060 12248 11112 12300
rect 2044 12180 2096 12232
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 3608 12180 3660 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9772 12180 9824 12232
rect 8208 12112 8260 12164
rect 2688 12044 2740 12096
rect 3976 12044 4028 12096
rect 5264 12044 5316 12096
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 10048 12044 10100 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 2964 11840 3016 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 8484 11840 8536 11892
rect 4068 11772 4120 11824
rect 6000 11772 6052 11824
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 3240 11636 3292 11688
rect 4712 11636 4764 11688
rect 2596 11568 2648 11620
rect 5356 11611 5408 11620
rect 5356 11577 5365 11611
rect 5365 11577 5399 11611
rect 5399 11577 5408 11611
rect 5356 11568 5408 11577
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 5080 11500 5132 11552
rect 6552 11500 6604 11552
rect 7012 11500 7064 11552
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 7748 11500 7800 11552
rect 9588 11500 9640 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10140 11500 10192 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11296 1728 11348
rect 2872 11296 2924 11348
rect 3056 11296 3108 11348
rect 4804 11296 4856 11348
rect 6920 11296 6972 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 8576 11296 8628 11348
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 9772 11296 9824 11348
rect 4712 11228 4764 11280
rect 9680 11228 9732 11280
rect 1860 11160 1912 11212
rect 2136 11160 2188 11212
rect 2596 11203 2648 11212
rect 2596 11169 2605 11203
rect 2605 11169 2639 11203
rect 2639 11169 2648 11203
rect 2596 11160 2648 11169
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 5448 11160 5500 11212
rect 7748 11160 7800 11212
rect 11060 11160 11112 11212
rect 12716 11203 12768 11212
rect 12716 11169 12725 11203
rect 12725 11169 12759 11203
rect 12759 11169 12768 11203
rect 12716 11160 12768 11169
rect 4804 11092 4856 11144
rect 5356 11092 5408 11144
rect 6644 11092 6696 11144
rect 8300 11092 8352 11144
rect 10048 11092 10100 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 2228 11024 2280 11076
rect 2780 11024 2832 11076
rect 3608 11024 3660 11076
rect 4160 11067 4212 11076
rect 4160 11033 4169 11067
rect 4169 11033 4203 11067
rect 4203 11033 4212 11067
rect 4160 11024 4212 11033
rect 5448 11024 5500 11076
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 4712 10752 4764 10804
rect 6828 10752 6880 10804
rect 7748 10752 7800 10804
rect 11060 10752 11112 10804
rect 11612 10752 11664 10804
rect 12716 10752 12768 10804
rect 5264 10727 5316 10736
rect 5264 10693 5273 10727
rect 5273 10693 5307 10727
rect 5307 10693 5316 10727
rect 5264 10684 5316 10693
rect 8392 10727 8444 10736
rect 8392 10693 8401 10727
rect 8401 10693 8435 10727
rect 8435 10693 8444 10727
rect 8392 10684 8444 10693
rect 5448 10616 5500 10668
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 2412 10591 2464 10600
rect 2412 10557 2446 10591
rect 2446 10557 2464 10591
rect 2412 10548 2464 10557
rect 2780 10548 2832 10600
rect 3240 10480 3292 10532
rect 5448 10480 5500 10532
rect 6368 10548 6420 10600
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 6000 10480 6052 10532
rect 7932 10480 7984 10532
rect 1860 10412 1912 10464
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 4620 10412 4672 10464
rect 9680 10480 9732 10532
rect 9864 10480 9916 10532
rect 10232 10480 10284 10532
rect 12440 10523 12492 10532
rect 12440 10489 12449 10523
rect 12449 10489 12483 10523
rect 12483 10489 12492 10523
rect 12440 10480 12492 10489
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2412 10208 2464 10260
rect 2504 10208 2556 10260
rect 4068 10208 4120 10260
rect 4804 10208 4856 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7472 10208 7524 10260
rect 9680 10208 9732 10260
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 2688 10140 2740 10192
rect 3240 10140 3292 10192
rect 4988 10140 5040 10192
rect 8208 10140 8260 10192
rect 7288 10072 7340 10124
rect 7564 10072 7616 10124
rect 10876 10072 10928 10124
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 3516 10004 3568 10056
rect 4068 10004 4120 10056
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9864 10004 9916 10056
rect 2136 9868 2188 9920
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 7288 9868 7340 9920
rect 8392 9868 8444 9920
rect 9128 9868 9180 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 3148 9707 3200 9716
rect 3148 9673 3157 9707
rect 3157 9673 3191 9707
rect 3191 9673 3200 9707
rect 3148 9664 3200 9673
rect 5356 9664 5408 9716
rect 2320 9596 2372 9648
rect 2964 9596 3016 9648
rect 5540 9639 5592 9648
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 7748 9664 7800 9716
rect 14096 9664 14148 9716
rect 14280 9664 14332 9716
rect 7564 9596 7616 9648
rect 8576 9639 8628 9648
rect 8576 9605 8585 9639
rect 8585 9605 8619 9639
rect 8619 9605 8628 9639
rect 8576 9596 8628 9605
rect 11704 9596 11756 9648
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2412 9460 2464 9512
rect 3148 9460 3200 9512
rect 7196 9528 7248 9580
rect 8392 9528 8444 9580
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 3516 9503 3568 9512
rect 3516 9469 3550 9503
rect 3550 9469 3568 9503
rect 3516 9460 3568 9469
rect 7748 9460 7800 9512
rect 8208 9460 8260 9512
rect 2228 9435 2280 9444
rect 2228 9401 2237 9435
rect 2237 9401 2271 9435
rect 2271 9401 2280 9435
rect 2228 9392 2280 9401
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 7472 9435 7524 9444
rect 7472 9401 7481 9435
rect 7481 9401 7515 9435
rect 7515 9401 7524 9435
rect 7472 9392 7524 9401
rect 7840 9392 7892 9444
rect 9036 9435 9088 9444
rect 9036 9401 9045 9435
rect 9045 9401 9079 9435
rect 9079 9401 9088 9435
rect 9036 9392 9088 9401
rect 10692 9392 10744 9444
rect 11244 9392 11296 9444
rect 4896 9324 4948 9376
rect 7656 9324 7708 9376
rect 11796 9324 11848 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2044 9120 2096 9172
rect 2412 9120 2464 9172
rect 3516 9120 3568 9172
rect 7288 9120 7340 9172
rect 2228 9052 2280 9104
rect 7380 9052 7432 9104
rect 8392 9120 8444 9172
rect 9772 9120 9824 9172
rect 10692 9120 10744 9172
rect 10876 9120 10928 9172
rect 11704 9120 11756 9172
rect 7656 9095 7708 9104
rect 7656 9061 7665 9095
rect 7665 9061 7699 9095
rect 7699 9061 7708 9095
rect 7656 9052 7708 9061
rect 7932 9052 7984 9104
rect 11612 9052 11664 9104
rect 1492 8984 1544 9036
rect 1952 8984 2004 9036
rect 2320 8984 2372 9036
rect 3148 8984 3200 9036
rect 4712 8984 4764 9036
rect 4896 9027 4948 9036
rect 4896 8993 4930 9027
rect 4930 8993 4948 9027
rect 4896 8984 4948 8993
rect 7840 8984 7892 9036
rect 9956 8984 10008 9036
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 4804 8780 4856 8832
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 7012 8780 7064 8832
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 10140 8780 10192 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1768 8576 1820 8628
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 7656 8576 7708 8628
rect 8300 8576 8352 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 2780 8508 2832 8560
rect 5540 8508 5592 8560
rect 7932 8551 7984 8560
rect 7932 8517 7941 8551
rect 7941 8517 7975 8551
rect 7975 8517 7984 8551
rect 7932 8508 7984 8517
rect 10232 8576 10284 8628
rect 10876 8576 10928 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 11704 8508 11756 8560
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4896 8440 4948 8492
rect 1768 8372 1820 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 5080 8372 5132 8424
rect 6000 8372 6052 8424
rect 5540 8347 5592 8356
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 7196 8440 7248 8492
rect 7748 8372 7800 8424
rect 8024 8372 8076 8424
rect 9772 8372 9824 8424
rect 9128 8304 9180 8356
rect 9496 8304 9548 8356
rect 10968 8304 11020 8356
rect 2688 8279 2740 8288
rect 2688 8245 2697 8279
rect 2697 8245 2731 8279
rect 2731 8245 2740 8279
rect 2688 8236 2740 8245
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 3516 8236 3568 8288
rect 7748 8236 7800 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1492 8032 1544 8084
rect 2964 8032 3016 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 7196 8032 7248 8084
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 11612 8075 11664 8084
rect 11612 8041 11621 8075
rect 11621 8041 11655 8075
rect 11655 8041 11664 8075
rect 11612 8032 11664 8041
rect 3056 7964 3108 8016
rect 4712 7964 4764 8016
rect 7748 8007 7800 8016
rect 7748 7973 7757 8007
rect 7757 7973 7791 8007
rect 7791 7973 7800 8007
rect 7748 7964 7800 7973
rect 9956 8007 10008 8016
rect 9956 7973 9990 8007
rect 9990 7973 10008 8007
rect 9956 7964 10008 7973
rect 2504 7896 2556 7948
rect 2780 7896 2832 7948
rect 3792 7896 3844 7948
rect 5080 7896 5132 7948
rect 6644 7896 6696 7948
rect 8208 7896 8260 7948
rect 9772 7896 9824 7948
rect 10692 7896 10744 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 7380 7760 7432 7812
rect 8484 7692 8536 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2596 7488 2648 7540
rect 3240 7488 3292 7540
rect 3792 7531 3844 7540
rect 3792 7497 3801 7531
rect 3801 7497 3835 7531
rect 3835 7497 3844 7531
rect 3792 7488 3844 7497
rect 6644 7531 6696 7540
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7748 7488 7800 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 6920 7463 6972 7472
rect 6920 7429 6929 7463
rect 6929 7429 6963 7463
rect 6963 7429 6972 7463
rect 6920 7420 6972 7429
rect 4344 7284 4396 7336
rect 8484 7284 8536 7336
rect 9772 7284 9824 7336
rect 2320 7216 2372 7268
rect 7196 7259 7248 7268
rect 7196 7225 7205 7259
rect 7205 7225 7239 7259
rect 7239 7225 7248 7259
rect 7196 7216 7248 7225
rect 7380 7259 7432 7268
rect 7380 7225 7389 7259
rect 7389 7225 7423 7259
rect 7423 7225 7432 7259
rect 7380 7216 7432 7225
rect 5540 7148 5592 7200
rect 10692 7148 10744 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2504 6987 2556 6996
rect 2504 6953 2513 6987
rect 2513 6953 2547 6987
rect 2547 6953 2556 6987
rect 2504 6944 2556 6953
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5080 6987 5132 6996
rect 5080 6953 5089 6987
rect 5089 6953 5123 6987
rect 5123 6953 5132 6987
rect 5080 6944 5132 6953
rect 7196 6944 7248 6996
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 4252 6876 4304 6928
rect 2872 6808 2924 6860
rect 3792 6808 3844 6860
rect 4528 6808 4580 6860
rect 5448 6808 5500 6860
rect 2044 6740 2096 6792
rect 5540 6740 5592 6792
rect 5724 6808 5776 6860
rect 7840 6876 7892 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10140 6808 10192 6860
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 10968 6808 11020 6860
rect 6828 6740 6880 6792
rect 4528 6672 4580 6724
rect 5632 6672 5684 6724
rect 3976 6604 4028 6656
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 6092 6604 6144 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3700 6443 3752 6452
rect 3700 6409 3709 6443
rect 3709 6409 3743 6443
rect 3743 6409 3752 6443
rect 3700 6400 3752 6409
rect 4252 6400 4304 6452
rect 7840 6400 7892 6452
rect 2780 6375 2832 6384
rect 2780 6341 2789 6375
rect 2789 6341 2823 6375
rect 2823 6341 2832 6375
rect 2780 6332 2832 6341
rect 3148 6264 3200 6316
rect 4160 6264 4212 6316
rect 10048 6400 10100 6452
rect 10140 6400 10192 6452
rect 10324 6332 10376 6384
rect 1860 6196 1912 6248
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 4528 6239 4580 6248
rect 4528 6205 4562 6239
rect 4562 6205 4580 6239
rect 4528 6196 4580 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 1400 6060 1452 6112
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1860 5856 1912 5908
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 5540 5856 5592 5908
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 7196 5856 7248 5908
rect 7840 5856 7892 5908
rect 4712 5831 4764 5840
rect 4712 5797 4721 5831
rect 4721 5797 4755 5831
rect 4755 5797 4764 5831
rect 4712 5788 4764 5797
rect 2504 5720 2556 5772
rect 3976 5720 4028 5772
rect 4528 5720 4580 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 3240 5584 3292 5636
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 2044 5108 2096 5160
rect 2872 5108 2924 5160
rect 4160 5108 4212 5160
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 4620 4972 4672 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 4160 4768 4212 4820
rect 1952 4632 2004 4684
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 3240 4564 3292 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2044 4471 2096 4480
rect 2044 4437 2053 4471
rect 2053 4437 2087 4471
rect 2087 4437 2096 4471
rect 2044 4428 2096 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1952 4224 2004 4276
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 2504 4156 2556 4208
rect 2320 4020 2372 4072
rect 2688 3952 2740 4004
rect 2964 3995 3016 4004
rect 2964 3961 2973 3995
rect 2973 3961 3007 3995
rect 3007 3961 3016 3995
rect 2964 3952 3016 3961
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1492 3680 1544 3732
rect 2136 3680 2188 3732
rect 2228 3544 2280 3596
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 1492 2932 1544 2984
rect 3240 2932 3292 2984
rect 2504 2864 2556 2916
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 2780 2524 2832 2576
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2688 2295 2740 2304
rect 2688 2261 2697 2295
rect 2697 2261 2731 2295
rect 2731 2261 2740 2295
rect 2688 2252 2740 2261
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27520 3110 28000
rect 3330 27704 3386 27713
rect 3330 27639 3386 27648
rect 308 23769 336 27520
rect 860 24954 888 27520
rect 848 24948 900 24954
rect 848 24890 900 24896
rect 294 23760 350 23769
rect 294 23695 350 23704
rect 1412 23610 1440 27520
rect 1964 25514 1992 27520
rect 1964 25498 2084 25514
rect 1964 25492 2096 25498
rect 1964 25486 2044 25492
rect 2044 25434 2096 25440
rect 1584 25424 1636 25430
rect 1584 25366 1636 25372
rect 1596 24614 1624 25366
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1412 23582 1532 23610
rect 1504 22166 1532 23582
rect 1596 23497 1624 24550
rect 1780 24410 1808 25298
rect 2516 24698 2544 27520
rect 3068 26568 3096 27520
rect 2884 26540 3096 26568
rect 2688 25492 2740 25498
rect 2688 25434 2740 25440
rect 2700 24886 2728 25434
rect 2780 25220 2832 25226
rect 2780 25162 2832 25168
rect 2792 24954 2820 25162
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 2688 24880 2740 24886
rect 2688 24822 2740 24828
rect 2516 24670 2728 24698
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 1780 23730 1808 24346
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 24154 2544 24210
rect 2424 24138 2544 24154
rect 2412 24132 2544 24138
rect 2464 24126 2544 24132
rect 2412 24074 2464 24080
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1676 23520 1728 23526
rect 1582 23488 1638 23497
rect 1676 23462 1728 23468
rect 1582 23423 1638 23432
rect 1584 22976 1636 22982
rect 1688 22964 1716 23462
rect 1636 22936 1716 22964
rect 1584 22918 1636 22924
rect 1596 22438 1624 22918
rect 1674 22808 1730 22817
rect 1674 22743 1730 22752
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1492 22160 1544 22166
rect 1492 22102 1544 22108
rect 1596 22012 1624 22374
rect 1504 21984 1624 22012
rect 1504 21418 1532 21984
rect 1492 21412 1544 21418
rect 1492 21354 1544 21360
rect 1504 20942 1532 21354
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1504 19718 1532 20878
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1596 18902 1624 21286
rect 1688 20602 1716 22743
rect 2148 22234 2268 22250
rect 2136 22228 2268 22234
rect 2188 22222 2268 22228
rect 2136 22170 2188 22176
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1872 21078 1900 21830
rect 2148 21690 2176 22034
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 1860 21072 1912 21078
rect 1860 21014 1912 21020
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1688 20330 1716 20538
rect 2240 20398 2268 22222
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 2332 20058 2360 24006
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2424 22438 2452 23258
rect 2516 22642 2544 24126
rect 2608 23322 2636 24550
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2700 22681 2728 24670
rect 2780 24676 2832 24682
rect 2780 24618 2832 24624
rect 2792 24585 2820 24618
rect 2778 24576 2834 24585
rect 2778 24511 2834 24520
rect 2778 24440 2834 24449
rect 2778 24375 2834 24384
rect 2792 24206 2820 24375
rect 2884 24342 2912 26540
rect 2962 26480 3018 26489
rect 2962 26415 3018 26424
rect 2872 24336 2924 24342
rect 2872 24278 2924 24284
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2792 24070 2820 24142
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2884 23866 2912 24278
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2780 22976 2832 22982
rect 2976 22930 3004 26415
rect 3238 25256 3294 25265
rect 3056 25220 3108 25226
rect 3238 25191 3294 25200
rect 3056 25162 3108 25168
rect 3068 24682 3096 25162
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3056 24676 3108 24682
rect 3056 24618 3108 24624
rect 3068 24206 3096 24618
rect 3056 24200 3108 24206
rect 3056 24142 3108 24148
rect 3056 23248 3108 23254
rect 3056 23190 3108 23196
rect 2780 22918 2832 22924
rect 2792 22778 2820 22918
rect 2884 22902 3004 22930
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2686 22672 2742 22681
rect 2504 22636 2556 22642
rect 2686 22607 2742 22616
rect 2504 22578 2556 22584
rect 2792 22556 2820 22714
rect 2700 22528 2820 22556
rect 2596 22500 2648 22506
rect 2596 22442 2648 22448
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2608 22234 2636 22442
rect 2596 22228 2648 22234
rect 2596 22170 2648 22176
rect 2700 22030 2728 22528
rect 2688 22024 2740 22030
rect 2502 21992 2558 22001
rect 2884 22012 2912 22902
rect 3068 22642 3096 23190
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3160 22234 3188 25094
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 2884 21984 3096 22012
rect 2688 21966 2740 21972
rect 2502 21927 2504 21936
rect 2556 21927 2558 21936
rect 2596 21956 2648 21962
rect 2504 21898 2556 21904
rect 2596 21898 2648 21904
rect 2608 20602 2636 21898
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2884 21418 2912 21830
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2884 21146 2912 21354
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2884 20754 2912 21082
rect 2700 20726 2912 20754
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2700 20466 2728 20726
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19174 1900 19858
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 19378 1992 19654
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1860 19168 1912 19174
rect 1860 19110 1912 19116
rect 1584 18896 1636 18902
rect 1584 18838 1636 18844
rect 1872 18601 1900 19110
rect 1858 18592 1914 18601
rect 1858 18527 1914 18536
rect 1964 18358 1992 19314
rect 2516 18873 2544 19994
rect 2688 19984 2740 19990
rect 2688 19926 2740 19932
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 2608 18970 2636 19722
rect 2700 19310 2728 19926
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2688 18896 2740 18902
rect 2502 18864 2558 18873
rect 2044 18828 2096 18834
rect 2688 18838 2740 18844
rect 2502 18799 2558 18808
rect 2044 18770 2096 18776
rect 1952 18352 2004 18358
rect 1952 18294 2004 18300
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1872 17270 1900 18022
rect 1964 17814 1992 18294
rect 2056 18290 2084 18770
rect 2134 18728 2190 18737
rect 2134 18663 2136 18672
rect 2188 18663 2190 18672
rect 2136 18634 2188 18640
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2700 17898 2728 18838
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2700 17882 2820 17898
rect 2700 17876 2832 17882
rect 2700 17870 2780 17876
rect 2780 17818 2832 17824
rect 1952 17808 2004 17814
rect 1952 17750 2004 17756
rect 2318 17776 2374 17785
rect 2318 17711 2374 17720
rect 2412 17740 2464 17746
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1872 17105 1900 17206
rect 1858 17096 1914 17105
rect 2332 17066 2360 17711
rect 2412 17682 2464 17688
rect 2424 17202 2452 17682
rect 2884 17610 2912 18770
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2976 17814 3004 18158
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 1858 17031 1914 17040
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 2424 16794 2452 17138
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2148 16250 2176 16390
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14482 1440 14962
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1492 14000 1544 14006
rect 1492 13942 1544 13948
rect 1504 9042 1532 13942
rect 1688 13326 1716 14418
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 11898 1716 13262
rect 1780 13258 1808 13738
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1872 12442 1900 13330
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1688 10810 1716 11290
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1872 10470 1900 11154
rect 1860 10464 1912 10470
rect 1766 10432 1822 10441
rect 1860 10406 1912 10412
rect 1766 10367 1822 10376
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8090 1532 8978
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1596 7585 1624 8502
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1688 7449 1716 8910
rect 1780 8634 1808 10367
rect 1872 8922 1900 10406
rect 1964 9042 1992 15914
rect 2148 15026 2176 16186
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2516 15366 2544 15574
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2148 12646 2176 13398
rect 2240 13297 2268 15302
rect 2608 14618 2636 16594
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15745 3004 15914
rect 2962 15736 3018 15745
rect 2962 15671 3018 15680
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 2700 15502 2728 15535
rect 2688 15496 2740 15502
rect 2872 15496 2924 15502
rect 2688 15438 2740 15444
rect 2870 15464 2872 15473
rect 2924 15464 2926 15473
rect 2870 15399 2926 15408
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 15201 2728 15302
rect 2686 15192 2742 15201
rect 2686 15127 2742 15136
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 13938 2636 14554
rect 2700 14226 2728 15127
rect 2884 14958 2912 15399
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14618 2912 14894
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 3068 14226 3096 21984
rect 3148 21956 3200 21962
rect 3148 21898 3200 21904
rect 3160 19786 3188 21898
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 3146 18864 3202 18873
rect 3252 18834 3280 25191
rect 3146 18799 3202 18808
rect 3240 18828 3292 18834
rect 3160 18630 3188 18799
rect 3240 18770 3292 18776
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3160 18329 3188 18566
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3160 17338 3188 18158
rect 3252 18154 3280 18566
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3160 16250 3188 17274
rect 3252 17202 3280 18090
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3344 16726 3372 27639
rect 3606 27520 3662 28000
rect 4158 27520 4214 28000
rect 4710 27520 4766 28000
rect 5262 27520 5318 28000
rect 5814 27520 5870 28000
rect 6366 27520 6422 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8114 27520 8170 28000
rect 8666 27520 8722 28000
rect 9218 27520 9274 28000
rect 9770 27520 9826 28000
rect 10322 27520 10378 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 15934 27520 15990 28000
rect 16486 27520 16542 28000
rect 17038 27520 17094 28000
rect 17590 27520 17646 28000
rect 18142 27520 18198 28000
rect 18694 27520 18750 28000
rect 19246 27520 19302 28000
rect 19798 27520 19854 28000
rect 20350 27520 20406 28000
rect 20902 27520 20958 28000
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3620 26058 3648 27520
rect 4066 27160 4122 27169
rect 4066 27095 4122 27104
rect 4080 26586 4108 27095
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 3620 26030 3832 26058
rect 3698 25936 3754 25945
rect 3698 25871 3754 25880
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3436 24818 3464 25230
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3436 24290 3464 24754
rect 3436 24262 3556 24290
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3436 24070 3464 24142
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3436 23594 3464 24006
rect 3528 23866 3556 24262
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3424 23588 3476 23594
rect 3424 23530 3476 23536
rect 3436 22982 3464 23530
rect 3528 23254 3556 23802
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3606 23080 3662 23089
rect 3606 23015 3662 23024
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3620 22778 3648 23015
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3514 20224 3570 20233
rect 3514 20159 3570 20168
rect 3528 20058 3556 20159
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3712 17134 3740 25871
rect 3804 23361 3832 26030
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 3896 24614 3924 24890
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3790 23352 3846 23361
rect 3790 23287 3846 23296
rect 3896 22506 3924 24550
rect 4172 24449 4200 27520
rect 4158 24440 4214 24449
rect 4158 24375 4214 24384
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4160 24064 4212 24070
rect 4066 24032 4122 24041
rect 4160 24006 4212 24012
rect 4066 23967 4122 23976
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3988 23186 4016 23598
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3988 22778 4016 23122
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 4080 22681 4108 23967
rect 4066 22672 4122 22681
rect 4066 22607 4122 22616
rect 3884 22500 3936 22506
rect 3884 22442 3936 22448
rect 4068 22500 4120 22506
rect 4172 22488 4200 24006
rect 4120 22460 4200 22488
rect 4068 22442 4120 22448
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3804 20330 3832 21626
rect 3882 21584 3938 21593
rect 3882 21519 3938 21528
rect 3792 20324 3844 20330
rect 3792 20266 3844 20272
rect 3804 20058 3832 20266
rect 3896 20097 3924 21519
rect 3988 20856 4016 22170
rect 4264 22030 4292 24142
rect 4434 23760 4490 23769
rect 4434 23695 4490 23704
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4448 21894 4476 23695
rect 4526 22264 4582 22273
rect 4526 22199 4582 22208
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4540 21690 4568 22199
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4632 21622 4660 21966
rect 4724 21876 4752 27520
rect 5170 23216 5226 23225
rect 5080 23180 5132 23186
rect 5170 23151 5226 23160
rect 5080 23122 5132 23128
rect 5092 22642 5120 23122
rect 5184 22778 5212 23151
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 5092 22234 5120 22578
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 5276 22148 5304 27520
rect 5828 25242 5856 27520
rect 5828 25214 6040 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24818 6040 25214
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 6092 24744 6144 24750
rect 6092 24686 6144 24692
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5368 23730 5396 24006
rect 5448 23792 5500 23798
rect 5448 23734 5500 23740
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5184 22120 5304 22148
rect 5184 22012 5212 22120
rect 4908 21984 5212 22012
rect 4724 21848 4844 21876
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4528 21072 4580 21078
rect 4528 21014 4580 21020
rect 4160 20868 4212 20874
rect 3988 20828 4160 20856
rect 4160 20810 4212 20816
rect 4252 20528 4304 20534
rect 4066 20496 4122 20505
rect 4540 20482 4568 21014
rect 4304 20476 4568 20482
rect 4252 20470 4568 20476
rect 4264 20454 4568 20470
rect 4066 20431 4122 20440
rect 3882 20088 3938 20097
rect 3792 20052 3844 20058
rect 3882 20023 3938 20032
rect 3792 19994 3844 20000
rect 4080 19825 4108 20431
rect 4540 19990 4568 20454
rect 4528 19984 4580 19990
rect 4528 19926 4580 19932
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4540 19446 4568 19926
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3804 18766 3832 19110
rect 4172 18986 4200 19110
rect 4080 18958 4200 18986
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3804 18630 3832 18702
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3804 18154 3832 18566
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 4080 17921 4108 18958
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4632 18426 4660 18838
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 4066 17912 4122 17921
rect 4172 17882 4200 18090
rect 4066 17847 4122 17856
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3974 16960 4030 16969
rect 3332 16720 3384 16726
rect 3252 16680 3332 16708
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 2700 14198 2820 14226
rect 3068 14198 3188 14226
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2410 13424 2466 13433
rect 2410 13359 2466 13368
rect 2226 13288 2282 13297
rect 2226 13223 2282 13232
rect 2424 12986 2452 13359
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 9518 2084 12174
rect 2148 11218 2176 12582
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 9178 2084 9454
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1872 8894 1992 8922
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1780 8430 1808 8570
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1674 7440 1730 7449
rect 1674 7375 1730 7384
rect 1872 6254 1900 7822
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 2689 1440 6054
rect 1872 5914 1900 6190
rect 1964 5953 1992 8894
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 6254 2084 6734
rect 2044 6248 2096 6254
rect 2042 6216 2044 6225
rect 2096 6216 2098 6225
rect 2042 6151 2098 6160
rect 1950 5944 2006 5953
rect 1860 5908 1912 5914
rect 1950 5879 2006 5888
rect 1860 5850 1912 5856
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 4690 1992 5646
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 3913 1624 4422
rect 1964 4282 1992 4626
rect 2056 4486 2084 5102
rect 2044 4480 2096 4486
rect 2042 4448 2044 4457
rect 2096 4448 2098 4457
rect 2042 4383 2098 4392
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1582 3904 1638 3913
rect 1582 3839 1638 3848
rect 2148 3738 2176 9862
rect 2240 9450 2268 11018
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10266 2452 10542
rect 2516 10266 2544 13194
rect 2608 12442 2636 13874
rect 2792 12442 2820 14198
rect 3160 14006 3188 14198
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3068 13802 3096 13942
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12782 2912 13126
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2608 11218 2636 11562
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 9654 2360 9998
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2424 9518 2452 10202
rect 2700 10198 2728 12038
rect 2884 11354 2912 12582
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11898 3004 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3068 11354 3096 13738
rect 3252 13530 3280 16680
rect 3332 16662 3384 16668
rect 3896 16114 3924 16934
rect 3974 16895 4030 16904
rect 3988 16153 4016 16895
rect 3974 16144 4030 16153
rect 3884 16108 3936 16114
rect 4172 16130 4200 17206
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4724 16726 4752 17002
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 3974 16079 4030 16088
rect 4080 16102 4200 16130
rect 3884 16050 3936 16056
rect 4080 16046 4108 16102
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3344 15706 3372 15914
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 4172 15570 4200 15914
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4632 15502 4660 16390
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14618 3556 14758
rect 3606 14648 3662 14657
rect 3516 14612 3568 14618
rect 3606 14583 3662 14592
rect 3516 14554 3568 14560
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3252 12646 3280 13466
rect 3344 12850 3372 13738
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10606 2820 11018
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 3252 10538 3280 11630
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3252 10198 3280 10474
rect 2688 10192 2740 10198
rect 2594 10160 2650 10169
rect 3240 10192 3292 10198
rect 3160 10152 3240 10180
rect 2740 10140 3096 10146
rect 2688 10134 3096 10140
rect 2700 10118 3096 10134
rect 2594 10095 2650 10104
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 9110 2268 9386
rect 2424 9178 2452 9454
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8634 2360 8978
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 4078 2360 7210
rect 2516 7002 2544 7890
rect 2608 7546 2636 10095
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2700 6361 2728 8230
rect 2792 7954 2820 8502
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2884 7041 2912 8774
rect 2976 8090 3004 9590
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3068 8022 3096 10118
rect 3160 9722 3188 10152
rect 3240 10134 3292 10140
rect 3436 10044 3464 14214
rect 3528 13938 3556 14554
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3528 13530 3556 13874
rect 3620 13802 3648 14583
rect 3896 14550 3924 15302
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 3884 14544 3936 14550
rect 3884 14486 3936 14492
rect 3988 14385 4016 14991
rect 4632 14793 4660 15438
rect 4724 15162 4752 15438
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4618 14784 4674 14793
rect 4618 14719 4674 14728
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3974 14376 4030 14385
rect 3974 14311 4030 14320
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3528 13326 3556 13466
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 4068 12980 4120 12986
rect 4264 12968 4292 14554
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 13530 4384 14350
rect 4448 14074 4476 14486
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4120 12940 4292 12968
rect 4068 12922 4120 12928
rect 4080 12442 4108 12922
rect 4448 12617 4476 13806
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4434 12608 4490 12617
rect 4434 12543 4490 12552
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4160 12368 4212 12374
rect 4066 12336 4122 12345
rect 4160 12310 4212 12316
rect 4066 12271 4068 12280
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 11558 3648 12174
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11082 3648 11494
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10062 3556 10406
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3252 10016 3464 10044
rect 3516 10056 3568 10062
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3160 9518 3188 9658
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 9042 3188 9454
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3160 7410 3188 8230
rect 3252 7546 3280 10016
rect 3804 10033 3832 10231
rect 3516 9998 3568 10004
rect 3790 10024 3846 10033
rect 3528 9518 3556 9998
rect 3790 9959 3846 9968
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3896 8809 3924 11319
rect 3988 9489 4016 12038
rect 4080 11830 4108 12242
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4172 11098 4200 12310
rect 4632 11150 4660 12786
rect 4816 12646 4844 21848
rect 4908 18034 4936 21984
rect 5368 21962 5396 23462
rect 5460 22556 5488 23734
rect 5552 23662 5580 24550
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 6000 23316 6052 23322
rect 6000 23258 6052 23264
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5722 22672 5778 22681
rect 5722 22607 5778 22616
rect 5540 22568 5592 22574
rect 5460 22528 5540 22556
rect 5460 22098 5488 22528
rect 5540 22510 5592 22516
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5000 21690 5028 21830
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 5000 21146 5028 21626
rect 5184 21486 5212 21830
rect 5448 21616 5500 21622
rect 5446 21584 5448 21593
rect 5500 21584 5502 21593
rect 5446 21519 5502 21528
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5276 21146 5304 21354
rect 5552 21185 5580 22102
rect 5736 22030 5764 22607
rect 6012 22438 6040 23258
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6104 22114 6132 24686
rect 6184 24336 6236 24342
rect 6184 24278 6236 24284
rect 6196 23594 6224 24278
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6184 23588 6236 23594
rect 6184 23530 6236 23536
rect 6196 23118 6224 23530
rect 6288 23254 6316 23666
rect 6276 23248 6328 23254
rect 6276 23190 6328 23196
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6196 22778 6224 23054
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6274 22536 6330 22545
rect 6274 22471 6276 22480
rect 6328 22471 6330 22480
rect 6276 22442 6328 22448
rect 6380 22386 6408 27520
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6095 22086 6132 22114
rect 6288 22358 6408 22386
rect 6095 22080 6123 22086
rect 6012 22052 6123 22080
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5538 21176 5594 21185
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 5264 21140 5316 21146
rect 5538 21111 5540 21120
rect 5264 21082 5316 21088
rect 5592 21111 5594 21120
rect 5540 21082 5592 21088
rect 5000 20602 5028 21082
rect 5736 21078 5764 21422
rect 6012 21418 6040 22052
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6104 21690 6132 21898
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5736 20856 5764 21014
rect 5552 20828 5764 20856
rect 5552 20602 5580 20828
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5000 19990 5028 20538
rect 5552 19990 5580 20538
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5000 19514 5028 19926
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5092 19378 5120 19654
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 5000 18170 5028 18770
rect 5092 18290 5120 19314
rect 5184 19242 5212 19790
rect 5460 19310 5488 19858
rect 5814 19816 5870 19825
rect 5814 19751 5816 19760
rect 5868 19751 5870 19760
rect 5816 19722 5868 19728
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 5000 18142 5120 18170
rect 5092 18086 5120 18142
rect 5080 18080 5132 18086
rect 4908 18006 5028 18034
rect 5080 18022 5132 18028
rect 4894 17912 4950 17921
rect 4894 17847 4950 17856
rect 4908 17066 4936 17847
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4908 15570 4936 16526
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 5000 13977 5028 18006
rect 5092 17678 5120 18022
rect 5276 17882 5304 18362
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5552 17814 5580 18906
rect 6012 18630 6040 19178
rect 6182 19136 6238 19145
rect 6182 19071 6238 19080
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18566
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6196 18193 6224 19071
rect 6182 18184 6238 18193
rect 6182 18119 6238 18128
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 17338 5120 17614
rect 5262 17368 5318 17377
rect 5080 17332 5132 17338
rect 5262 17303 5318 17312
rect 5080 17274 5132 17280
rect 5092 16998 5120 17274
rect 5276 17134 5304 17303
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16658 5120 16934
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5276 15706 5304 16594
rect 5368 15722 5396 17750
rect 5552 17338 5580 17750
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5460 16182 5488 17206
rect 6090 17096 6146 17105
rect 6090 17031 6092 17040
rect 6144 17031 6146 17040
rect 6092 17002 6144 17008
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5264 15700 5316 15706
rect 5368 15694 5488 15722
rect 5644 15706 5672 15846
rect 5264 15642 5316 15648
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4986 13968 5042 13977
rect 4896 13932 4948 13938
rect 4986 13903 5042 13912
rect 4896 13874 4948 13880
rect 4908 13462 4936 13874
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4908 12986 4936 13398
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4908 12782 4936 12922
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5000 12646 5028 13126
rect 4804 12640 4856 12646
rect 4710 12608 4766 12617
rect 4804 12582 4856 12588
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4710 12543 4766 12552
rect 4724 12442 4752 12543
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4724 11694 4752 12378
rect 5000 12306 5028 12582
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4816 11354 4844 11834
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4712 11280 4764 11286
rect 4710 11248 4712 11257
rect 4764 11248 4766 11257
rect 4710 11183 4766 11192
rect 4080 11082 4200 11098
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4080 11076 4212 11082
rect 4080 11070 4160 11076
rect 4080 10266 4108 11070
rect 4160 11018 4212 11024
rect 4632 10470 4660 11086
rect 4724 10810 4752 11183
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3882 8800 3938 8809
rect 3882 8735 3938 8744
rect 4080 8498 4108 9998
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3882 8392 3938 8401
rect 4080 8378 4108 8434
rect 3882 8327 3938 8336
rect 3988 8350 4108 8378
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2870 7032 2926 7041
rect 3528 7002 3556 8230
rect 3896 8090 3924 8327
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3804 7546 3832 7890
rect 3792 7540 3844 7546
rect 3712 7500 3792 7528
rect 2870 6967 2926 6976
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2780 6384 2832 6390
rect 2686 6352 2742 6361
rect 2780 6326 2832 6332
rect 2686 6287 2742 6296
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2516 5681 2544 5714
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2516 5370 2544 5607
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2792 5250 2820 6326
rect 2516 5222 2820 5250
rect 2516 4690 2544 5222
rect 2884 5166 2912 6802
rect 3712 6458 3740 7500
rect 3792 7482 3844 7488
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3054 5944 3110 5953
rect 3160 5914 3188 6258
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3054 5879 3110 5888
rect 3148 5908 3200 5914
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2516 4214 2544 4626
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2962 4040 3018 4049
rect 2688 4004 2740 4010
rect 2962 3975 2964 3984
rect 2688 3946 2740 3952
rect 3016 3975 3018 3984
rect 2964 3946 3016 3952
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 1504 2990 1532 3674
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1952 3528 2004 3534
rect 2240 3505 2268 3538
rect 1952 3470 2004 3476
rect 2226 3496 2282 3505
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1398 2680 1454 2689
rect 1964 2650 1992 3470
rect 2226 3431 2282 3440
rect 2240 3194 2268 3431
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 1398 2615 1454 2624
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2516 2514 2544 2858
rect 2700 2666 2728 3946
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 3194 2912 3295
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2700 2638 2820 2666
rect 2792 2582 2820 2638
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 1596 1465 1624 2246
rect 2700 2145 2728 2246
rect 2686 2136 2742 2145
rect 2686 2071 2742 2080
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 3068 377 3096 5879
rect 3148 5850 3200 5856
rect 3252 5642 3280 6054
rect 3804 5914 3832 6802
rect 3988 6662 4016 8350
rect 4264 8090 4292 8366
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4264 7426 4292 8026
rect 4264 7398 4384 7426
rect 4356 7342 4384 7398
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6322 4200 6598
rect 4264 6458 4292 6870
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4540 6730 4568 6802
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4264 5953 4292 6394
rect 4540 6254 4568 6666
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4250 5944 4306 5953
rect 3792 5908 3844 5914
rect 4250 5879 4306 5888
rect 3792 5850 3844 5856
rect 3606 5808 3662 5817
rect 4540 5778 4568 6190
rect 3606 5743 3662 5752
rect 3976 5772 4028 5778
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3160 4593 3188 4966
rect 3240 4616 3292 4622
rect 3146 4584 3202 4593
rect 3240 4558 3292 4564
rect 3146 4519 3202 4528
rect 3252 3194 3280 4558
rect 3620 4282 3648 5743
rect 3976 5714 4028 5720
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 3988 5370 4016 5714
rect 4632 5710 4660 10406
rect 4816 10266 4844 11086
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 5000 10198 5028 12242
rect 5092 11558 5120 13670
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4724 8634 4752 8978
rect 4816 8838 4844 9862
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 9042 4936 9318
rect 5092 9081 5120 11494
rect 5078 9072 5134 9081
rect 4896 9036 4948 9042
rect 5078 9007 5134 9016
rect 4896 8978 4948 8984
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4724 8022 4752 8570
rect 4908 8498 4936 8978
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 5092 7954 5120 8366
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5092 7002 5120 7890
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4712 5840 4764 5846
rect 4710 5808 4712 5817
rect 4764 5808 4766 5817
rect 4710 5743 4766 5752
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4250 5128 4306 5137
rect 4172 4826 4200 5102
rect 4250 5063 4306 5072
rect 4264 5030 4292 5063
rect 4632 5030 4660 5646
rect 4724 5370 4752 5743
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3252 2990 3280 3130
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4264 921 4292 2246
rect 4250 912 4306 921
rect 4250 847 4306 856
rect 4632 480 4660 4966
rect 5184 4049 5212 15302
rect 5262 15192 5318 15201
rect 5368 15162 5396 15574
rect 5262 15127 5264 15136
rect 5316 15127 5318 15136
rect 5356 15156 5408 15162
rect 5264 15098 5316 15104
rect 5356 15098 5408 15104
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14521 5304 14826
rect 5262 14512 5318 14521
rect 5262 14447 5264 14456
rect 5316 14447 5318 14456
rect 5264 14418 5316 14424
rect 5368 14346 5396 15098
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5460 13376 5488 15694
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15026 6040 15574
rect 6090 15192 6146 15201
rect 6090 15127 6146 15136
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6012 14618 6040 14962
rect 6104 14890 6132 15127
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 13870 6040 14418
rect 6090 14104 6146 14113
rect 6090 14039 6092 14048
rect 6144 14039 6146 14048
rect 6092 14010 6144 14016
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5368 13348 5488 13376
rect 5368 12186 5396 13348
rect 6012 13297 6040 13806
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6196 13326 6224 13466
rect 6184 13320 6236 13326
rect 5446 13288 5502 13297
rect 5446 13223 5502 13232
rect 5998 13288 6054 13297
rect 6184 13262 6236 13268
rect 5998 13223 6054 13232
rect 5460 12782 5488 13223
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6196 12986 6224 13262
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5368 12158 5488 12186
rect 5264 12096 5316 12102
rect 5316 12056 5396 12084
rect 5264 12038 5316 12044
rect 5368 11626 5396 12056
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 11529 5396 11562
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5368 11150 5396 11455
rect 5460 11218 5488 12158
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11830 6040 12718
rect 6196 12374 6224 12922
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6196 11898 6224 12310
rect 6288 11937 6316 22358
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6380 19514 6408 19790
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6380 18970 6408 19450
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6472 17338 6500 17682
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15638 6408 16390
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 14822 6500 15506
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6366 14512 6422 14521
rect 6366 14447 6422 14456
rect 6274 11928 6330 11937
rect 6184 11892 6236 11898
rect 6274 11863 6330 11872
rect 6184 11834 6236 11840
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5814 11384 5870 11393
rect 5814 11319 5870 11328
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5828 11082 5856 11319
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5276 10033 5304 10678
rect 5460 10674 5488 11018
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 10577 5764 10610
rect 6380 10606 6408 14447
rect 6472 13870 6500 14758
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6564 12889 6592 24754
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 6656 23526 6684 24210
rect 6932 24138 6960 27520
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 7194 23760 7250 23769
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6656 22098 6684 23462
rect 6840 23322 6868 23734
rect 7194 23695 7250 23704
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21554 6776 21830
rect 6840 21690 6868 22170
rect 6932 21962 6960 23462
rect 7102 23352 7158 23361
rect 7102 23287 7158 23296
rect 7116 22710 7144 23287
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7116 22574 7144 22646
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7208 22166 7236 23695
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 7208 21690 7236 22102
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6932 21457 6960 21558
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6918 21448 6974 21457
rect 6918 21383 6974 21392
rect 7116 21146 7144 21490
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 20330 6684 20742
rect 7116 20398 7144 21082
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6656 18222 6684 20266
rect 7116 20058 7144 20334
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7208 18834 7236 19178
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 6918 18728 6974 18737
rect 6918 18663 6920 18672
rect 6972 18663 6974 18672
rect 6920 18634 6972 18640
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6748 18154 6776 18566
rect 7208 18426 7236 18770
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6748 17882 6776 18090
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6748 17746 6776 17818
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6550 12880 6606 12889
rect 6550 12815 6606 12824
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6368 10600 6420 10606
rect 5722 10568 5778 10577
rect 5448 10532 5500 10538
rect 6368 10542 6420 10548
rect 5722 10503 5778 10512
rect 6000 10532 6052 10538
rect 5448 10474 5500 10480
rect 6000 10474 6052 10480
rect 5460 10266 5488 10474
rect 5448 10260 5500 10266
rect 5368 10220 5448 10248
rect 5262 10024 5318 10033
rect 5262 9959 5318 9968
rect 5368 9722 5396 10220
rect 5448 10202 5500 10208
rect 5448 10056 5500 10062
rect 5500 10016 5580 10044
rect 5448 9998 5500 10004
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5552 9654 5580 10016
rect 6012 9926 6040 10474
rect 6472 10441 6500 12650
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12306 6592 12582
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 11558 6592 12242
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6656 11150 6684 17138
rect 6748 16794 6776 17682
rect 7024 17338 7052 17750
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15609 6868 15846
rect 6826 15600 6882 15609
rect 6826 15535 6882 15544
rect 7010 15464 7066 15473
rect 7010 15399 7012 15408
rect 7064 15399 7066 15408
rect 7012 15370 7064 15376
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6748 13530 6776 15030
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6748 12714 6776 13466
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6748 12442 6776 12650
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 7116 12345 7144 17274
rect 7300 15008 7328 26522
rect 7576 24410 7604 27520
rect 8128 24834 8156 27520
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 7852 24806 8156 24834
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7392 22778 7420 23666
rect 7654 23624 7710 23633
rect 7654 23559 7710 23568
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7472 22568 7524 22574
rect 7378 22536 7434 22545
rect 7472 22510 7524 22516
rect 7378 22471 7380 22480
rect 7432 22471 7434 22480
rect 7380 22442 7432 22448
rect 7484 22098 7512 22510
rect 7668 22234 7696 23559
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21593 7420 21830
rect 7378 21584 7434 21593
rect 7378 21519 7434 21528
rect 7392 21418 7420 21519
rect 7576 21486 7604 22034
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7576 21146 7604 21422
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7668 20058 7696 21626
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7484 18086 7512 18702
rect 7668 18630 7696 19994
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 17882 7512 18022
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17134 7420 17614
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7484 17066 7512 17818
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7576 16794 7604 17070
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7300 14980 7696 15008
rect 7562 14920 7618 14929
rect 7380 14884 7432 14890
rect 7562 14855 7618 14864
rect 7380 14826 7432 14832
rect 7194 14784 7250 14793
rect 7194 14719 7250 14728
rect 7208 13258 7236 14719
rect 7392 14414 7420 14826
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 14278 7420 14350
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 14074 7420 14214
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7102 12336 7158 12345
rect 7102 12271 7158 12280
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6828 10804 6880 10810
rect 6932 10792 6960 11290
rect 7024 11014 7052 11494
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6880 10764 6960 10792
rect 6828 10746 6880 10752
rect 7024 10606 7052 10950
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6458 10432 6514 10441
rect 6458 10367 6514 10376
rect 7300 10130 7328 13942
rect 7576 13938 7604 14855
rect 7668 14550 7696 14980
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7668 14006 7696 14486
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7656 13456 7708 13462
rect 7654 13424 7656 13433
rect 7708 13424 7710 13433
rect 7654 13359 7710 13368
rect 7760 11801 7788 24074
rect 7852 17338 7880 24806
rect 8116 24744 8168 24750
rect 8114 24712 8116 24721
rect 8220 24732 8248 25366
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 8168 24712 8248 24732
rect 8170 24704 8248 24712
rect 8312 24682 8340 25298
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8114 24647 8170 24656
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8588 24410 8616 25230
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 7932 22976 7984 22982
rect 7932 22918 7984 22924
rect 7944 22642 7972 22918
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7930 20088 7986 20097
rect 7930 20023 7986 20032
rect 7944 19854 7972 20023
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7944 19514 7972 19790
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7944 17610 7972 18838
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 13394 7880 15846
rect 7930 14920 7986 14929
rect 7930 14855 7986 14864
rect 7944 14550 7972 14855
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 12442 7880 13330
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7930 12336 7986 12345
rect 7930 12271 7986 12280
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7746 11792 7802 11801
rect 7746 11727 7802 11736
rect 7748 11552 7800 11558
rect 7852 11540 7880 12038
rect 7800 11512 7880 11540
rect 7748 11494 7800 11500
rect 7760 11218 7788 11494
rect 7944 11354 7972 12271
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10266 7512 10950
rect 7760 10810 7788 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7378 10024 7434 10033
rect 7378 9959 7434 9968
rect 6000 9920 6052 9926
rect 5998 9888 6000 9897
rect 7288 9920 7340 9926
rect 6052 9888 6054 9897
rect 5622 9820 5918 9840
rect 7288 9862 7340 9868
rect 5998 9823 6054 9832
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 8401 5580 8502
rect 6012 8430 6040 8774
rect 6000 8424 6052 8430
rect 5538 8392 5594 8401
rect 5538 8327 5540 8336
rect 5592 8327 5594 8336
rect 5722 8392 5778 8401
rect 6000 8366 6052 8372
rect 6090 8392 6146 8401
rect 5722 8327 5724 8336
rect 5540 8298 5592 8304
rect 5776 8327 5778 8336
rect 6090 8327 6146 8336
rect 5724 8298 5776 8304
rect 5538 8256 5594 8265
rect 5538 8191 5594 8200
rect 5552 7528 5580 8191
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5552 7500 5672 7528
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6882 5580 7142
rect 5460 6866 5580 6882
rect 5448 6860 5580 6866
rect 5500 6854 5580 6860
rect 5448 6802 5500 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 5914 5580 6734
rect 5644 6730 5672 7500
rect 5722 7440 5778 7449
rect 5722 7375 5778 7384
rect 5736 6866 5764 7375
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 6104 6662 6132 8327
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7546 6684 7890
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6840 6254 6868 6734
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5914 6868 6190
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6932 5681 6960 7414
rect 6918 5672 6974 5681
rect 6918 5607 6974 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 7024 3505 7052 8774
rect 7208 8498 7236 9522
rect 7300 9450 7328 9862
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 9178 7328 9386
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7392 9110 7420 9959
rect 7484 9450 7512 10202
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9654 7604 10066
rect 7760 10062 7788 10746
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9722 7788 9998
rect 7838 9888 7894 9897
rect 7838 9823 7894 9832
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9110 7696 9318
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7668 8634 7696 9046
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 8090 7236 8434
rect 7760 8430 7788 9454
rect 7852 9450 7880 9823
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7852 9042 7880 9386
rect 7944 9110 7972 10474
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7944 8566 7972 9046
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 8036 8430 8064 24346
rect 8680 23474 8708 27520
rect 9232 24834 9260 27520
rect 9404 25220 9456 25226
rect 9404 25162 9456 25168
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 8404 23446 8708 23474
rect 8772 24806 9260 24834
rect 8208 22704 8260 22710
rect 8206 22672 8208 22681
rect 8260 22672 8262 22681
rect 8206 22607 8262 22616
rect 8300 20800 8352 20806
rect 8220 20748 8300 20754
rect 8220 20742 8352 20748
rect 8220 20726 8340 20742
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 19854 8156 20198
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8128 19446 8156 19790
rect 8220 19786 8248 20726
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 8128 19224 8156 19382
rect 8300 19236 8352 19242
rect 8128 19196 8300 19224
rect 8220 18970 8248 19196
rect 8300 19178 8352 19184
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8116 18624 8168 18630
rect 8300 18624 8352 18630
rect 8116 18566 8168 18572
rect 8220 18572 8300 18578
rect 8220 18566 8352 18572
rect 8128 16726 8156 18566
rect 8220 18550 8340 18566
rect 8220 16794 8248 18550
rect 8404 17785 8432 23446
rect 8484 21616 8536 21622
rect 8482 21584 8484 21593
rect 8536 21584 8538 21593
rect 8482 21519 8538 21528
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8496 21146 8524 21354
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8312 16658 8340 16934
rect 8484 16720 8536 16726
rect 8390 16688 8446 16697
rect 8300 16652 8352 16658
rect 8220 16612 8300 16640
rect 8220 16250 8248 16612
rect 8484 16662 8536 16668
rect 8390 16623 8446 16632
rect 8300 16594 8352 16600
rect 8404 16590 8432 16623
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 16250 8432 16526
rect 8496 16250 8524 16662
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8114 15736 8170 15745
rect 8114 15671 8116 15680
rect 8168 15671 8170 15680
rect 8116 15642 8168 15648
rect 8680 15162 8708 15982
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8772 14657 8800 24806
rect 9324 24682 9352 25094
rect 8944 24676 8996 24682
rect 8944 24618 8996 24624
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 8956 24585 8984 24618
rect 9128 24608 9180 24614
rect 8942 24576 8998 24585
rect 9128 24550 9180 24556
rect 8942 24511 8998 24520
rect 8956 24070 8984 24511
rect 8944 24064 8996 24070
rect 8944 24006 8996 24012
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8864 22166 8892 23802
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21554 8984 21830
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8864 20806 8892 21286
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8956 20330 8984 21490
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 18426 9076 18770
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9140 17882 9168 24550
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9232 23186 9260 23598
rect 9324 23594 9352 24618
rect 9416 24410 9444 25162
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9312 23588 9364 23594
rect 9312 23530 9364 23536
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9232 22778 9260 23122
rect 9324 22982 9352 23530
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9324 22098 9352 22918
rect 9588 22568 9640 22574
rect 9692 22556 9720 24822
rect 9640 22528 9720 22556
rect 9588 22510 9640 22516
rect 9600 22234 9628 22510
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9324 21146 9352 22034
rect 9508 21690 9536 22102
rect 9784 21944 9812 27520
rect 10336 25786 10364 27520
rect 9968 25758 10364 25786
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9692 21916 9812 21944
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9310 20496 9366 20505
rect 9310 20431 9312 20440
rect 9364 20431 9366 20440
rect 9312 20402 9364 20408
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9416 20058 9444 20266
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9416 19514 9444 19994
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18086 9536 19110
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9508 17728 9536 18022
rect 9600 17882 9628 18090
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9588 17740 9640 17746
rect 9508 17700 9588 17728
rect 9588 17682 9640 17688
rect 9600 17202 9628 17682
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9692 16810 9720 21916
rect 9876 21486 9904 24006
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 21049 9812 21286
rect 9876 21146 9904 21422
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9770 21040 9826 21049
rect 9770 20975 9826 20984
rect 9770 18864 9826 18873
rect 9770 18799 9826 18808
rect 9784 18698 9812 18799
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9876 17134 9904 21082
rect 9968 17921 9996 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10152 24818 10180 25298
rect 10244 24954 10272 25366
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10428 24886 10456 25230
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 10060 21962 10088 24618
rect 10152 24410 10180 24754
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24410 10732 24618
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10152 23866 10180 24346
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10152 23254 10180 23802
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10152 22574 10180 23190
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10152 21706 10180 21966
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10060 21678 10180 21706
rect 10060 21146 10088 21678
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10060 18329 10088 21082
rect 10152 19310 10180 21558
rect 10704 21554 10732 21830
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21078 10732 21490
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10704 20602 10732 21014
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20538
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 19514 10548 19790
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10520 19310 10548 19450
rect 10888 19360 10916 27520
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 10980 23304 11008 24822
rect 11060 23316 11112 23322
rect 10980 23276 11060 23304
rect 11060 23258 11112 23264
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10980 22506 11008 23122
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 10980 21078 11008 22442
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 10980 20584 11008 21014
rect 11060 20596 11112 20602
rect 10980 20556 11060 20584
rect 10980 20505 11008 20556
rect 11060 20538 11112 20544
rect 10966 20496 11022 20505
rect 10966 20431 11022 20440
rect 10796 19332 10916 19360
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10046 18320 10102 18329
rect 10046 18255 10102 18264
rect 9954 17912 10010 17921
rect 9954 17847 10010 17856
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9772 16992 9824 16998
rect 9770 16960 9772 16969
rect 9824 16960 9826 16969
rect 9770 16895 9826 16904
rect 9692 16782 9812 16810
rect 9876 16794 9904 17070
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9586 16552 9642 16561
rect 9586 16487 9642 16496
rect 9600 16250 9628 16487
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 8758 14648 8814 14657
rect 9140 14618 9168 15506
rect 9508 14618 9536 15574
rect 9600 15366 9628 15914
rect 9692 15910 9720 16594
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15434 9720 15846
rect 9784 15586 9812 16782
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9968 16658 9996 17682
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10060 16266 10088 18255
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 10152 16726 10180 17206
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16810 10824 19332
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 10968 19168 11020 19174
rect 10966 19136 10968 19145
rect 11020 19136 11022 19145
rect 10966 19071 11022 19080
rect 11348 18970 11376 19246
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18086 11100 18702
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10888 17338 10916 18022
rect 11072 17882 11100 18022
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10966 17096 11022 17105
rect 10966 17031 11022 17040
rect 10704 16782 10824 16810
rect 10980 16794 11008 17031
rect 10968 16788 11020 16794
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10060 16238 10180 16266
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10060 15706 10088 16050
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15638 10180 16238
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15632 10192 15638
rect 9784 15558 9996 15586
rect 10140 15574 10192 15580
rect 10322 15600 10378 15609
rect 9864 15496 9916 15502
rect 9784 15456 9864 15484
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 15360 9640 15366
rect 9640 15308 9720 15314
rect 9588 15302 9720 15308
rect 9600 15286 9720 15302
rect 9692 14822 9720 15286
rect 9784 15094 9812 15456
rect 9864 15438 9916 15444
rect 9968 15201 9996 15558
rect 10322 15535 10324 15544
rect 10376 15535 10378 15544
rect 10324 15506 10376 15512
rect 9954 15192 10010 15201
rect 9954 15127 10010 15136
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 8758 14583 8814 14592
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9692 14482 9720 14758
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 13870 8248 14350
rect 9692 14074 9720 14418
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8128 13190 8156 13738
rect 8220 13530 8248 13806
rect 9784 13705 9812 15030
rect 10336 14958 10364 15506
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 10324 14952 10376 14958
rect 10704 14929 10732 16782
rect 10968 16730 11020 16736
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10796 15638 10824 16662
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11164 16114 11192 16594
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10324 14894 10376 14900
rect 10690 14920 10746 14929
rect 9876 14414 9904 14894
rect 10690 14855 10746 14864
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 14113 11376 14214
rect 11334 14104 11390 14113
rect 11334 14039 11390 14048
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 10138 13968 10194 13977
rect 9770 13696 9826 13705
rect 9770 13631 9826 13640
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12782 8156 13126
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8208 12640 8260 12646
rect 9036 12640 9088 12646
rect 8208 12582 8260 12588
rect 9034 12608 9036 12617
rect 9088 12608 9090 12617
rect 8220 12170 8248 12582
rect 9034 12543 9090 12552
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9588 12436 9640 12442
rect 9692 12424 9720 12854
rect 9640 12396 9720 12424
rect 9588 12378 9640 12384
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8484 12232 8536 12238
rect 8482 12200 8484 12209
rect 8536 12200 8538 12209
rect 8208 12164 8260 12170
rect 8482 12135 8538 12144
rect 8208 12106 8260 12112
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 10169 8156 12038
rect 8496 11898 8524 12135
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8390 11520 8446 11529
rect 8390 11455 8446 11464
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10588 8340 11086
rect 8404 10742 8432 11455
rect 8588 11354 8616 12242
rect 8864 11354 8892 12378
rect 9784 12322 9812 13330
rect 9876 12481 9904 13942
rect 10138 13903 10194 13912
rect 10152 13870 10180 13903
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 10060 13190 10088 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9600 12306 9812 12322
rect 9588 12300 9812 12306
rect 9640 12294 9812 12300
rect 9588 12242 9640 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11558 9812 12174
rect 10060 12102 10088 13126
rect 10520 12986 10548 13330
rect 11256 13297 11284 13670
rect 11242 13288 11298 13297
rect 11242 13223 11298 13232
rect 11440 13002 11468 27520
rect 11612 24336 11664 24342
rect 11612 24278 11664 24284
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11532 23769 11560 24142
rect 11624 23866 11652 24278
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11716 23866 11744 24142
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11518 23760 11574 23769
rect 11518 23695 11520 23704
rect 11572 23695 11574 23704
rect 11520 23666 11572 23672
rect 11624 23633 11652 23802
rect 11610 23624 11666 23633
rect 11610 23559 11666 23568
rect 11716 23526 11744 23802
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11702 22672 11758 22681
rect 11702 22607 11758 22616
rect 11716 22030 11744 22607
rect 11886 22536 11942 22545
rect 11886 22471 11942 22480
rect 11900 22098 11928 22471
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11716 21690 11744 21966
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11900 21350 11928 22034
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11716 19990 11744 21286
rect 11704 19984 11756 19990
rect 11518 19952 11574 19961
rect 11704 19926 11756 19932
rect 11518 19887 11520 19896
rect 11572 19887 11574 19896
rect 11520 19858 11572 19864
rect 11532 19514 11560 19858
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11716 18902 11744 19926
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18086 11836 18770
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11624 16250 11652 16730
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11808 16017 11836 18022
rect 11794 16008 11850 16017
rect 11794 15943 11850 15952
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11164 12974 11468 13002
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12096 10100 12102
rect 10704 12073 10732 12854
rect 10980 12442 11008 12922
rect 11058 12880 11114 12889
rect 11058 12815 11060 12824
rect 11112 12815 11114 12824
rect 11060 12786 11112 12792
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11072 12306 11100 12650
rect 11164 12646 11192 12974
rect 11992 12764 12020 27520
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12452 24410 12480 24686
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12452 23338 12480 24210
rect 12360 23322 12480 23338
rect 12348 23316 12480 23322
rect 12400 23310 12480 23316
rect 12348 23258 12400 23264
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12176 22506 12204 23054
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 12360 21962 12388 23258
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12452 21185 12480 21966
rect 12438 21176 12494 21185
rect 12438 21111 12494 21120
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 20482 12388 20742
rect 12452 20602 12480 20878
rect 12544 20874 12572 27520
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12728 23186 12756 23462
rect 12716 23180 12768 23186
rect 12716 23122 12768 23128
rect 12728 22438 12756 23122
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12728 22098 12756 22374
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12728 21622 12756 22034
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12820 21486 12848 25230
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12912 24682 12940 24754
rect 13004 24682 13032 24822
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 12912 21690 12940 24618
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13004 22506 13032 23462
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12992 21956 13044 21962
rect 12992 21898 13044 21904
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 21146 12848 21422
rect 12912 21146 12940 21490
rect 13004 21418 13032 21898
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12360 20454 12572 20482
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 19854 12388 20334
rect 12544 20330 12572 20454
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12544 20058 12572 20266
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12176 19174 12204 19790
rect 12544 19666 12572 19994
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12360 19638 12572 19666
rect 12360 19310 12388 19638
rect 12728 19378 12756 19790
rect 13004 19718 13032 21014
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12348 19304 12400 19310
rect 12992 19304 13044 19310
rect 12348 19246 12400 19252
rect 12990 19272 12992 19281
rect 13044 19272 13046 19281
rect 12990 19207 13046 19216
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18970 12204 19110
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12268 18426 12296 18838
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12452 17882 12480 18702
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17134 12204 17614
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12176 16658 12204 17070
rect 12452 16998 12480 17818
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16726 12480 16934
rect 12544 16794 12572 17070
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12452 15706 12480 16662
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 11256 12736 12020 12764
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10048 12038 10100 12044
rect 10690 12064 10746 12073
rect 10060 11558 10088 12038
rect 10690 11999 10746 12008
rect 10690 11928 10746 11937
rect 10690 11863 10746 11872
rect 10230 11792 10286 11801
rect 10230 11727 10286 11736
rect 10244 11694 10272 11727
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9588 11552 9640 11558
rect 9772 11552 9824 11558
rect 9588 11494 9640 11500
rect 9678 11520 9734 11529
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8312 10560 8432 10588
rect 8298 10296 8354 10305
rect 8298 10231 8354 10240
rect 8208 10192 8260 10198
rect 8114 10160 8170 10169
rect 8208 10134 8260 10140
rect 8114 10095 8170 10104
rect 8220 9518 8248 10134
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8312 8634 8340 10231
rect 8404 9926 8432 10560
rect 9600 10520 9628 11494
rect 9772 11494 9824 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9678 11455 9734 11464
rect 9692 11286 9720 11455
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 10060 11150 10088 11494
rect 10048 11144 10100 11150
rect 10152 11121 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11257 10732 11863
rect 10690 11248 10746 11257
rect 10690 11183 10746 11192
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10232 11144 10284 11150
rect 10048 11086 10100 11092
rect 10138 11112 10194 11121
rect 10232 11086 10284 11092
rect 10138 11047 10194 11056
rect 10244 10538 10272 11086
rect 11072 10810 11100 11154
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 9680 10532 9732 10538
rect 9600 10492 9680 10520
rect 9680 10474 9732 10480
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 9692 10266 9720 10474
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 9128 9920 9180 9926
rect 9692 9897 9720 10202
rect 9876 10062 9904 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9128 9862 9180 9868
rect 9678 9888 9734 9897
rect 8404 9586 8432 9862
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8404 9178 8432 9522
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8514 8432 9114
rect 8220 8486 8432 8514
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7760 8294 7788 8366
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7748 8016 7800 8022
rect 7746 7984 7748 7993
rect 7800 7984 7802 7993
rect 8220 7954 8248 8486
rect 8588 8401 8616 9590
rect 9140 9586 9168 9862
rect 9678 9823 9734 9832
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9034 9480 9090 9489
rect 9034 9415 9036 9424
rect 9088 9415 9090 9424
rect 9036 9386 9088 9392
rect 8574 8392 8630 8401
rect 9140 8362 9168 9522
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8362 9536 8774
rect 9784 8634 9812 9114
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8514 9904 9998
rect 10888 9586 10916 10066
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9353 10732 9386
rect 10690 9344 10746 9353
rect 10289 9276 10585 9296
rect 10690 9279 10746 9288
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10690 9208 10746 9217
rect 10888 9178 10916 9522
rect 11256 9450 11284 12736
rect 11334 12200 11390 12209
rect 11334 12135 11390 12144
rect 11348 11762 11376 12135
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 12714 11248 12770 11257
rect 12714 11183 12716 11192
rect 12768 11183 12770 11192
rect 12716 11154 12768 11160
rect 12728 10810 12756 11154
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 11624 10266 11652 10746
rect 12438 10568 12494 10577
rect 12438 10503 12440 10512
rect 12492 10503 12494 10512
rect 12440 10474 12492 10480
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10690 9143 10692 9152
rect 10744 9143 10746 9152
rect 10876 9172 10928 9178
rect 10692 9114 10744 9120
rect 10876 9114 10928 9120
rect 10230 9072 10286 9081
rect 9956 9036 10008 9042
rect 10230 9007 10286 9016
rect 9956 8978 10008 8984
rect 9784 8486 9904 8514
rect 9784 8430 9812 8486
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 8574 8327 8630 8336
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9784 7954 9812 8366
rect 9968 8022 9996 8978
rect 10244 8974 10272 9007
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 7746 7919 7802 7928
rect 8208 7948 8260 7954
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7274 7420 7754
rect 7760 7546 7788 7919
rect 8208 7890 8260 7896
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7208 7002 7236 7210
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7208 5914 7236 6938
rect 7852 6934 7880 7822
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7342 8524 7686
rect 9784 7342 9812 7890
rect 9968 7546 9996 7958
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 8496 7002 8524 7278
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7852 6458 7880 6870
rect 10152 6866 10180 8774
rect 10244 8634 10272 8910
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7954 10732 8774
rect 10888 8634 10916 9114
rect 11624 9110 11652 10202
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11716 9178 11744 9590
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 8106 11008 8298
rect 10980 8090 11100 8106
rect 10980 8084 11112 8090
rect 10980 8078 11060 8084
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10704 7206 10732 7890
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7852 5914 7880 6394
rect 9784 6225 9812 6598
rect 10060 6458 10088 6802
rect 10152 6458 10180 6802
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10336 6390 10364 6802
rect 10324 6384 10376 6390
rect 10704 6361 10732 7142
rect 10980 6866 11008 8078
rect 11060 8026 11112 8032
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10324 6326 10376 6332
rect 10690 6352 10746 6361
rect 10690 6287 10746 6296
rect 9770 6216 9826 6225
rect 9770 6151 9826 6160
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 11348 4593 11376 8774
rect 11624 8090 11652 9046
rect 11716 8566 11744 9114
rect 11808 8974 11836 9318
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8634 11836 8910
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 12820 5817 12848 17274
rect 13004 16726 13032 18226
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13004 16250 13032 16662
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13096 7993 13124 27520
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13280 24410 13308 24550
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13372 23866 13400 24618
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13372 22778 13400 23802
rect 13464 23594 13492 24006
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13464 22982 13492 23530
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13174 21312 13230 21321
rect 13174 21247 13230 21256
rect 13188 20806 13216 21247
rect 13280 21078 13308 22374
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21350 13400 21966
rect 13464 21554 13492 22918
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 21894 13584 22374
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13268 20868 13320 20874
rect 13268 20810 13320 20816
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13188 18426 13216 18770
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13174 16824 13230 16833
rect 13174 16759 13230 16768
rect 13188 15978 13216 16759
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13188 15706 13216 15914
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 9217 13308 20810
rect 13372 12753 13400 21286
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18193 13492 18566
rect 13450 18184 13506 18193
rect 13450 18119 13506 18128
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 17134 13584 17478
rect 13648 17338 13676 27520
rect 13726 24168 13782 24177
rect 13726 24103 13782 24112
rect 13740 22098 13768 24103
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 14016 21486 14044 22102
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 14016 21049 14044 21422
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14002 21040 14058 21049
rect 13820 21004 13872 21010
rect 14002 20975 14058 20984
rect 13820 20946 13872 20952
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13740 20058 13768 20878
rect 13832 20602 13860 20946
rect 14108 20806 14136 21354
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20641 14136 20742
rect 14094 20632 14150 20641
rect 13820 20596 13872 20602
rect 14094 20567 14150 20576
rect 13820 20538 13872 20544
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13740 19310 13768 19994
rect 13832 19990 13860 20198
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 18426 13952 19246
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 18154 14044 18702
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14016 17542 14044 18090
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 14016 16794 14044 17478
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14292 14550 14320 27520
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14384 23769 14412 24618
rect 14370 23760 14426 23769
rect 14370 23695 14426 23704
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14568 21350 14596 22170
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 21554 14688 21830
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14568 20806 14596 21286
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14660 20330 14688 21490
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14660 20058 14688 20266
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14660 17338 14688 17818
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15609 14504 15846
rect 14462 15600 14518 15609
rect 14462 15535 14518 15544
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 13358 12744 13414 12753
rect 13358 12679 13414 12688
rect 14108 9722 14136 14486
rect 14844 11121 14872 27520
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24426 15332 25094
rect 15396 24834 15424 27520
rect 15396 24806 15700 24834
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15304 24398 15424 24426
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23526 15332 24210
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15304 23225 15332 23462
rect 15290 23216 15346 23225
rect 15396 23186 15424 24398
rect 15580 23254 15608 24686
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15290 23151 15346 23160
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22778 15424 23122
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15488 22001 15516 22034
rect 15474 21992 15530 22001
rect 15474 21927 15530 21936
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15488 21690 15516 21927
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 15028 21146 15056 21558
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15120 21185 15148 21286
rect 15106 21176 15162 21185
rect 15016 21140 15068 21146
rect 15106 21111 15162 21120
rect 15016 21082 15068 21088
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 18902 15332 20742
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 19514 15424 20266
rect 15488 19718 15516 20946
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15488 19281 15516 19654
rect 15474 19272 15530 19281
rect 15474 19207 15530 19216
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18426 15332 18702
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15304 18306 15332 18362
rect 15212 18278 15332 18306
rect 15212 17882 15240 18278
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 16794 15332 18090
rect 15580 18086 15608 18770
rect 15568 18080 15620 18086
rect 15566 18048 15568 18057
rect 15620 18048 15622 18057
rect 15566 17983 15622 17992
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15396 17338 15424 17682
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15672 12345 15700 24806
rect 15948 23798 15976 27520
rect 16500 24682 16528 27520
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 17052 24410 17080 27520
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16592 23866 16620 24210
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 16854 23760 16910 23769
rect 16854 23695 16910 23704
rect 16868 23662 16896 23695
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16040 23118 16068 23598
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23168 16528 23530
rect 17604 23322 17632 27520
rect 18156 23746 18184 27520
rect 17788 23718 18184 23746
rect 18418 23760 18474 23769
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 16580 23180 16632 23186
rect 16500 23140 16580 23168
rect 16580 23122 16632 23128
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 16028 23112 16080 23118
rect 16026 23080 16028 23089
rect 16080 23080 16082 23089
rect 16026 23015 16082 23024
rect 16592 22778 16620 23122
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 17696 22506 17724 23122
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 22166 16252 22374
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16210 21584 16266 21593
rect 16684 21554 16712 22442
rect 17788 22438 17816 23718
rect 18418 23695 18474 23704
rect 17866 23488 17922 23497
rect 17866 23423 17922 23432
rect 17880 23322 17908 23423
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17880 22098 17908 22510
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 16210 21519 16212 21528
rect 16264 21519 16266 21528
rect 16672 21548 16724 21554
rect 16212 21490 16264 21496
rect 16672 21490 16724 21496
rect 17144 21486 17172 21966
rect 17132 21480 17184 21486
rect 17130 21448 17132 21457
rect 17184 21448 17186 21457
rect 17130 21383 17186 21392
rect 17788 21350 17816 21966
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17776 21344 17828 21350
rect 17774 21312 17776 21321
rect 17828 21312 17830 21321
rect 17774 21247 17830 21256
rect 17500 21072 17552 21078
rect 16486 21040 16542 21049
rect 16486 20975 16542 20984
rect 17498 21040 17500 21049
rect 17552 21040 17554 21049
rect 17498 20975 17554 20984
rect 17592 21004 17644 21010
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16040 19990 16068 20538
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16224 19854 16252 20334
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16224 19242 16252 19790
rect 16212 19236 16264 19242
rect 16132 19196 16212 19224
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15948 18426 15976 18838
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16132 17746 16160 19196
rect 16212 19178 16264 19184
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16210 18456 16266 18465
rect 16210 18391 16212 18400
rect 16264 18391 16266 18400
rect 16212 18362 16264 18368
rect 16316 18154 16344 18566
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16794 15792 17070
rect 16026 16960 16082 16969
rect 16026 16895 16082 16904
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16040 16250 16068 16895
rect 16132 16658 16160 17682
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16500 15978 16528 20975
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17052 20262 17080 20878
rect 17512 20602 17540 20975
rect 17592 20946 17644 20952
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16592 19310 16620 19926
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 18154 16712 18634
rect 17052 18329 17080 20198
rect 17604 20058 17632 20946
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17788 19378 17816 20198
rect 17972 20058 18000 20742
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18834 17816 19178
rect 18064 19145 18092 21422
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 18156 19310 18184 19926
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18432 19242 18460 23695
rect 18708 22778 18736 27520
rect 19062 23624 19118 23633
rect 19062 23559 19118 23568
rect 19076 23322 19104 23559
rect 19260 23497 19288 27520
rect 19812 25786 19840 27520
rect 19536 25758 19840 25786
rect 19246 23488 19302 23497
rect 19246 23423 19302 23432
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18800 22438 18828 23122
rect 19536 22778 19564 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19982 24848 20038 24857
rect 19982 24783 20038 24792
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18800 21078 18828 22374
rect 19168 21554 19196 22510
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19352 21622 19380 22034
rect 19996 21690 20024 24783
rect 20364 21962 20392 27520
rect 20916 23633 20944 27520
rect 21560 24857 21588 27520
rect 21546 24848 21602 24857
rect 21546 24783 21602 24792
rect 21914 24440 21970 24449
rect 21914 24375 21970 24384
rect 21928 24342 21956 24375
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21270 23896 21326 23905
rect 21270 23831 21326 23840
rect 20902 23624 20958 23633
rect 20902 23559 20958 23568
rect 21086 23624 21142 23633
rect 21086 23559 21142 23568
rect 20626 23488 20682 23497
rect 20626 23423 20682 23432
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20640 21690 20668 23423
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20466 18736 20742
rect 19076 20602 19104 20946
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19352 20466 19380 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 20058 18644 20198
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18708 19174 18736 20402
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20456 19990 20484 21422
rect 21100 21146 21128 23559
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21100 20466 21128 20946
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19076 19378 19104 19858
rect 20732 19825 20760 20198
rect 21284 20058 21312 23831
rect 21652 23769 21680 24142
rect 21928 23866 21956 24278
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21638 23760 21694 23769
rect 21638 23695 21694 23704
rect 22006 23760 22062 23769
rect 22006 23695 22008 23704
rect 22060 23695 22062 23704
rect 22008 23666 22060 23672
rect 22112 23497 22140 27520
rect 22190 23760 22246 23769
rect 22190 23695 22246 23704
rect 22098 23488 22154 23497
rect 22098 23423 22154 23432
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22112 22438 22140 23122
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 21100 19514 21128 19858
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 19154 19408 19210 19417
rect 19064 19372 19116 19378
rect 19154 19343 19210 19352
rect 19064 19314 19116 19320
rect 18696 19168 18748 19174
rect 18050 19136 18106 19145
rect 18696 19110 18748 19116
rect 18050 19071 18106 19080
rect 18708 18902 18736 19110
rect 19076 19009 19104 19314
rect 19062 19000 19118 19009
rect 19168 18970 19196 19343
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19062 18935 19118 18944
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18696 18896 18748 18902
rect 20456 18873 20484 19110
rect 21100 18902 21128 19450
rect 21088 18896 21140 18902
rect 18696 18838 18748 18844
rect 20442 18864 20498 18873
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 18426 17816 18770
rect 18142 18728 18198 18737
rect 18142 18663 18198 18672
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17038 18320 17094 18329
rect 17038 18255 17094 18264
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16776 17882 16804 18090
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16776 17134 16804 17818
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17788 17338 17816 17614
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 18156 17270 18184 18663
rect 18340 18426 18368 18838
rect 21088 18838 21140 18844
rect 20442 18799 20498 18808
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20916 18601 20944 18770
rect 22112 18737 22140 22374
rect 22204 19174 22232 23695
rect 22664 23633 22692 27520
rect 23018 24168 23074 24177
rect 23018 24103 23020 24112
rect 23072 24103 23074 24112
rect 23020 24074 23072 24080
rect 23216 23905 23244 27520
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23202 23896 23258 23905
rect 23202 23831 23258 23840
rect 23480 23656 23532 23662
rect 22650 23624 22706 23633
rect 23480 23598 23532 23604
rect 22650 23559 22706 23568
rect 23492 23254 23520 23598
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23584 22642 23612 23530
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22098 18728 22154 18737
rect 22098 18663 22154 18672
rect 20902 18592 20958 18601
rect 20902 18527 20958 18536
rect 20916 18426 20944 18527
rect 22296 18465 22324 22510
rect 23676 22148 23704 25162
rect 23768 23769 23796 27520
rect 24320 25226 24348 27520
rect 24308 25220 24360 25226
rect 24308 25162 24360 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23754 23760 23810 23769
rect 23754 23695 23810 23704
rect 23952 23662 23980 24006
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24044 23594 24072 24210
rect 24122 24168 24178 24177
rect 24122 24103 24178 24112
rect 24136 23866 24164 24103
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24872 23746 24900 27520
rect 25424 24410 25452 27520
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25976 24177 26004 27520
rect 25962 24168 26018 24177
rect 25962 24103 26018 24112
rect 26528 23866 26556 27520
rect 26516 23860 26568 23866
rect 26516 23802 26568 23808
rect 24872 23718 25084 23746
rect 24860 23656 24912 23662
rect 24780 23604 24860 23610
rect 24780 23598 24912 23604
rect 24032 23588 24084 23594
rect 24032 23530 24084 23536
rect 24780 23582 24900 23598
rect 24780 23254 24808 23582
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23768 22420 23796 23122
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 23848 22432 23900 22438
rect 23768 22392 23848 22420
rect 23848 22374 23900 22380
rect 23400 22120 23704 22148
rect 23400 20058 23428 22120
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22848 19174 22876 19858
rect 22926 19408 22982 19417
rect 22926 19343 22982 19352
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22282 18456 22338 18465
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 20904 18420 20956 18426
rect 22282 18391 22338 18400
rect 20904 18362 20956 18368
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21730 18184 21786 18193
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 18616 16998 18644 17478
rect 21284 17105 21312 18158
rect 21730 18119 21786 18128
rect 21744 17746 21772 18119
rect 22756 18086 22784 18770
rect 22848 18290 22876 19110
rect 22940 18970 22968 19343
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22100 18080 22152 18086
rect 22020 18028 22100 18034
rect 22020 18022 22152 18028
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22020 18006 22140 18022
rect 22020 17814 22048 18006
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 17338 21772 17682
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 17408 16992 17460 16998
rect 18604 16992 18656 16998
rect 17408 16934 17460 16940
rect 18602 16960 18604 16969
rect 18656 16960 18658 16969
rect 16868 16658 16896 16934
rect 17420 16833 17448 16934
rect 18602 16895 18658 16904
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 17406 16824 17462 16833
rect 19622 16816 19918 16836
rect 17406 16759 17408 16768
rect 17460 16759 17462 16768
rect 17408 16730 17460 16736
rect 17420 16699 17448 16730
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16592 16250 16620 16594
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16868 16114 16896 16594
rect 23860 16561 23888 22374
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24122 21040 24178 21049
rect 24122 20975 24178 20984
rect 23846 16552 23902 16561
rect 23846 16487 23902 16496
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15065 15792 15846
rect 16500 15706 16528 15914
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 15750 15056 15806 15065
rect 15750 14991 15806 15000
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 24136 14521 24164 20975
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 25056 19417 25084 23718
rect 27080 21457 27108 27520
rect 27632 24449 27660 27520
rect 27618 24440 27674 24449
rect 27618 24375 27674 24384
rect 27066 21448 27122 21457
rect 27066 21383 27122 21392
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24122 14512 24178 14521
rect 24122 14447 24178 14456
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 15658 12336 15714 12345
rect 15658 12271 15714 12280
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14292 9353 14320 9658
rect 13910 9344 13966 9353
rect 13910 9279 13966 9288
rect 14278 9344 14334 9353
rect 14278 9279 14334 9288
rect 13266 9208 13322 9217
rect 13266 9143 13322 9152
rect 13082 7984 13138 7993
rect 13082 7919 13138 7928
rect 12806 5808 12862 5817
rect 12806 5743 12862 5752
rect 11334 4584 11390 4593
rect 11334 4519 11390 4528
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 7010 3496 7066 3505
rect 7010 3431 7066 3440
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 13924 480 13952 9279
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 23478 9072 23534 9081
rect 23478 9007 23534 9016
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 23492 7041 23520 9007
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23478 7032 23534 7041
rect 23478 6967 23534 6976
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 23202 6352 23258 6361
rect 23202 6287 23258 6296
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 23216 480 23244 6287
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 3054 368 3110 377
rect 3054 303 3110 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
<< via2 >>
rect 3330 27648 3386 27704
rect 294 23704 350 23760
rect 1582 23432 1638 23488
rect 1674 22752 1730 22808
rect 2778 24520 2834 24576
rect 2778 24384 2834 24440
rect 2962 26424 3018 26480
rect 3238 25200 3294 25256
rect 2686 22616 2742 22672
rect 2502 21956 2558 21992
rect 2502 21936 2504 21956
rect 2504 21936 2556 21956
rect 2556 21936 2558 21956
rect 1858 18536 1914 18592
rect 2502 18808 2558 18864
rect 2134 18692 2190 18728
rect 2134 18672 2136 18692
rect 2136 18672 2188 18692
rect 2188 18672 2190 18692
rect 2318 17720 2374 17776
rect 1858 17040 1914 17096
rect 1766 10376 1822 10432
rect 1582 7520 1638 7576
rect 2962 15680 3018 15736
rect 2686 15544 2742 15600
rect 2870 15444 2872 15464
rect 2872 15444 2924 15464
rect 2924 15444 2926 15464
rect 2870 15408 2926 15444
rect 2686 15136 2742 15192
rect 3146 18808 3202 18864
rect 3146 18264 3202 18320
rect 4066 27104 4122 27160
rect 3698 25880 3754 25936
rect 3606 23024 3662 23080
rect 3514 20168 3570 20224
rect 3790 23296 3846 23352
rect 4158 24384 4214 24440
rect 4066 23976 4122 24032
rect 4066 22616 4122 22672
rect 3882 21528 3938 21584
rect 4434 23704 4490 23760
rect 4526 22208 4582 22264
rect 5170 23160 5226 23216
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4066 20440 4122 20496
rect 3882 20032 3938 20088
rect 4066 19760 4122 19816
rect 4066 17856 4122 17912
rect 2410 13368 2466 13424
rect 2226 13232 2282 13288
rect 1674 7384 1730 7440
rect 2042 6196 2044 6216
rect 2044 6196 2096 6216
rect 2096 6196 2098 6216
rect 2042 6160 2098 6196
rect 1950 5888 2006 5944
rect 2042 4428 2044 4448
rect 2044 4428 2096 4448
rect 2096 4428 2098 4448
rect 2042 4392 2098 4428
rect 1582 3848 1638 3904
rect 3974 16904 4030 16960
rect 3974 16088 4030 16144
rect 3606 14592 3662 14648
rect 2594 10104 2650 10160
rect 3974 15000 4030 15056
rect 4618 14728 4674 14784
rect 3974 14320 4030 14376
rect 4434 12552 4490 12608
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 3882 11328 3938 11384
rect 3790 10240 3846 10296
rect 3790 9968 3846 10024
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5722 22616 5778 22672
rect 5446 21564 5448 21584
rect 5448 21564 5500 21584
rect 5500 21564 5502 21584
rect 5446 21528 5502 21564
rect 6274 22500 6330 22536
rect 6274 22480 6276 22500
rect 6276 22480 6328 22500
rect 6328 22480 6330 22500
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5538 21140 5594 21176
rect 5538 21120 5540 21140
rect 5540 21120 5592 21140
rect 5592 21120 5594 21140
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5814 19780 5870 19816
rect 5814 19760 5816 19780
rect 5816 19760 5868 19780
rect 5868 19760 5870 19780
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4894 17856 4950 17912
rect 6182 19080 6238 19136
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6182 18128 6238 18184
rect 5262 17312 5318 17368
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6090 17060 6146 17096
rect 6090 17040 6092 17060
rect 6092 17040 6144 17060
rect 6144 17040 6146 17060
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4986 13912 5042 13968
rect 4710 12552 4766 12608
rect 4710 11228 4712 11248
rect 4712 11228 4764 11248
rect 4764 11228 4766 11248
rect 4710 11192 4766 11228
rect 3974 9424 4030 9480
rect 3882 8744 3938 8800
rect 3882 8336 3938 8392
rect 2870 6976 2926 7032
rect 2686 6296 2742 6352
rect 2502 5616 2558 5672
rect 3054 5888 3110 5944
rect 2962 4004 3018 4040
rect 2962 3984 2964 4004
rect 2964 3984 3016 4004
rect 3016 3984 3018 4004
rect 1398 2624 1454 2680
rect 2226 3440 2282 3496
rect 2870 3304 2926 3360
rect 2686 2080 2742 2136
rect 1582 1400 1638 1456
rect 4250 5888 4306 5944
rect 3606 5752 3662 5808
rect 3146 4528 3202 4584
rect 5078 9016 5134 9072
rect 4710 5788 4712 5808
rect 4712 5788 4764 5808
rect 4764 5788 4766 5808
rect 4710 5752 4766 5788
rect 4250 5072 4306 5128
rect 4250 856 4306 912
rect 5262 15156 5318 15192
rect 5262 15136 5264 15156
rect 5264 15136 5316 15156
rect 5316 15136 5318 15156
rect 5262 14476 5318 14512
rect 5262 14456 5264 14476
rect 5264 14456 5316 14476
rect 5316 14456 5318 14476
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6090 15136 6146 15192
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6090 14068 6146 14104
rect 6090 14048 6092 14068
rect 6092 14048 6144 14068
rect 6144 14048 6146 14068
rect 5446 13232 5502 13288
rect 5998 13232 6054 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5354 11464 5410 11520
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6366 14456 6422 14512
rect 6274 11872 6330 11928
rect 5814 11328 5870 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 7194 23704 7250 23760
rect 7102 23296 7158 23352
rect 6918 21392 6974 21448
rect 6918 18692 6974 18728
rect 6918 18672 6920 18692
rect 6920 18672 6972 18692
rect 6972 18672 6974 18692
rect 6550 12824 6606 12880
rect 5722 10512 5778 10568
rect 5262 9968 5318 10024
rect 6826 15544 6882 15600
rect 7010 15428 7066 15464
rect 7010 15408 7012 15428
rect 7012 15408 7064 15428
rect 7064 15408 7066 15428
rect 7654 23568 7710 23624
rect 7378 22500 7434 22536
rect 7378 22480 7380 22500
rect 7380 22480 7432 22500
rect 7432 22480 7434 22500
rect 7378 21528 7434 21584
rect 7562 14864 7618 14920
rect 7194 14728 7250 14784
rect 7102 12280 7158 12336
rect 6458 10376 6514 10432
rect 7654 13404 7656 13424
rect 7656 13404 7708 13424
rect 7708 13404 7710 13424
rect 7654 13368 7710 13404
rect 8114 24692 8116 24712
rect 8116 24692 8168 24712
rect 8168 24692 8170 24712
rect 8114 24656 8170 24692
rect 7930 20032 7986 20088
rect 7930 14864 7986 14920
rect 7930 12280 7986 12336
rect 7746 11736 7802 11792
rect 7378 9968 7434 10024
rect 5998 9868 6000 9888
rect 6000 9868 6052 9888
rect 6052 9868 6054 9888
rect 5998 9832 6054 9868
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5538 8356 5594 8392
rect 5538 8336 5540 8356
rect 5540 8336 5592 8356
rect 5592 8336 5594 8356
rect 5722 8356 5778 8392
rect 5722 8336 5724 8356
rect 5724 8336 5776 8356
rect 5776 8336 5778 8356
rect 6090 8336 6146 8392
rect 5538 8200 5594 8256
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5722 7384 5778 7440
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6918 5616 6974 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5170 3984 5226 4040
rect 7838 9832 7894 9888
rect 8206 22652 8208 22672
rect 8208 22652 8260 22672
rect 8260 22652 8262 22672
rect 8206 22616 8262 22652
rect 8482 21564 8484 21584
rect 8484 21564 8536 21584
rect 8536 21564 8538 21584
rect 8482 21528 8538 21564
rect 8390 17720 8446 17776
rect 8390 16632 8446 16688
rect 8114 15700 8170 15736
rect 8114 15680 8116 15700
rect 8116 15680 8168 15700
rect 8168 15680 8170 15700
rect 8942 24520 8998 24576
rect 9310 20460 9366 20496
rect 9310 20440 9312 20460
rect 9312 20440 9364 20460
rect 9364 20440 9366 20460
rect 9770 20984 9826 21040
rect 9770 18808 9826 18864
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10966 20440 11022 20496
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10046 18264 10102 18320
rect 9954 17856 10010 17912
rect 9770 16940 9772 16960
rect 9772 16940 9824 16960
rect 9824 16940 9826 16960
rect 9770 16904 9826 16940
rect 9586 16496 9642 16552
rect 8758 14592 8814 14648
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10966 19116 10968 19136
rect 10968 19116 11020 19136
rect 11020 19116 11022 19136
rect 10966 19080 11022 19116
rect 10966 17040 11022 17096
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10322 15564 10378 15600
rect 10322 15544 10324 15564
rect 10324 15544 10376 15564
rect 10376 15544 10378 15564
rect 9954 15136 10010 15192
rect 10690 14864 10746 14920
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 11334 14048 11390 14104
rect 9770 13640 9826 13696
rect 9034 12588 9036 12608
rect 9036 12588 9088 12608
rect 9088 12588 9090 12608
rect 9034 12552 9090 12588
rect 8482 12180 8484 12200
rect 8484 12180 8536 12200
rect 8536 12180 8538 12200
rect 8482 12144 8538 12180
rect 8390 11464 8446 11520
rect 10138 13912 10194 13968
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9862 12416 9918 12472
rect 11242 13232 11298 13288
rect 11518 23724 11574 23760
rect 11518 23704 11520 23724
rect 11520 23704 11572 23724
rect 11572 23704 11574 23724
rect 11610 23568 11666 23624
rect 11702 22616 11758 22672
rect 11886 22480 11942 22536
rect 11518 19916 11574 19952
rect 11518 19896 11520 19916
rect 11520 19896 11572 19916
rect 11572 19896 11574 19916
rect 11794 15952 11850 16008
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11058 12844 11114 12880
rect 11058 12824 11060 12844
rect 11060 12824 11112 12844
rect 11112 12824 11114 12844
rect 12438 21120 12494 21176
rect 12990 19252 12992 19272
rect 12992 19252 13044 19272
rect 13044 19252 13046 19272
rect 12990 19216 13046 19252
rect 10690 12008 10746 12064
rect 10690 11872 10746 11928
rect 10230 11736 10286 11792
rect 8298 10240 8354 10296
rect 8114 10104 8170 10160
rect 9678 11464 9734 11520
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10690 11192 10746 11248
rect 10138 11056 10194 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 7746 7964 7748 7984
rect 7748 7964 7800 7984
rect 7800 7964 7802 7984
rect 7746 7928 7802 7964
rect 9678 9832 9734 9888
rect 9034 9444 9090 9480
rect 9034 9424 9036 9444
rect 9036 9424 9088 9444
rect 9088 9424 9090 9444
rect 8574 8336 8630 8392
rect 10690 9288 10746 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10690 9172 10746 9208
rect 11334 12144 11390 12200
rect 12714 11212 12770 11248
rect 12714 11192 12716 11212
rect 12716 11192 12768 11212
rect 12768 11192 12770 11212
rect 12438 10532 12494 10568
rect 12438 10512 12440 10532
rect 12440 10512 12492 10532
rect 12492 10512 12494 10532
rect 10690 9152 10692 9172
rect 10692 9152 10744 9172
rect 10744 9152 10746 9172
rect 10230 9016 10286 9072
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10690 6296 10746 6352
rect 9770 6160 9826 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 13174 21256 13230 21312
rect 13174 16768 13230 16824
rect 13450 18128 13506 18184
rect 13726 24112 13782 24168
rect 14002 20984 14058 21040
rect 14094 20576 14150 20632
rect 14370 23704 14426 23760
rect 14462 15544 14518 15600
rect 13358 12688 13414 12744
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15290 23160 15346 23216
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15474 21936 15530 21992
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15106 21120 15162 21176
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15474 19216 15530 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15566 18028 15568 18048
rect 15568 18028 15620 18048
rect 15620 18028 15622 18048
rect 15566 17992 15622 18028
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 16854 23704 16910 23760
rect 16026 23060 16028 23080
rect 16028 23060 16080 23080
rect 16080 23060 16082 23080
rect 16026 23024 16082 23060
rect 16210 21548 16266 21584
rect 18418 23704 18474 23760
rect 17866 23432 17922 23488
rect 16210 21528 16212 21548
rect 16212 21528 16264 21548
rect 16264 21528 16266 21548
rect 17130 21428 17132 21448
rect 17132 21428 17184 21448
rect 17184 21428 17186 21448
rect 17130 21392 17186 21428
rect 17774 21292 17776 21312
rect 17776 21292 17828 21312
rect 17828 21292 17830 21312
rect 17774 21256 17830 21292
rect 16486 20984 16542 21040
rect 17498 21020 17500 21040
rect 17500 21020 17552 21040
rect 17552 21020 17554 21040
rect 17498 20984 17554 21020
rect 16210 18420 16266 18456
rect 16210 18400 16212 18420
rect 16212 18400 16264 18420
rect 16264 18400 16266 18420
rect 16026 16904 16082 16960
rect 19062 23568 19118 23624
rect 19246 23432 19302 23488
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19982 24792 20038 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 21546 24792 21602 24848
rect 21914 24384 21970 24440
rect 21270 23840 21326 23896
rect 20902 23568 20958 23624
rect 21086 23568 21142 23624
rect 20626 23432 20682 23488
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 21638 23704 21694 23760
rect 22006 23724 22062 23760
rect 22006 23704 22008 23724
rect 22008 23704 22060 23724
rect 22060 23704 22062 23724
rect 22190 23704 22246 23760
rect 22098 23432 22154 23488
rect 20718 19760 20774 19816
rect 19154 19352 19210 19408
rect 18050 19080 18106 19136
rect 19062 18944 19118 19000
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 18142 18672 18198 18728
rect 17038 18264 17094 18320
rect 20442 18808 20498 18864
rect 23018 24132 23074 24168
rect 23018 24112 23020 24132
rect 23020 24112 23072 24132
rect 23072 24112 23074 24132
rect 23202 23840 23258 23896
rect 22650 23568 22706 23624
rect 22098 18672 22154 18728
rect 20902 18536 20958 18592
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 23754 23704 23810 23760
rect 24122 24112 24178 24168
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25962 24112 26018 24168
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 22926 19352 22982 19408
rect 22282 18400 22338 18456
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 21730 18128 21786 18184
rect 21270 17040 21326 17096
rect 18602 16940 18604 16960
rect 18604 16940 18656 16960
rect 18656 16940 18658 16960
rect 18602 16904 18658 16940
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 17406 16788 17462 16824
rect 17406 16768 17408 16788
rect 17408 16768 17460 16788
rect 17460 16768 17462 16788
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24122 20984 24178 21040
rect 23846 16496 23902 16552
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 15750 15000 15806 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 27618 24384 27674 24440
rect 27066 21392 27122 21448
rect 25042 19352 25098 19408
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24122 14456 24178 14512
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 15658 12280 15714 12336
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 14830 11056 14886 11112
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 13910 9288 13966 9344
rect 14278 9288 14334 9344
rect 13266 9152 13322 9208
rect 13082 7928 13138 7984
rect 12806 5752 12862 5808
rect 11334 4528 11390 4584
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 7010 3440 7066 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 23478 9016 23534 9072
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23478 6976 23534 7032
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23202 6296 23258 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 3054 312 3110 368
<< metal3 >>
rect 0 27706 480 27736
rect 3325 27706 3391 27709
rect 0 27704 3391 27706
rect 0 27648 3330 27704
rect 3386 27648 3391 27704
rect 0 27646 3391 27648
rect 0 27616 480 27646
rect 3325 27643 3391 27646
rect 0 27162 480 27192
rect 4061 27162 4127 27165
rect 0 27160 4127 27162
rect 0 27104 4066 27160
rect 4122 27104 4127 27160
rect 0 27102 4127 27104
rect 0 27072 480 27102
rect 4061 27099 4127 27102
rect 0 26482 480 26512
rect 2957 26482 3023 26485
rect 0 26480 3023 26482
rect 0 26424 2962 26480
rect 3018 26424 3023 26480
rect 0 26422 3023 26424
rect 0 26392 480 26422
rect 2957 26419 3023 26422
rect 0 25938 480 25968
rect 3693 25938 3759 25941
rect 0 25936 3759 25938
rect 0 25880 3698 25936
rect 3754 25880 3759 25936
rect 0 25878 3759 25880
rect 0 25848 480 25878
rect 3693 25875 3759 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25258 480 25288
rect 3233 25258 3299 25261
rect 0 25256 3299 25258
rect 0 25200 3238 25256
rect 3294 25200 3299 25256
rect 0 25198 3299 25200
rect 0 25168 480 25198
rect 3233 25195 3299 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 19977 24850 20043 24853
rect 21541 24850 21607 24853
rect 19977 24848 21607 24850
rect 19977 24792 19982 24848
rect 20038 24792 21546 24848
rect 21602 24792 21607 24848
rect 19977 24790 21607 24792
rect 19977 24787 20043 24790
rect 21541 24787 21607 24790
rect 0 24714 480 24744
rect 8109 24714 8175 24717
rect 0 24712 8175 24714
rect 0 24656 8114 24712
rect 8170 24656 8175 24712
rect 0 24654 8175 24656
rect 0 24624 480 24654
rect 8109 24651 8175 24654
rect 2773 24578 2839 24581
rect 8937 24578 9003 24581
rect 2773 24576 9003 24578
rect 2773 24520 2778 24576
rect 2834 24520 8942 24576
rect 8998 24520 9003 24576
rect 2773 24518 9003 24520
rect 2773 24515 2839 24518
rect 8937 24515 9003 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 2773 24442 2839 24445
rect 4153 24442 4219 24445
rect 2773 24440 4219 24442
rect 2773 24384 2778 24440
rect 2834 24384 4158 24440
rect 4214 24384 4219 24440
rect 2773 24382 4219 24384
rect 2773 24379 2839 24382
rect 4153 24379 4219 24382
rect 21909 24442 21975 24445
rect 27613 24442 27679 24445
rect 21909 24440 27679 24442
rect 21909 24384 21914 24440
rect 21970 24384 27618 24440
rect 27674 24384 27679 24440
rect 21909 24382 27679 24384
rect 21909 24379 21975 24382
rect 27613 24379 27679 24382
rect 13721 24170 13787 24173
rect 23013 24170 23079 24173
rect 13721 24168 23079 24170
rect 13721 24112 13726 24168
rect 13782 24112 23018 24168
rect 23074 24112 23079 24168
rect 13721 24110 23079 24112
rect 13721 24107 13787 24110
rect 23013 24107 23079 24110
rect 24117 24170 24183 24173
rect 25957 24170 26023 24173
rect 24117 24168 26023 24170
rect 24117 24112 24122 24168
rect 24178 24112 25962 24168
rect 26018 24112 26023 24168
rect 24117 24110 26023 24112
rect 24117 24107 24183 24110
rect 25957 24107 26023 24110
rect 0 24034 480 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 480 23974
rect 4061 23971 4127 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 21265 23898 21331 23901
rect 23197 23898 23263 23901
rect 21265 23896 23263 23898
rect 21265 23840 21270 23896
rect 21326 23840 23202 23896
rect 23258 23840 23263 23896
rect 21265 23838 23263 23840
rect 21265 23835 21331 23838
rect 23197 23835 23263 23838
rect 289 23762 355 23765
rect 4429 23762 4495 23765
rect 289 23760 4495 23762
rect 289 23704 294 23760
rect 350 23704 4434 23760
rect 4490 23704 4495 23760
rect 289 23702 4495 23704
rect 289 23699 355 23702
rect 4429 23699 4495 23702
rect 7189 23762 7255 23765
rect 11513 23762 11579 23765
rect 7189 23760 11579 23762
rect 7189 23704 7194 23760
rect 7250 23704 11518 23760
rect 11574 23704 11579 23760
rect 7189 23702 11579 23704
rect 7189 23699 7255 23702
rect 11513 23699 11579 23702
rect 14365 23762 14431 23765
rect 16849 23762 16915 23765
rect 14365 23760 16915 23762
rect 14365 23704 14370 23760
rect 14426 23704 16854 23760
rect 16910 23704 16915 23760
rect 14365 23702 16915 23704
rect 14365 23699 14431 23702
rect 16849 23699 16915 23702
rect 18413 23762 18479 23765
rect 21633 23762 21699 23765
rect 22001 23762 22067 23765
rect 18413 23760 22067 23762
rect 18413 23704 18418 23760
rect 18474 23704 21638 23760
rect 21694 23704 22006 23760
rect 22062 23704 22067 23760
rect 18413 23702 22067 23704
rect 18413 23699 18479 23702
rect 21633 23699 21699 23702
rect 22001 23699 22067 23702
rect 22185 23762 22251 23765
rect 23749 23762 23815 23765
rect 22185 23760 23815 23762
rect 22185 23704 22190 23760
rect 22246 23704 23754 23760
rect 23810 23704 23815 23760
rect 22185 23702 23815 23704
rect 22185 23699 22251 23702
rect 23749 23699 23815 23702
rect 7649 23626 7715 23629
rect 11605 23626 11671 23629
rect 7649 23624 11671 23626
rect 7649 23568 7654 23624
rect 7710 23568 11610 23624
rect 11666 23568 11671 23624
rect 7649 23566 11671 23568
rect 7649 23563 7715 23566
rect 11605 23563 11671 23566
rect 19057 23626 19123 23629
rect 20897 23626 20963 23629
rect 19057 23624 20963 23626
rect 19057 23568 19062 23624
rect 19118 23568 20902 23624
rect 20958 23568 20963 23624
rect 19057 23566 20963 23568
rect 19057 23563 19123 23566
rect 20897 23563 20963 23566
rect 21081 23626 21147 23629
rect 22645 23626 22711 23629
rect 21081 23624 22711 23626
rect 21081 23568 21086 23624
rect 21142 23568 22650 23624
rect 22706 23568 22711 23624
rect 21081 23566 22711 23568
rect 21081 23563 21147 23566
rect 22645 23563 22711 23566
rect 0 23490 480 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 480 23430
rect 1577 23427 1643 23430
rect 17861 23490 17927 23493
rect 19241 23490 19307 23493
rect 17861 23488 19307 23490
rect 17861 23432 17866 23488
rect 17922 23432 19246 23488
rect 19302 23432 19307 23488
rect 17861 23430 19307 23432
rect 17861 23427 17927 23430
rect 19241 23427 19307 23430
rect 20621 23490 20687 23493
rect 22093 23490 22159 23493
rect 20621 23488 22159 23490
rect 20621 23432 20626 23488
rect 20682 23432 22098 23488
rect 22154 23432 22159 23488
rect 20621 23430 22159 23432
rect 20621 23427 20687 23430
rect 22093 23427 22159 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 3785 23354 3851 23357
rect 7097 23354 7163 23357
rect 3785 23352 7163 23354
rect 3785 23296 3790 23352
rect 3846 23296 7102 23352
rect 7158 23296 7163 23352
rect 3785 23294 7163 23296
rect 3785 23291 3851 23294
rect 7097 23291 7163 23294
rect 5165 23218 5231 23221
rect 15285 23218 15351 23221
rect 5165 23216 15351 23218
rect 5165 23160 5170 23216
rect 5226 23160 15290 23216
rect 15346 23160 15351 23216
rect 5165 23158 15351 23160
rect 5165 23155 5231 23158
rect 15285 23155 15351 23158
rect 3601 23082 3667 23085
rect 16021 23082 16087 23085
rect 3601 23080 16087 23082
rect 3601 23024 3606 23080
rect 3662 23024 16026 23080
rect 16082 23024 16087 23080
rect 3601 23022 16087 23024
rect 3601 23019 3667 23022
rect 16021 23019 16087 23022
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1669 22810 1735 22813
rect 0 22808 1735 22810
rect 0 22752 1674 22808
rect 1730 22752 1735 22808
rect 0 22750 1735 22752
rect 0 22720 480 22750
rect 1669 22747 1735 22750
rect 2681 22674 2747 22677
rect 4061 22674 4127 22677
rect 5717 22674 5783 22677
rect 2681 22672 3986 22674
rect 2681 22616 2686 22672
rect 2742 22616 3986 22672
rect 2681 22614 3986 22616
rect 2681 22611 2747 22614
rect 3926 22538 3986 22614
rect 4061 22672 5783 22674
rect 4061 22616 4066 22672
rect 4122 22616 5722 22672
rect 5778 22616 5783 22672
rect 4061 22614 5783 22616
rect 4061 22611 4127 22614
rect 5717 22611 5783 22614
rect 8201 22674 8267 22677
rect 11697 22674 11763 22677
rect 8201 22672 11763 22674
rect 8201 22616 8206 22672
rect 8262 22616 11702 22672
rect 11758 22616 11763 22672
rect 8201 22614 11763 22616
rect 8201 22611 8267 22614
rect 11697 22611 11763 22614
rect 6269 22538 6335 22541
rect 3926 22536 6335 22538
rect 3926 22480 6274 22536
rect 6330 22480 6335 22536
rect 3926 22478 6335 22480
rect 6269 22475 6335 22478
rect 7373 22538 7439 22541
rect 11881 22538 11947 22541
rect 7373 22536 11947 22538
rect 7373 22480 7378 22536
rect 7434 22480 11886 22536
rect 11942 22480 11947 22536
rect 7373 22478 11947 22480
rect 7373 22475 7439 22478
rect 11881 22475 11947 22478
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 4521 22266 4587 22269
rect 0 22264 4587 22266
rect 0 22208 4526 22264
rect 4582 22208 4587 22264
rect 0 22206 4587 22208
rect 0 22176 480 22206
rect 4521 22203 4587 22206
rect 2497 21994 2563 21997
rect 15469 21994 15535 21997
rect 2497 21992 15535 21994
rect 2497 21936 2502 21992
rect 2558 21936 15474 21992
rect 15530 21936 15535 21992
rect 2497 21934 15535 21936
rect 2497 21931 2563 21934
rect 15469 21931 15535 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21586 480 21616
rect 3877 21586 3943 21589
rect 0 21584 3943 21586
rect 0 21528 3882 21584
rect 3938 21528 3943 21584
rect 0 21526 3943 21528
rect 0 21496 480 21526
rect 3877 21523 3943 21526
rect 5441 21586 5507 21589
rect 7373 21586 7439 21589
rect 5441 21584 7439 21586
rect 5441 21528 5446 21584
rect 5502 21528 7378 21584
rect 7434 21528 7439 21584
rect 5441 21526 7439 21528
rect 5441 21523 5507 21526
rect 7373 21523 7439 21526
rect 8477 21586 8543 21589
rect 16205 21586 16271 21589
rect 8477 21584 16271 21586
rect 8477 21528 8482 21584
rect 8538 21528 16210 21584
rect 16266 21528 16271 21584
rect 8477 21526 16271 21528
rect 8477 21523 8543 21526
rect 16205 21523 16271 21526
rect 6913 21450 6979 21453
rect 17125 21450 17191 21453
rect 27061 21450 27127 21453
rect 6913 21448 17191 21450
rect 6913 21392 6918 21448
rect 6974 21392 17130 21448
rect 17186 21392 17191 21448
rect 6913 21390 17191 21392
rect 6913 21387 6979 21390
rect 17125 21387 17191 21390
rect 17910 21448 27127 21450
rect 17910 21392 27066 21448
rect 27122 21392 27127 21448
rect 17910 21390 27127 21392
rect 13169 21314 13235 21317
rect 17769 21314 17835 21317
rect 13169 21312 17835 21314
rect 13169 21256 13174 21312
rect 13230 21256 17774 21312
rect 17830 21256 17835 21312
rect 13169 21254 17835 21256
rect 13169 21251 13235 21254
rect 17769 21251 17835 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 5533 21178 5599 21181
rect 12433 21178 12499 21181
rect 15101 21178 15167 21181
rect 17910 21178 17970 21390
rect 27061 21387 27127 21390
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 5533 21176 10058 21178
rect 5533 21120 5538 21176
rect 5594 21120 10058 21176
rect 5533 21118 10058 21120
rect 5533 21115 5599 21118
rect 0 21042 480 21072
rect 9765 21042 9831 21045
rect 0 21040 9831 21042
rect 0 20984 9770 21040
rect 9826 20984 9831 21040
rect 0 20982 9831 20984
rect 9998 21042 10058 21118
rect 12433 21176 15026 21178
rect 12433 21120 12438 21176
rect 12494 21120 15026 21176
rect 12433 21118 15026 21120
rect 12433 21115 12499 21118
rect 13997 21042 14063 21045
rect 9998 21040 14063 21042
rect 9998 20984 14002 21040
rect 14058 20984 14063 21040
rect 9998 20982 14063 20984
rect 14966 21042 15026 21118
rect 15101 21176 17970 21178
rect 15101 21120 15106 21176
rect 15162 21120 17970 21176
rect 15101 21118 17970 21120
rect 15101 21115 15167 21118
rect 16481 21042 16547 21045
rect 17493 21042 17559 21045
rect 14966 21040 17559 21042
rect 14966 20984 16486 21040
rect 16542 20984 17498 21040
rect 17554 20984 17559 21040
rect 14966 20982 17559 20984
rect 0 20952 480 20982
rect 9765 20979 9831 20982
rect 13997 20979 14063 20982
rect 16481 20979 16547 20982
rect 17493 20979 17559 20982
rect 24117 21042 24183 21045
rect 27520 21042 28000 21072
rect 24117 21040 28000 21042
rect 24117 20984 24122 21040
rect 24178 20984 28000 21040
rect 24117 20982 28000 20984
rect 24117 20979 24183 20982
rect 27520 20952 28000 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 14089 20634 14155 20637
rect 6134 20632 14155 20634
rect 6134 20576 14094 20632
rect 14150 20576 14155 20632
rect 6134 20574 14155 20576
rect 4061 20498 4127 20501
rect 6134 20498 6194 20574
rect 14089 20571 14155 20574
rect 4061 20496 6194 20498
rect 4061 20440 4066 20496
rect 4122 20440 6194 20496
rect 4061 20438 6194 20440
rect 9305 20498 9371 20501
rect 10961 20498 11027 20501
rect 9305 20496 11027 20498
rect 9305 20440 9310 20496
rect 9366 20440 10966 20496
rect 11022 20440 11027 20496
rect 9305 20438 11027 20440
rect 4061 20435 4127 20438
rect 9305 20435 9371 20438
rect 10961 20435 11027 20438
rect 0 20362 480 20392
rect 0 20302 3434 20362
rect 9622 20328 9628 20364
rect 0 20272 480 20302
rect 3374 19954 3434 20302
rect 9308 20300 9628 20328
rect 9692 20300 9698 20364
rect 9308 20268 9690 20300
rect 3509 20226 3575 20229
rect 9308 20226 9368 20268
rect 3509 20224 9368 20226
rect 3509 20168 3514 20224
rect 3570 20168 9368 20224
rect 3509 20166 9368 20168
rect 3509 20163 3575 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 3877 20090 3943 20093
rect 7925 20090 7991 20093
rect 3877 20088 7991 20090
rect 3877 20032 3882 20088
rect 3938 20032 7930 20088
rect 7986 20032 7991 20088
rect 3877 20030 7991 20032
rect 3877 20027 3943 20030
rect 7925 20027 7991 20030
rect 11513 19954 11579 19957
rect 3374 19952 11579 19954
rect 3374 19896 11518 19952
rect 11574 19896 11579 19952
rect 3374 19894 11579 19896
rect 11513 19891 11579 19894
rect 0 19818 480 19848
rect 4061 19818 4127 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 480 19758
rect 4061 19755 4127 19758
rect 5809 19818 5875 19821
rect 20713 19818 20779 19821
rect 5809 19816 20779 19818
rect 5809 19760 5814 19816
rect 5870 19760 20718 19816
rect 20774 19760 20779 19816
rect 5809 19758 20779 19760
rect 5809 19755 5875 19758
rect 20713 19755 20779 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 9622 19348 9628 19412
rect 9692 19410 9698 19412
rect 19149 19410 19215 19413
rect 9692 19408 19215 19410
rect 9692 19352 19154 19408
rect 19210 19352 19215 19408
rect 9692 19350 19215 19352
rect 9692 19348 9698 19350
rect 19149 19347 19215 19350
rect 22921 19410 22987 19413
rect 25037 19410 25103 19413
rect 22921 19408 25103 19410
rect 22921 19352 22926 19408
rect 22982 19352 25042 19408
rect 25098 19352 25103 19408
rect 22921 19350 25103 19352
rect 22921 19347 22987 19350
rect 25037 19347 25103 19350
rect 12985 19274 13051 19277
rect 15469 19274 15535 19277
rect 6502 19214 10794 19274
rect 0 19138 480 19168
rect 6177 19138 6243 19141
rect 0 19136 6243 19138
rect 0 19080 6182 19136
rect 6238 19080 6243 19136
rect 0 19078 6243 19080
rect 0 19048 480 19078
rect 6177 19075 6243 19078
rect 2497 18866 2563 18869
rect 3141 18866 3207 18869
rect 2497 18864 3207 18866
rect 2497 18808 2502 18864
rect 2558 18808 3146 18864
rect 3202 18808 3207 18864
rect 2497 18806 3207 18808
rect 2497 18803 2563 18806
rect 3141 18803 3207 18806
rect 2129 18730 2195 18733
rect 6502 18730 6562 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 10734 19002 10794 19214
rect 12985 19272 15535 19274
rect 12985 19216 12990 19272
rect 13046 19216 15474 19272
rect 15530 19216 15535 19272
rect 12985 19214 15535 19216
rect 12985 19211 13051 19214
rect 15469 19211 15535 19214
rect 10961 19138 11027 19141
rect 18045 19138 18111 19141
rect 10961 19136 18111 19138
rect 10961 19080 10966 19136
rect 11022 19080 18050 19136
rect 18106 19080 18111 19136
rect 10961 19078 18111 19080
rect 10961 19075 11027 19078
rect 18045 19075 18111 19078
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 19057 19002 19123 19005
rect 10734 19000 19123 19002
rect 10734 18944 19062 19000
rect 19118 18944 19123 19000
rect 10734 18942 19123 18944
rect 19057 18939 19123 18942
rect 9765 18866 9831 18869
rect 20437 18866 20503 18869
rect 9765 18864 20503 18866
rect 9765 18808 9770 18864
rect 9826 18808 20442 18864
rect 20498 18808 20503 18864
rect 9765 18806 20503 18808
rect 9765 18803 9831 18806
rect 20437 18803 20503 18806
rect 2129 18728 6562 18730
rect 2129 18672 2134 18728
rect 2190 18672 6562 18728
rect 2129 18670 6562 18672
rect 6913 18730 6979 18733
rect 18137 18730 18203 18733
rect 22093 18730 22159 18733
rect 6913 18728 17970 18730
rect 6913 18672 6918 18728
rect 6974 18672 17970 18728
rect 6913 18670 17970 18672
rect 2129 18667 2195 18670
rect 6913 18667 6979 18670
rect 0 18594 480 18624
rect 1853 18594 1919 18597
rect 0 18592 1919 18594
rect 0 18536 1858 18592
rect 1914 18536 1919 18592
rect 0 18534 1919 18536
rect 17910 18594 17970 18670
rect 18137 18728 22159 18730
rect 18137 18672 18142 18728
rect 18198 18672 22098 18728
rect 22154 18672 22159 18728
rect 18137 18670 22159 18672
rect 18137 18667 18203 18670
rect 22093 18667 22159 18670
rect 20897 18594 20963 18597
rect 17910 18592 20963 18594
rect 17910 18536 20902 18592
rect 20958 18536 20963 18592
rect 17910 18534 20963 18536
rect 0 18504 480 18534
rect 1853 18531 1919 18534
rect 20897 18531 20963 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 16205 18458 16271 18461
rect 22277 18458 22343 18461
rect 16205 18456 22343 18458
rect 16205 18400 16210 18456
rect 16266 18400 22282 18456
rect 22338 18400 22343 18456
rect 16205 18398 22343 18400
rect 16205 18395 16271 18398
rect 22277 18395 22343 18398
rect 3141 18322 3207 18325
rect 10041 18322 10107 18325
rect 17033 18322 17099 18325
rect 3141 18320 10107 18322
rect 3141 18264 3146 18320
rect 3202 18264 10046 18320
rect 10102 18264 10107 18320
rect 3141 18262 10107 18264
rect 3141 18259 3207 18262
rect 10041 18259 10107 18262
rect 13310 18320 17099 18322
rect 13310 18264 17038 18320
rect 17094 18264 17099 18320
rect 13310 18262 17099 18264
rect 6177 18186 6243 18189
rect 13310 18186 13370 18262
rect 17033 18259 17099 18262
rect 6177 18184 13370 18186
rect 6177 18128 6182 18184
rect 6238 18128 13370 18184
rect 6177 18126 13370 18128
rect 13445 18186 13511 18189
rect 21725 18186 21791 18189
rect 13445 18184 21791 18186
rect 13445 18128 13450 18184
rect 13506 18128 21730 18184
rect 21786 18128 21791 18184
rect 13445 18126 21791 18128
rect 6177 18123 6243 18126
rect 13445 18123 13511 18126
rect 21725 18123 21791 18126
rect 15561 18052 15627 18053
rect 15510 17988 15516 18052
rect 15580 18050 15627 18052
rect 15580 18048 15672 18050
rect 15622 17992 15672 18048
rect 15580 17990 15672 17992
rect 15580 17988 15627 17990
rect 15561 17987 15627 17988
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 4061 17914 4127 17917
rect 0 17912 4127 17914
rect 0 17856 4066 17912
rect 4122 17856 4127 17912
rect 0 17854 4127 17856
rect 0 17824 480 17854
rect 4061 17851 4127 17854
rect 4889 17914 4955 17917
rect 9949 17914 10015 17917
rect 4889 17912 10015 17914
rect 4889 17856 4894 17912
rect 4950 17856 9954 17912
rect 10010 17856 10015 17912
rect 4889 17854 10015 17856
rect 4889 17851 4955 17854
rect 9949 17851 10015 17854
rect 2313 17778 2379 17781
rect 8385 17778 8451 17781
rect 2313 17776 8451 17778
rect 2313 17720 2318 17776
rect 2374 17720 8390 17776
rect 8446 17720 8451 17776
rect 2313 17718 8451 17720
rect 2313 17715 2379 17718
rect 8385 17715 8451 17718
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 5257 17370 5323 17373
rect 0 17368 5323 17370
rect 0 17312 5262 17368
rect 5318 17312 5323 17368
rect 0 17310 5323 17312
rect 0 17280 480 17310
rect 5257 17307 5323 17310
rect 1853 17098 1919 17101
rect 6085 17098 6151 17101
rect 1853 17096 6151 17098
rect 1853 17040 1858 17096
rect 1914 17040 6090 17096
rect 6146 17040 6151 17096
rect 1853 17038 6151 17040
rect 1853 17035 1919 17038
rect 6085 17035 6151 17038
rect 10961 17098 11027 17101
rect 21265 17098 21331 17101
rect 10961 17096 21331 17098
rect 10961 17040 10966 17096
rect 11022 17040 21270 17096
rect 21326 17040 21331 17096
rect 10961 17038 21331 17040
rect 10961 17035 11027 17038
rect 21265 17035 21331 17038
rect 3969 16962 4035 16965
rect 9765 16962 9831 16965
rect 3969 16960 9831 16962
rect 3969 16904 3974 16960
rect 4030 16904 9770 16960
rect 9826 16904 9831 16960
rect 3969 16902 9831 16904
rect 3969 16899 4035 16902
rect 9765 16899 9831 16902
rect 16021 16962 16087 16965
rect 18597 16962 18663 16965
rect 16021 16960 18663 16962
rect 16021 16904 16026 16960
rect 16082 16904 18602 16960
rect 18658 16904 18663 16960
rect 16021 16902 18663 16904
rect 16021 16899 16087 16902
rect 18597 16899 18663 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 13169 16826 13235 16829
rect 17401 16826 17467 16829
rect 13169 16824 17467 16826
rect 13169 16768 13174 16824
rect 13230 16768 17406 16824
rect 17462 16768 17467 16824
rect 13169 16766 17467 16768
rect 13169 16763 13235 16766
rect 17401 16763 17467 16766
rect 0 16690 480 16720
rect 8385 16690 8451 16693
rect 0 16688 8451 16690
rect 0 16632 8390 16688
rect 8446 16632 8451 16688
rect 0 16630 8451 16632
rect 0 16600 480 16630
rect 8385 16627 8451 16630
rect 9581 16554 9647 16557
rect 23841 16554 23907 16557
rect 9581 16552 23907 16554
rect 9581 16496 9586 16552
rect 9642 16496 23846 16552
rect 23902 16496 23907 16552
rect 9581 16494 23907 16496
rect 9581 16491 9647 16494
rect 23841 16491 23907 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16146 480 16176
rect 3969 16146 4035 16149
rect 0 16144 4035 16146
rect 0 16088 3974 16144
rect 4030 16088 4035 16144
rect 0 16086 4035 16088
rect 0 16056 480 16086
rect 3969 16083 4035 16086
rect 11789 16010 11855 16013
rect 2500 16008 11855 16010
rect 2500 15952 11794 16008
rect 11850 15952 11855 16008
rect 2500 15950 11855 15952
rect 0 15466 480 15496
rect 2500 15466 2560 15950
rect 11789 15947 11855 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 2957 15738 3023 15741
rect 8109 15738 8175 15741
rect 2957 15736 8175 15738
rect 2957 15680 2962 15736
rect 3018 15680 8114 15736
rect 8170 15680 8175 15736
rect 2957 15678 8175 15680
rect 2957 15675 3023 15678
rect 8109 15675 8175 15678
rect 2681 15602 2747 15605
rect 6821 15602 6887 15605
rect 2681 15600 6887 15602
rect 2681 15544 2686 15600
rect 2742 15544 6826 15600
rect 6882 15544 6887 15600
rect 2681 15542 6887 15544
rect 2681 15539 2747 15542
rect 6821 15539 6887 15542
rect 10317 15602 10383 15605
rect 14457 15602 14523 15605
rect 10317 15600 14523 15602
rect 10317 15544 10322 15600
rect 10378 15544 14462 15600
rect 14518 15544 14523 15600
rect 10317 15542 14523 15544
rect 10317 15539 10383 15542
rect 14457 15539 14523 15542
rect 0 15406 2560 15466
rect 2865 15466 2931 15469
rect 7005 15466 7071 15469
rect 2865 15464 7071 15466
rect 2865 15408 2870 15464
rect 2926 15408 7010 15464
rect 7066 15408 7071 15464
rect 2865 15406 7071 15408
rect 0 15376 480 15406
rect 2865 15403 2931 15406
rect 7005 15403 7071 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 2681 15194 2747 15197
rect 5257 15194 5323 15197
rect 2681 15192 5323 15194
rect 2681 15136 2686 15192
rect 2742 15136 5262 15192
rect 5318 15136 5323 15192
rect 2681 15134 5323 15136
rect 2681 15131 2747 15134
rect 5257 15131 5323 15134
rect 6085 15194 6151 15197
rect 9949 15194 10015 15197
rect 6085 15192 10015 15194
rect 6085 15136 6090 15192
rect 6146 15136 9954 15192
rect 10010 15136 10015 15192
rect 6085 15134 10015 15136
rect 6085 15131 6151 15134
rect 9949 15131 10015 15134
rect 3969 15058 4035 15061
rect 15745 15058 15811 15061
rect 3969 15056 15811 15058
rect 3969 15000 3974 15056
rect 4030 15000 15750 15056
rect 15806 15000 15811 15056
rect 3969 14998 15811 15000
rect 3969 14995 4035 14998
rect 15745 14995 15811 14998
rect 0 14922 480 14952
rect 3918 14922 3924 14924
rect 0 14862 3924 14922
rect 0 14832 480 14862
rect 3918 14860 3924 14862
rect 3988 14860 3994 14924
rect 7557 14922 7623 14925
rect 7925 14922 7991 14925
rect 10685 14922 10751 14925
rect 7557 14920 10751 14922
rect 7557 14864 7562 14920
rect 7618 14864 7930 14920
rect 7986 14864 10690 14920
rect 10746 14864 10751 14920
rect 7557 14862 10751 14864
rect 7557 14859 7623 14862
rect 7925 14859 7991 14862
rect 10685 14859 10751 14862
rect 4613 14786 4679 14789
rect 7189 14786 7255 14789
rect 4613 14784 7255 14786
rect 4613 14728 4618 14784
rect 4674 14728 7194 14784
rect 7250 14728 7255 14784
rect 4613 14726 7255 14728
rect 4613 14723 4679 14726
rect 7189 14723 7255 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3601 14650 3667 14653
rect 8753 14650 8819 14653
rect 3601 14648 8819 14650
rect 3601 14592 3606 14648
rect 3662 14592 8758 14648
rect 8814 14592 8819 14648
rect 3601 14590 8819 14592
rect 3601 14587 3667 14590
rect 8753 14587 8819 14590
rect 5257 14514 5323 14517
rect 6361 14514 6427 14517
rect 24117 14514 24183 14517
rect 5257 14512 24183 14514
rect 5257 14456 5262 14512
rect 5318 14456 6366 14512
rect 6422 14456 24122 14512
rect 24178 14456 24183 14512
rect 5257 14454 24183 14456
rect 5257 14451 5323 14454
rect 6361 14451 6427 14454
rect 24117 14451 24183 14454
rect 0 14378 480 14408
rect 3969 14378 4035 14381
rect 0 14376 4035 14378
rect 0 14320 3974 14376
rect 4030 14320 4035 14376
rect 0 14318 4035 14320
rect 0 14288 480 14318
rect 3969 14315 4035 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6085 14106 6151 14109
rect 11329 14106 11395 14109
rect 6085 14104 11395 14106
rect 6085 14048 6090 14104
rect 6146 14048 11334 14104
rect 11390 14048 11395 14104
rect 6085 14046 11395 14048
rect 6085 14043 6151 14046
rect 11329 14043 11395 14046
rect 4981 13970 5047 13973
rect 10133 13970 10199 13973
rect 4981 13968 10199 13970
rect 4981 13912 4986 13968
rect 5042 13912 10138 13968
rect 10194 13912 10199 13968
rect 4981 13910 10199 13912
rect 4981 13907 5047 13910
rect 10133 13907 10199 13910
rect 0 13698 480 13728
rect 9765 13698 9831 13701
rect 0 13696 9831 13698
rect 0 13640 9770 13696
rect 9826 13640 9831 13696
rect 0 13638 9831 13640
rect 0 13608 480 13638
rect 9765 13635 9831 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 2405 13426 2471 13429
rect 7649 13426 7715 13429
rect 2405 13424 7715 13426
rect 2405 13368 2410 13424
rect 2466 13368 7654 13424
rect 7710 13368 7715 13424
rect 2405 13366 7715 13368
rect 2405 13363 2471 13366
rect 7649 13363 7715 13366
rect 2221 13290 2287 13293
rect 5441 13290 5507 13293
rect 2221 13288 5507 13290
rect 2221 13232 2226 13288
rect 2282 13232 5446 13288
rect 5502 13232 5507 13288
rect 2221 13230 5507 13232
rect 2221 13227 2287 13230
rect 5441 13227 5507 13230
rect 5993 13290 6059 13293
rect 11237 13290 11303 13293
rect 5993 13288 11303 13290
rect 5993 13232 5998 13288
rect 6054 13232 11242 13288
rect 11298 13232 11303 13288
rect 5993 13230 11303 13232
rect 5993 13227 6059 13230
rect 11237 13227 11303 13230
rect 0 13154 480 13184
rect 0 13094 4906 13154
rect 0 13064 480 13094
rect 4846 12746 4906 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6545 12882 6611 12885
rect 11053 12882 11119 12885
rect 6545 12880 11119 12882
rect 6545 12824 6550 12880
rect 6606 12824 11058 12880
rect 11114 12824 11119 12880
rect 6545 12822 11119 12824
rect 6545 12819 6611 12822
rect 11053 12819 11119 12822
rect 13353 12746 13419 12749
rect 4846 12744 13419 12746
rect 4846 12688 13358 12744
rect 13414 12688 13419 12744
rect 4846 12686 13419 12688
rect 13353 12683 13419 12686
rect 4429 12610 4495 12613
rect 4705 12610 4771 12613
rect 9029 12610 9095 12613
rect 4429 12608 9095 12610
rect 4429 12552 4434 12608
rect 4490 12552 4710 12608
rect 4766 12552 9034 12608
rect 9090 12552 9095 12608
rect 4429 12550 9095 12552
rect 4429 12547 4495 12550
rect 4705 12547 4771 12550
rect 9029 12547 9095 12550
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 9857 12474 9923 12477
rect 0 12472 9923 12474
rect 0 12416 9862 12472
rect 9918 12416 9923 12472
rect 0 12414 9923 12416
rect 0 12384 480 12414
rect 9857 12411 9923 12414
rect 4061 12338 4127 12341
rect 7097 12338 7163 12341
rect 4061 12336 7163 12338
rect 4061 12280 4066 12336
rect 4122 12280 7102 12336
rect 7158 12280 7163 12336
rect 4061 12278 7163 12280
rect 4061 12275 4127 12278
rect 7097 12275 7163 12278
rect 7925 12338 7991 12341
rect 15653 12338 15719 12341
rect 7925 12336 15719 12338
rect 7925 12280 7930 12336
rect 7986 12280 15658 12336
rect 15714 12280 15719 12336
rect 7925 12278 15719 12280
rect 7925 12275 7991 12278
rect 15653 12275 15719 12278
rect 8477 12202 8543 12205
rect 11329 12202 11395 12205
rect 4846 12142 6056 12202
rect 0 11930 480 11960
rect 4846 11930 4906 12142
rect 5996 12066 6056 12142
rect 8477 12200 11395 12202
rect 8477 12144 8482 12200
rect 8538 12144 11334 12200
rect 11390 12144 11395 12200
rect 8477 12142 11395 12144
rect 8477 12139 8543 12142
rect 11329 12139 11395 12142
rect 10685 12066 10751 12069
rect 5996 12064 10751 12066
rect 5996 12008 10690 12064
rect 10746 12008 10751 12064
rect 5996 12006 10751 12008
rect 10685 12003 10751 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11870 4906 11930
rect 6269 11930 6335 11933
rect 10685 11930 10751 11933
rect 6269 11928 10751 11930
rect 6269 11872 6274 11928
rect 6330 11872 10690 11928
rect 10746 11872 10751 11928
rect 6269 11870 10751 11872
rect 0 11840 480 11870
rect 6269 11867 6335 11870
rect 10685 11867 10751 11870
rect 7741 11794 7807 11797
rect 10225 11794 10291 11797
rect 7741 11792 10291 11794
rect 7741 11736 7746 11792
rect 7802 11736 10230 11792
rect 10286 11736 10291 11792
rect 7741 11734 10291 11736
rect 7741 11731 7807 11734
rect 10225 11731 10291 11734
rect 3972 11598 9690 11658
rect 3972 11522 4032 11598
rect 9630 11556 9690 11598
rect 9630 11525 9736 11556
rect 3742 11462 4032 11522
rect 5349 11522 5415 11525
rect 8385 11522 8451 11525
rect 5349 11520 8451 11522
rect 5349 11464 5354 11520
rect 5410 11464 8390 11520
rect 8446 11464 8451 11520
rect 9630 11520 9739 11525
rect 9630 11496 9678 11520
rect 5349 11462 8451 11464
rect 0 11250 480 11280
rect 3742 11250 3802 11462
rect 5349 11459 5415 11462
rect 8385 11459 8451 11462
rect 9673 11464 9678 11496
rect 9734 11464 9739 11520
rect 9673 11459 9739 11464
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3877 11386 3943 11389
rect 5809 11386 5875 11389
rect 3877 11384 5875 11386
rect 3877 11328 3882 11384
rect 3938 11328 5814 11384
rect 5870 11328 5875 11384
rect 3877 11326 5875 11328
rect 3877 11323 3943 11326
rect 5809 11323 5875 11326
rect 0 11190 3802 11250
rect 4705 11250 4771 11253
rect 10685 11250 10751 11253
rect 12709 11250 12775 11253
rect 4705 11248 10426 11250
rect 4705 11192 4710 11248
rect 4766 11192 10426 11248
rect 4705 11190 10426 11192
rect 0 11160 480 11190
rect 4705 11187 4771 11190
rect 10133 11114 10199 11117
rect 4846 11112 10199 11114
rect 4846 11056 10138 11112
rect 10194 11056 10199 11112
rect 4846 11054 10199 11056
rect 10366 11114 10426 11190
rect 10685 11248 12775 11250
rect 10685 11192 10690 11248
rect 10746 11192 12714 11248
rect 12770 11192 12775 11248
rect 10685 11190 12775 11192
rect 10685 11187 10751 11190
rect 12709 11187 12775 11190
rect 14825 11114 14891 11117
rect 10366 11112 14891 11114
rect 10366 11056 14830 11112
rect 14886 11056 14891 11112
rect 10366 11054 14891 11056
rect 0 10706 480 10736
rect 4846 10706 4906 11054
rect 10133 11051 10199 11054
rect 14825 11051 14891 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10646 4906 10706
rect 0 10616 480 10646
rect 5717 10570 5783 10573
rect 12433 10570 12499 10573
rect 5717 10568 12499 10570
rect 5717 10512 5722 10568
rect 5778 10512 12438 10568
rect 12494 10512 12499 10568
rect 5717 10510 12499 10512
rect 5717 10507 5783 10510
rect 12433 10507 12499 10510
rect 1761 10434 1827 10437
rect 6453 10434 6519 10437
rect 1761 10432 6519 10434
rect 1761 10376 1766 10432
rect 1822 10376 6458 10432
rect 6514 10376 6519 10432
rect 1761 10374 6519 10376
rect 1761 10371 1827 10374
rect 6453 10371 6519 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3785 10298 3851 10301
rect 8293 10298 8359 10301
rect 3785 10296 8359 10298
rect 3785 10240 3790 10296
rect 3846 10240 8298 10296
rect 8354 10240 8359 10296
rect 3785 10238 8359 10240
rect 3785 10235 3851 10238
rect 8293 10235 8359 10238
rect 2589 10162 2655 10165
rect 8109 10162 8175 10165
rect 2589 10160 8175 10162
rect 2589 10104 2594 10160
rect 2650 10104 8114 10160
rect 8170 10104 8175 10160
rect 2589 10102 8175 10104
rect 2589 10099 2655 10102
rect 8109 10099 8175 10102
rect 0 10026 480 10056
rect 3785 10026 3851 10029
rect 0 10024 3851 10026
rect 0 9968 3790 10024
rect 3846 9968 3851 10024
rect 0 9966 3851 9968
rect 0 9936 480 9966
rect 3785 9963 3851 9966
rect 5257 10026 5323 10029
rect 7373 10026 7439 10029
rect 5257 10024 7439 10026
rect 5257 9968 5262 10024
rect 5318 9968 7378 10024
rect 7434 9968 7439 10024
rect 5257 9966 7439 9968
rect 5257 9963 5323 9966
rect 7373 9963 7439 9966
rect 5993 9890 6059 9893
rect 7833 9890 7899 9893
rect 9673 9890 9739 9893
rect 5993 9888 9739 9890
rect 5993 9832 5998 9888
rect 6054 9832 7838 9888
rect 7894 9832 9678 9888
rect 9734 9832 9739 9888
rect 5993 9830 9739 9832
rect 5993 9827 6059 9830
rect 7833 9827 7899 9830
rect 9673 9827 9739 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9482 480 9512
rect 3969 9482 4035 9485
rect 0 9480 4035 9482
rect 0 9424 3974 9480
rect 4030 9424 4035 9480
rect 0 9422 4035 9424
rect 0 9392 480 9422
rect 3969 9419 4035 9422
rect 9029 9482 9095 9485
rect 9029 9480 14106 9482
rect 9029 9424 9034 9480
rect 9090 9424 14106 9480
rect 9029 9422 14106 9424
rect 9029 9419 9095 9422
rect 10685 9346 10751 9349
rect 13905 9346 13971 9349
rect 10685 9344 13971 9346
rect 10685 9288 10690 9344
rect 10746 9288 13910 9344
rect 13966 9288 13971 9344
rect 10685 9286 13971 9288
rect 14046 9346 14106 9422
rect 14273 9346 14339 9349
rect 14046 9344 14339 9346
rect 14046 9288 14278 9344
rect 14334 9288 14339 9344
rect 14046 9286 14339 9288
rect 10685 9283 10751 9286
rect 13905 9283 13971 9286
rect 14273 9283 14339 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 10685 9210 10751 9213
rect 13261 9210 13327 9213
rect 10685 9208 13327 9210
rect 10685 9152 10690 9208
rect 10746 9152 13266 9208
rect 13322 9152 13327 9208
rect 10685 9150 13327 9152
rect 10685 9147 10751 9150
rect 13261 9147 13327 9150
rect 5073 9074 5139 9077
rect 10225 9074 10291 9077
rect 23473 9074 23539 9077
rect 5073 9072 23539 9074
rect 5073 9016 5078 9072
rect 5134 9016 10230 9072
rect 10286 9016 23478 9072
rect 23534 9016 23539 9072
rect 5073 9014 23539 9016
rect 5073 9011 5139 9014
rect 10225 9011 10291 9014
rect 23473 9011 23539 9014
rect 0 8802 480 8832
rect 3877 8802 3943 8805
rect 0 8800 3943 8802
rect 0 8744 3882 8800
rect 3938 8744 3943 8800
rect 0 8742 3943 8744
rect 0 8712 480 8742
rect 3877 8739 3943 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 3877 8394 3943 8397
rect 5533 8394 5599 8397
rect 3877 8392 5599 8394
rect 3877 8336 3882 8392
rect 3938 8336 5538 8392
rect 5594 8336 5599 8392
rect 3877 8334 5599 8336
rect 3877 8331 3943 8334
rect 5533 8331 5599 8334
rect 5717 8394 5783 8397
rect 6085 8394 6151 8397
rect 8569 8394 8635 8397
rect 5717 8392 8635 8394
rect 5717 8336 5722 8392
rect 5778 8336 6090 8392
rect 6146 8336 8574 8392
rect 8630 8336 8635 8392
rect 5717 8334 8635 8336
rect 5717 8331 5783 8334
rect 6085 8331 6151 8334
rect 8569 8331 8635 8334
rect 0 8258 480 8288
rect 5533 8258 5599 8261
rect 0 8256 5599 8258
rect 0 8200 5538 8256
rect 5594 8200 5599 8256
rect 0 8198 5599 8200
rect 0 8168 480 8198
rect 5533 8195 5599 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 7741 7986 7807 7989
rect 13077 7986 13143 7989
rect 7741 7984 13143 7986
rect 7741 7928 7746 7984
rect 7802 7928 13082 7984
rect 13138 7928 13143 7984
rect 7741 7926 13143 7928
rect 7741 7923 7807 7926
rect 13077 7923 13143 7926
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 480 7518
rect 1577 7515 1643 7518
rect 1669 7442 1735 7445
rect 5717 7442 5783 7445
rect 1669 7440 5783 7442
rect 1669 7384 1674 7440
rect 1730 7384 5722 7440
rect 5778 7384 5783 7440
rect 1669 7382 5783 7384
rect 1669 7379 1735 7382
rect 5717 7379 5783 7382
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2865 7034 2931 7037
rect 0 7032 2931 7034
rect 0 6976 2870 7032
rect 2926 6976 2931 7032
rect 0 6974 2931 6976
rect 0 6944 480 6974
rect 2865 6971 2931 6974
rect 23473 7034 23539 7037
rect 27520 7034 28000 7064
rect 23473 7032 28000 7034
rect 23473 6976 23478 7032
rect 23534 6976 28000 7032
rect 23473 6974 28000 6976
rect 23473 6971 23539 6974
rect 27520 6944 28000 6974
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 2681 6354 2747 6357
rect 0 6352 2747 6354
rect 0 6296 2686 6352
rect 2742 6296 2747 6352
rect 0 6294 2747 6296
rect 0 6264 480 6294
rect 2681 6291 2747 6294
rect 10685 6354 10751 6357
rect 23197 6354 23263 6357
rect 10685 6352 23263 6354
rect 10685 6296 10690 6352
rect 10746 6296 23202 6352
rect 23258 6296 23263 6352
rect 10685 6294 23263 6296
rect 10685 6291 10751 6294
rect 23197 6291 23263 6294
rect 2037 6218 2103 6221
rect 9765 6218 9831 6221
rect 2037 6216 9831 6218
rect 2037 6160 2042 6216
rect 2098 6160 9770 6216
rect 9826 6160 9831 6216
rect 2037 6158 9831 6160
rect 2037 6155 2103 6158
rect 9765 6155 9831 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1945 5946 2011 5949
rect 3049 5946 3115 5949
rect 4245 5946 4311 5949
rect 1945 5944 4311 5946
rect 1945 5888 1950 5944
rect 2006 5888 3054 5944
rect 3110 5888 4250 5944
rect 4306 5888 4311 5944
rect 1945 5886 4311 5888
rect 1945 5883 2011 5886
rect 3049 5883 3115 5886
rect 4245 5883 4311 5886
rect 0 5810 480 5840
rect 3601 5810 3667 5813
rect 0 5808 3667 5810
rect 0 5752 3606 5808
rect 3662 5752 3667 5808
rect 0 5750 3667 5752
rect 0 5720 480 5750
rect 3601 5747 3667 5750
rect 4705 5810 4771 5813
rect 12801 5810 12867 5813
rect 4705 5808 12867 5810
rect 4705 5752 4710 5808
rect 4766 5752 12806 5808
rect 12862 5752 12867 5808
rect 4705 5750 12867 5752
rect 4705 5747 4771 5750
rect 12801 5747 12867 5750
rect 2497 5674 2563 5677
rect 6913 5674 6979 5677
rect 2497 5672 6979 5674
rect 2497 5616 2502 5672
rect 2558 5616 6918 5672
rect 6974 5616 6979 5672
rect 2497 5614 6979 5616
rect 2497 5611 2563 5614
rect 6913 5611 6979 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5130 480 5160
rect 4245 5130 4311 5133
rect 0 5128 4311 5130
rect 0 5072 4250 5128
rect 4306 5072 4311 5128
rect 0 5070 4311 5072
rect 0 5040 480 5070
rect 4245 5067 4311 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4586 480 4616
rect 3141 4586 3207 4589
rect 11329 4586 11395 4589
rect 0 4584 3207 4586
rect 0 4528 3146 4584
rect 3202 4528 3207 4584
rect 0 4526 3207 4528
rect 0 4496 480 4526
rect 3141 4523 3207 4526
rect 5398 4584 11395 4586
rect 5398 4528 11334 4584
rect 11390 4528 11395 4584
rect 5398 4526 11395 4528
rect 2037 4450 2103 4453
rect 5398 4450 5458 4526
rect 11329 4523 11395 4526
rect 2037 4448 5458 4450
rect 2037 4392 2042 4448
rect 2098 4392 5458 4448
rect 2037 4390 5458 4392
rect 2037 4387 2103 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 2957 4042 3023 4045
rect 5165 4042 5231 4045
rect 2957 4040 5231 4042
rect 2957 3984 2962 4040
rect 3018 3984 5170 4040
rect 5226 3984 5231 4040
rect 2957 3982 5231 3984
rect 2957 3979 3023 3982
rect 5165 3979 5231 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2221 3498 2287 3501
rect 7005 3498 7071 3501
rect 2221 3496 7071 3498
rect 2221 3440 2226 3496
rect 2282 3440 7010 3496
rect 7066 3440 7071 3496
rect 2221 3438 7071 3440
rect 2221 3435 2287 3438
rect 7005 3435 7071 3438
rect 0 3362 480 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 480 3302
rect 2865 3299 2931 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1393 2682 1459 2685
rect 0 2680 1459 2682
rect 0 2624 1398 2680
rect 1454 2624 1459 2680
rect 0 2622 1459 2624
rect 0 2592 480 2622
rect 1393 2619 1459 2622
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 2681 2138 2747 2141
rect 0 2136 2747 2138
rect 0 2080 2686 2136
rect 2742 2080 2747 2136
rect 0 2078 2747 2080
rect 0 2048 480 2078
rect 2681 2075 2747 2078
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 0 914 480 944
rect 4245 914 4311 917
rect 0 912 4311 914
rect 0 856 4250 912
rect 4306 856 4311 912
rect 0 854 4311 856
rect 0 824 480 854
rect 4245 851 4311 854
rect 0 370 480 400
rect 3049 370 3115 373
rect 0 368 3115 370
rect 0 312 3054 368
rect 3110 312 3115 368
rect 0 310 3115 312
rect 0 280 480 310
rect 3049 307 3115 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 9628 20300 9692 20364
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 9628 19348 9692 19412
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 15516 18048 15580 18052
rect 15516 17992 15566 18048
rect 15566 17992 15580 18048
rect 15516 17988 15580 17992
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 3924 14860 3988 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9627 20364 9693 20365
rect 9627 20300 9628 20364
rect 9692 20300 9693 20364
rect 9627 20299 9693 20300
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 9630 19413 9690 20299
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9627 19412 9693 19413
rect 9627 19348 9628 19412
rect 9692 19348 9693 19412
rect 9627 19347 9693 19348
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 3923 14924 3989 14925
rect 3923 14860 3924 14924
rect 3988 14860 3989 14924
rect 3923 14859 3989 14860
rect 3926 14738 3986 14859
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 15518 14738 15578 17987
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 3838 14502 4074 14738
rect 15430 14502 15666 14738
<< metal5 >>
rect 3796 14738 15708 14780
rect 3796 14502 3838 14738
rect 4074 14502 15430 14738
rect 15666 14502 15708 14738
rect 3796 14460 15708 14502
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _086_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_19
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_37 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_40
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_52
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_49
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_60
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_buf_4  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_13
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_25
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_45
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_21
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_28
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 590 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_13
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_42
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _056_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_buf_4  mux_left_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_12
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_57
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 1786 592
use scs8hd_buf_4  mux_left_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_26
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_buf_4  mux_left_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_9
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_13
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_25
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _067_
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _058_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_77
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_8  FILLER_16_118
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _066_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_116
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_16
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_12
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_26
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 1786 592
use scs8hd_buf_4  mux_left_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_33
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_50
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_67
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_26
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_139
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_34
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_24
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_6  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_38.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_113
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_160
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 866 592
use scs8hd_buf_4  mux_left_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_9
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_13
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_26
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 314 592
use scs8hd_conb_1  _062_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_38.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 130 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_36.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_48
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_28.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_89
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_99
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_30.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_106
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_103
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_30.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_36.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_238
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_38
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_118
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_173
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_200
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_4  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_223
timestamp 1586364061
transform 1 0 21620 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_242
timestamp 1586364061
transform 1 0 23368 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_254
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_266
timestamp 1586364061
transform 1 0 25576 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_52
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_128
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_155
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_34.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_30.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 590 592
use scs8hd_decap_6  FILLER_29_237
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_243
timestamp 1586364061
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_54
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_28.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11776 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_115
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_34.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_146
timestamp 1586364061
transform 1 0 14536 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_171
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_30_179
timestamp 1586364061
transform 1 0 17572 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 22724 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_221
timestamp 1586364061
transform 1 0 21436 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_233
timestamp 1586364061
transform 1 0 22540 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 1786 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4508 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_33
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_65
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_100
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_128
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 130 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 1786 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_28.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_203
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_207
timestamp 1586364061
transform 1 0 20148 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_218
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 21896 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_238
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4140 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_42
timestamp 1586364061
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_78
timestamp 1586364061
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_82
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_97
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_118
timestamp 1586364061
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_122
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_158
timestamp 1586364061
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_162
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18124 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_187
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_191
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 406 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 21068 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 22264 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_221
timestamp 1586364061
transform 1 0 21436 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_229
timestamp 1586364061
transform 1 0 22172 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_234
timestamp 1586364061
transform 1 0 22632 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_246
timestamp 1586364061
transform 1 0 23736 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_258
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_270
timestamp 1586364061
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_26
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_34_49
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_87
timestamp 1586364061
transform 1 0 9108 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_98
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_164
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_181
timestamp 1586364061
transform 1 0 17756 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_195
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 590 592
use scs8hd_decap_6  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_211
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_207
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 590 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_221
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_225
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_219
timestamp 1586364061
transform 1 0 21252 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_231
timestamp 1586364061
transform 1 0 22356 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_255
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 1786 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_8
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_116
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 590 592
use scs8hd_buf_4  mux_top_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_172
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_176
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_190
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_194
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_202
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_214
timestamp 1586364061
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_10
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4692 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_41
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_71
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_82
timestamp 1586364061
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_86
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13524 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_127
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_148
timestamp 1586364061
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16744 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_162
timestamp 1586364061
transform 1 0 16008 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_36_176
timestamp 1586364061
transform 1 0 17296 0 -1 22304
box -38 -48 774 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_18
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_85
timestamp 1586364061
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_170
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_174
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 590 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 406 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19688 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_216
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_34.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_249
timestamp 1586364061
transform 1 0 24012 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_261
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_273
timestamp 1586364061
transform 1 0 26220 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1786 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3312 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_22
timestamp 1586364061
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_26
timestamp 1586364061
transform 1 0 3496 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_51
timestamp 1586364061
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_55
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_78
timestamp 1586364061
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_86
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_90
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_112
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12144 0 -1 23392
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_139
timestamp 1586364061
transform 1 0 13892 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_38_151
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_160
timestamp 1586364061
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_164
timestamp 1586364061
transform 1 0 16192 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_172
timestamp 1586364061
transform 1 0 16928 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 406 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_184
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_192
timestamp 1586364061
transform 1 0 18768 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_197
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_209
timestamp 1586364061
transform 1 0 20332 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_36.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_237
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_4  mux_top_track_38.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_11
timestamp 1586364061
transform 1 0 2116 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_36
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_40
timestamp 1586364061
transform 1 0 4784 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_50
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_40_78
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_121
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_134
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_138
timestamp 1586364061
transform 1 0 13800 0 -1 24480
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 590 592
use scs8hd_buf_4  mux_top_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_153
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_160
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_172
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_184
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_196
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_208
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21620 0 -1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_242
timestamp 1586364061
transform 1 0 23368 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_256
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_252
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 23920 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_254
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_266
timestamp 1586364061
transform 1 0 25576 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_264
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_268
timestamp 1586364061
transform 1 0 25760 0 1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_276
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_31
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 5428 0 1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_41_43
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_41_50
timestamp 1586364061
transform 1 0 5704 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_41_58
timestamp 1586364061
transform 1 0 6440 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_41_70
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_90
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_96
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_107
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_111
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_115
timestamp 1586364061
transform 1 0 11684 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12512 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_133
timestamp 1586364061
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_137
timestamp 1586364061
transform 1 0 13708 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14076 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2760 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_12
timestamp 1586364061
transform 1 0 2208 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_16
timestamp 1586364061
transform 1 0 2576 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_20
timestamp 1586364061
transform 1 0 2944 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_24
timestamp 1586364061
transform 1 0 3312 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_30
timestamp 1586364061
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_89
timestamp 1586364061
transform 1 0 9292 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_115
timestamp 1586364061
transform 1 0 11684 0 -1 25568
box -38 -48 774 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_123
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_128
timestamp 1586364061
transform 1 0 12880 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_140
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_42_152
timestamp 1586364061
transform 1 0 15088 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 27618 27520 27674 28000 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 25168 480 25288 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 19728 480 19848 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 20272 480 20392 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 20952 480 21072 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 21496 480 21616 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 22176 480 22296 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 22720 480 22840 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 23400 480 23520 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 23944 480 24064 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 24624 480 24744 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 17280 480 17400 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 10616 480 10736 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4710 27520 4766 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10322 27520 10378 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5262 27520 5318 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8666 27520 8722 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9218 27520 9274 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16486 27520 16542 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18142 27520 18198 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19246 27520 19302 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 82 nsew default input
rlabel metal2 s 4618 0 4674 480 6 left_top_grid_pin_42_
port 83 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_43_
port 84 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 left_top_grid_pin_44_
port 85 nsew default input
rlabel metal2 s 13910 0 13966 480 6 left_top_grid_pin_45_
port 86 nsew default input
rlabel metal3 s 0 26392 480 26512 6 left_top_grid_pin_46_
port 87 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_47_
port 88 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_48_
port 89 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 left_top_grid_pin_49_
port 90 nsew default input
rlabel metal2 s 23202 0 23258 480 6 prog_clk
port 91 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 92 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 93 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 94 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_37_
port 95 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_38_
port 96 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 top_left_grid_pin_39_
port 97 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 top_left_grid_pin_40_
port 98 nsew default input
rlabel metal2 s 4158 27520 4214 28000 6 top_left_grid_pin_41_
port 99 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 101 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
